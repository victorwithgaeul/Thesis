// Product (AN) Code SEC l-LUT
// SEC_lLUT52bits.v
// Received single error location l, output remainder r.
module SEC_lLUT52bits(l, r);
input	signed	[7:0]	l;
output	reg	[15:0]	r;
always@(*) begin
	case(l)
		1: r = 1;
		-1: r = 50860;
		2: r = 2;
		-2: r = 50859;
		3: r = 4;
		-3: r = 50857;
		4: r = 8;
		-4: r = 50853;
		5: r = 16;
		-5: r = 50845;
		6: r = 32;
		-6: r = 50829;
		7: r = 64;
		-7: r = 50797;
		8: r = 128;
		-8: r = 50733;
		9: r = 256;
		-9: r = 50605;
		10: r = 512;
		-10: r = 50349;
		11: r = 1024;
		-11: r = 49837;
		12: r = 2048;
		-12: r = 48813;
		13: r = 4096;
		-13: r = 46765;
		14: r = 8192;
		-14: r = 42669;
		15: r = 16384;
		-15: r = 34477;
		16: r = 32768;
		-16: r = 18093;
		17: r = 14675;
		-17: r = 36186;
		18: r = 29350;
		-18: r = 21511;
		19: r = 7839;
		-19: r = 43022;
		20: r = 15678;
		-20: r = 35183;
		21: r = 31356;
		-21: r = 19505;
		22: r = 11851;
		-22: r = 39010;
		23: r = 23702;
		-23: r = 27159;
		24: r = 47404;
		-24: r = 3457;
		25: r = 43947;
		-25: r = 6914;
		26: r = 37033;
		-26: r = 13828;
		27: r = 23205;
		-27: r = 27656;
		28: r = 46410;
		-28: r = 4451;
		29: r = 41959;
		-29: r = 8902;
		30: r = 33057;
		-30: r = 17804;
		31: r = 15253;
		-31: r = 35608;
		32: r = 30506;
		-32: r = 20355;
		33: r = 10151;
		-33: r = 40710;
		34: r = 20302;
		-34: r = 30559;
		35: r = 40604;
		-35: r = 10257;
		36: r = 30347;
		-36: r = 20514;
		37: r = 9833;
		-37: r = 41028;
		38: r = 19666;
		-38: r = 31195;
		39: r = 39332;
		-39: r = 11529;
		40: r = 27803;
		-40: r = 23058;
		41: r = 4745;
		-41: r = 46116;
		42: r = 9490;
		-42: r = 41371;
		43: r = 18980;
		-43: r = 31881;
		44: r = 37960;
		-44: r = 12901;
		45: r = 25059;
		-45: r = 25802;
		46: r = 50118;
		-46: r = 743;
		47: r = 49375;
		-47: r = 1486;
		48: r = 47889;
		-48: r = 2972;
		49: r = 44917;
		-49: r = 5944;
		50: r = 38973;
		-50: r = 11888;
		51: r = 27085;
		-51: r = 23776;
		52: r = 3309;
		-52: r = 47552;
		53: r = 6618;
		-53: r = 44243;
		54: r = 13236;
		-54: r = 37625;
		55: r = 26472;
		-55: r = 24389;
		56: r = 2083;
		-56: r = 48778;
		57: r = 4166;
		-57: r = 46695;
		58: r = 8332;
		-58: r = 42529;
		59: r = 16664;
		-59: r = 34197;
		60: r = 33328;
		-60: r = 17533;
		61: r = 15795;
		-61: r = 35066;
		62: r = 31590;
		-62: r = 19271;
		63: r = 12319;
		-63: r = 38542;
		64: r = 24638;
		-64: r = 26223;
		65: r = 49276;
		-65: r = 1585;
		66: r = 47691;
		-66: r = 3170;
		67: r = 44521;
		-67: r = 6340;
		68: r = 38181;
		-68: r = 12680;
		default: r = 0;
	endcase
end

endmodule

// Product (AN) Code SEC_LUT_Decoder
// SEC_LUT_Decoder30bits.v
// Received codeword W = AN + e, e is single arithmetic weight error (AWE), +2^i or -2^i.
module SEC_LUT_Decoder30bits(W, N);
input 	[44:0]	W;
output	[29:0]	N;
parameter A = 18613;

wire 	[29:0]	Q;
wire 	[14:0]	R;
assign Q = W / A;
assign R = W - (A * Q);

reg	signed	[45:0]	Delta;
always@(*) begin
	case(R)
		1: Delta = 46'sb0000000000000000000000000000000000000000000001;
		18612: Delta = 46'sb1111111111111111111111111111111111111111111111;
		2: Delta = 46'sb0000000000000000000000000000000000000000000010;
		18611: Delta = 46'sb1111111111111111111111111111111111111111111110;
		4: Delta = 46'sb0000000000000000000000000000000000000000000100;
		18609: Delta = 46'sb1111111111111111111111111111111111111111111100;
		8: Delta = 46'sb0000000000000000000000000000000000000000001000;
		18605: Delta = 46'sb1111111111111111111111111111111111111111111000;
		16: Delta = 46'sb0000000000000000000000000000000000000000010000;
		18597: Delta = 46'sb1111111111111111111111111111111111111111110000;
		32: Delta = 46'sb0000000000000000000000000000000000000000100000;
		18581: Delta = 46'sb1111111111111111111111111111111111111111100000;
		64: Delta = 46'sb0000000000000000000000000000000000000001000000;
		18549: Delta = 46'sb1111111111111111111111111111111111111111000000;
		128: Delta = 46'sb0000000000000000000000000000000000000010000000;
		18485: Delta = 46'sb1111111111111111111111111111111111111110000000;
		256: Delta = 46'sb0000000000000000000000000000000000000100000000;
		18357: Delta = 46'sb1111111111111111111111111111111111111100000000;
		512: Delta = 46'sb0000000000000000000000000000000000001000000000;
		18101: Delta = 46'sb1111111111111111111111111111111111111000000000;
		1024: Delta = 46'sb0000000000000000000000000000000000010000000000;
		17589: Delta = 46'sb1111111111111111111111111111111111110000000000;
		2048: Delta = 46'sb0000000000000000000000000000000000100000000000;
		16565: Delta = 46'sb1111111111111111111111111111111111100000000000;
		4096: Delta = 46'sb0000000000000000000000000000000001000000000000;
		14517: Delta = 46'sb1111111111111111111111111111111111000000000000;
		8192: Delta = 46'sb0000000000000000000000000000000010000000000000;
		10421: Delta = 46'sb1111111111111111111111111111111110000000000000;
		16384: Delta = 46'sb0000000000000000000000000000000100000000000000;
		2229: Delta = 46'sb1111111111111111111111111111111100000000000000;
		14155: Delta = 46'sb0000000000000000000000000000001000000000000000;
		4458: Delta = 46'sb1111111111111111111111111111111000000000000000;
		9697: Delta = 46'sb0000000000000000000000000000010000000000000000;
		8916: Delta = 46'sb1111111111111111111111111111110000000000000000;
		781: Delta = 46'sb0000000000000000000000000000100000000000000000;
		17832: Delta = 46'sb1111111111111111111111111111100000000000000000;
		1562: Delta = 46'sb0000000000000000000000000001000000000000000000;
		17051: Delta = 46'sb1111111111111111111111111111000000000000000000;
		3124: Delta = 46'sb0000000000000000000000000010000000000000000000;
		15489: Delta = 46'sb1111111111111111111111111110000000000000000000;
		6248: Delta = 46'sb0000000000000000000000000100000000000000000000;
		12365: Delta = 46'sb1111111111111111111111111100000000000000000000;
		12496: Delta = 46'sb0000000000000000000000001000000000000000000000;
		6117: Delta = 46'sb1111111111111111111111111000000000000000000000;
		6379: Delta = 46'sb0000000000000000000000010000000000000000000000;
		12234: Delta = 46'sb1111111111111111111111110000000000000000000000;
		12758: Delta = 46'sb0000000000000000000000100000000000000000000000;
		5855: Delta = 46'sb1111111111111111111111100000000000000000000000;
		6903: Delta = 46'sb0000000000000000000001000000000000000000000000;
		11710: Delta = 46'sb1111111111111111111111000000000000000000000000;
		13806: Delta = 46'sb0000000000000000000010000000000000000000000000;
		4807: Delta = 46'sb1111111111111111111110000000000000000000000000;
		8999: Delta = 46'sb0000000000000000000100000000000000000000000000;
		9614: Delta = 46'sb1111111111111111111100000000000000000000000000;
		17998: Delta = 46'sb0000000000000000001000000000000000000000000000;
		615: Delta = 46'sb1111111111111111111000000000000000000000000000;
		17383: Delta = 46'sb0000000000000000010000000000000000000000000000;
		1230: Delta = 46'sb1111111111111111110000000000000000000000000000;
		16153: Delta = 46'sb0000000000000000100000000000000000000000000000;
		2460: Delta = 46'sb1111111111111111100000000000000000000000000000;
		13693: Delta = 46'sb0000000000000001000000000000000000000000000000;
		4920: Delta = 46'sb1111111111111111000000000000000000000000000000;
		8773: Delta = 46'sb0000000000000010000000000000000000000000000000;
		9840: Delta = 46'sb1111111111111110000000000000000000000000000000;
		17546: Delta = 46'sb0000000000000100000000000000000000000000000000;
		1067: Delta = 46'sb1111111111111100000000000000000000000000000000;
		16479: Delta = 46'sb0000000000001000000000000000000000000000000000;
		2134: Delta = 46'sb1111111111111000000000000000000000000000000000;
		14345: Delta = 46'sb0000000000010000000000000000000000000000000000;
		4268: Delta = 46'sb1111111111110000000000000000000000000000000000;
		10077: Delta = 46'sb0000000000100000000000000000000000000000000000;
		8536: Delta = 46'sb1111111111100000000000000000000000000000000000;
		1541: Delta = 46'sb0000000001000000000000000000000000000000000000;
		17072: Delta = 46'sb1111111111000000000000000000000000000000000000;
		3082: Delta = 46'sb0000000010000000000000000000000000000000000000;
		15531: Delta = 46'sb1111111110000000000000000000000000000000000000;
		6164: Delta = 46'sb0000000100000000000000000000000000000000000000;
		12449: Delta = 46'sb1111111100000000000000000000000000000000000000;
		12328: Delta = 46'sb0000001000000000000000000000000000000000000000;
		6285: Delta = 46'sb1111111000000000000000000000000000000000000000;
		6043: Delta = 46'sb0000010000000000000000000000000000000000000000;
		12570: Delta = 46'sb1111110000000000000000000000000000000000000000;
		12086: Delta = 46'sb0000100000000000000000000000000000000000000000;
		6527: Delta = 46'sb1111100000000000000000000000000000000000000000;
		5559: Delta = 46'sb0001000000000000000000000000000000000000000000;
		13054: Delta = 46'sb1111000000000000000000000000000000000000000000;
		11118: Delta = 46'sb0010000000000000000000000000000000000000000000;
		7495: Delta = 46'sb1110000000000000000000000000000000000000000000;
		3623: Delta = 46'sb0100000000000000000000000000000000000000000000;
		14990: Delta = 46'sb1100000000000000000000000000000000000000000000;
		default: Delta =46'sb0;
	endcase
end

assign N = (W - Delta) / A;

endmodule

// Product (AN) Code DEC r-LUT
// DEC_rLUT24bits.v
// Used to do DEC, but corrected errors by locations, not AWE
// Received remainder r, output two error locations.
module DEC_rLUT24bits(r, l_1, l_2);
input 	[13:0]	r;
output	reg	signed	[6:0]	l_1;
output	reg	signed	[6:0]	l_2;
always@(*) begin
	case(r)
		1: begin l_1 = -1;
				 l_2 = +2; end
		13836: begin l_1 = +1;
				 l_2 = -2; end
		2: begin l_1 = +1;
				 l_2 = +1; end
		13835: begin l_1 = -1;
				 l_2 = -1; end
		4: begin l_1 = +2;
				 l_2 = +2; end
		13833: begin l_1 = -2;
				 l_2 = -2; end
		8: begin l_1 = +3;
				 l_2 = +3; end
		13829: begin l_1 = -3;
				 l_2 = -3; end
		16: begin l_1 = +4;
				 l_2 = +4; end
		13821: begin l_1 = -4;
				 l_2 = -4; end
		32: begin l_1 = +5;
				 l_2 = +5; end
		13805: begin l_1 = -5;
				 l_2 = -5; end
		64: begin l_1 = +6;
				 l_2 = +6; end
		13773: begin l_1 = -6;
				 l_2 = -6; end
		128: begin l_1 = +7;
				 l_2 = +7; end
		13709: begin l_1 = -7;
				 l_2 = -7; end
		256: begin l_1 = +8;
				 l_2 = +8; end
		13581: begin l_1 = -8;
				 l_2 = -8; end
		512: begin l_1 = +9;
				 l_2 = +9; end
		13325: begin l_1 = -9;
				 l_2 = -9; end
		1024: begin l_1 = +10;
				 l_2 = +10; end
		12813: begin l_1 = -10;
				 l_2 = -10; end
		2048: begin l_1 = +11;
				 l_2 = +11; end
		11789: begin l_1 = -11;
				 l_2 = -11; end
		4096: begin l_1 = +12;
				 l_2 = +12; end
		9741: begin l_1 = -12;
				 l_2 = -12; end
		8192: begin l_1 = +13;
				 l_2 = +13; end
		5645: begin l_1 = -13;
				 l_2 = -13; end
		2547: begin l_1 = +14;
				 l_2 = +14; end
		11290: begin l_1 = -14;
				 l_2 = -14; end
		5094: begin l_1 = +15;
				 l_2 = +15; end
		8743: begin l_1 = -15;
				 l_2 = -15; end
		10188: begin l_1 = +16;
				 l_2 = +16; end
		3649: begin l_1 = -16;
				 l_2 = -16; end
		6539: begin l_1 = +17;
				 l_2 = +17; end
		7298: begin l_1 = -17;
				 l_2 = -17; end
		13078: begin l_1 = +18;
				 l_2 = +18; end
		759: begin l_1 = -18;
				 l_2 = -18; end
		12319: begin l_1 = +19;
				 l_2 = +19; end
		1518: begin l_1 = -19;
				 l_2 = -19; end
		10801: begin l_1 = +20;
				 l_2 = +20; end
		3036: begin l_1 = -20;
				 l_2 = -20; end
		7765: begin l_1 = +21;
				 l_2 = +21; end
		6072: begin l_1 = -21;
				 l_2 = -21; end
		1693: begin l_1 = +22;
				 l_2 = +22; end
		12144: begin l_1 = -22;
				 l_2 = -22; end
		3386: begin l_1 = +23;
				 l_2 = +23; end
		10451: begin l_1 = -23;
				 l_2 = -23; end
		6772: begin l_1 = +24;
				 l_2 = +24; end
		7065: begin l_1 = -24;
				 l_2 = -24; end
		13544: begin l_1 = +25;
				 l_2 = +25; end
		293: begin l_1 = -25;
				 l_2 = -25; end
		13251: begin l_1 = +26;
				 l_2 = +26; end
		586: begin l_1 = -26;
				 l_2 = -26; end
		12665: begin l_1 = +27;
				 l_2 = +27; end
		1172: begin l_1 = -27;
				 l_2 = -27; end
		11493: begin l_1 = +28;
				 l_2 = +28; end
		2344: begin l_1 = -28;
				 l_2 = -28; end
		9149: begin l_1 = +29;
				 l_2 = +29; end
		4688: begin l_1 = -29;
				 l_2 = -29; end
		4461: begin l_1 = +30;
				 l_2 = +30; end
		9376: begin l_1 = -30;
				 l_2 = -30; end
		8922: begin l_1 = +31;
				 l_2 = +31; end
		4915: begin l_1 = -31;
				 l_2 = -31; end
		4007: begin l_1 = +32;
				 l_2 = +32; end
		9830: begin l_1 = -32;
				 l_2 = -32; end
		8014: begin l_1 = +33;
				 l_2 = +33; end
		5823: begin l_1 = -33;
				 l_2 = -33; end
		2191: begin l_1 = +34;
				 l_2 = +34; end
		11646: begin l_1 = -34;
				 l_2 = -34; end
		4382: begin l_1 = +35;
				 l_2 = +35; end
		9455: begin l_1 = -35;
				 l_2 = -35; end
		8764: begin l_1 = +36;
				 l_2 = +36; end
		5073: begin l_1 = -36;
				 l_2 = -36; end
		3691: begin l_1 = +37;
				 l_2 = +37; end
		10146: begin l_1 = -37;
				 l_2 = -37; end
		3: begin l_1 = -1;
				 l_2 = +3; end
		13834: begin l_1 = -1;
				 l_2 = -2; end
		5: begin l_1 = +1;
				 l_2 = +3; end
		13832: begin l_1 = -1;
				 l_2 = -3; end
		9: begin l_1 = +1;
				 l_2 = +4; end
		13830: begin l_1 = +1;
				 l_2 = -4; end
		7: begin l_1 = -1;
				 l_2 = +4; end
		13828: begin l_1 = -1;
				 l_2 = -4; end
		17: begin l_1 = +1;
				 l_2 = +5; end
		13822: begin l_1 = +1;
				 l_2 = -5; end
		15: begin l_1 = -1;
				 l_2 = +5; end
		13820: begin l_1 = -1;
				 l_2 = -5; end
		33: begin l_1 = +1;
				 l_2 = +6; end
		13806: begin l_1 = +1;
				 l_2 = -6; end
		31: begin l_1 = -1;
				 l_2 = +6; end
		13804: begin l_1 = -1;
				 l_2 = -6; end
		65: begin l_1 = +1;
				 l_2 = +7; end
		13774: begin l_1 = +1;
				 l_2 = -7; end
		63: begin l_1 = -1;
				 l_2 = +7; end
		13772: begin l_1 = -1;
				 l_2 = -7; end
		129: begin l_1 = +1;
				 l_2 = +8; end
		13710: begin l_1 = +1;
				 l_2 = -8; end
		127: begin l_1 = -1;
				 l_2 = +8; end
		13708: begin l_1 = -1;
				 l_2 = -8; end
		257: begin l_1 = +1;
				 l_2 = +9; end
		13582: begin l_1 = +1;
				 l_2 = -9; end
		255: begin l_1 = -1;
				 l_2 = +9; end
		13580: begin l_1 = -1;
				 l_2 = -9; end
		513: begin l_1 = +1;
				 l_2 = +10; end
		13326: begin l_1 = +1;
				 l_2 = -10; end
		511: begin l_1 = -1;
				 l_2 = +10; end
		13324: begin l_1 = -1;
				 l_2 = -10; end
		1025: begin l_1 = +1;
				 l_2 = +11; end
		12814: begin l_1 = +1;
				 l_2 = -11; end
		1023: begin l_1 = -1;
				 l_2 = +11; end
		12812: begin l_1 = -1;
				 l_2 = -11; end
		2049: begin l_1 = +1;
				 l_2 = +12; end
		11790: begin l_1 = +1;
				 l_2 = -12; end
		2047: begin l_1 = -1;
				 l_2 = +12; end
		11788: begin l_1 = -1;
				 l_2 = -12; end
		4097: begin l_1 = +1;
				 l_2 = +13; end
		9742: begin l_1 = +1;
				 l_2 = -13; end
		4095: begin l_1 = -1;
				 l_2 = +13; end
		9740: begin l_1 = -1;
				 l_2 = -13; end
		8193: begin l_1 = +1;
				 l_2 = +14; end
		5646: begin l_1 = +1;
				 l_2 = -14; end
		8191: begin l_1 = -1;
				 l_2 = +14; end
		5644: begin l_1 = -1;
				 l_2 = -14; end
		2548: begin l_1 = +1;
				 l_2 = +15; end
		11291: begin l_1 = +1;
				 l_2 = -15; end
		2546: begin l_1 = -1;
				 l_2 = +15; end
		11289: begin l_1 = -1;
				 l_2 = -15; end
		5095: begin l_1 = +1;
				 l_2 = +16; end
		8744: begin l_1 = +1;
				 l_2 = -16; end
		5093: begin l_1 = -1;
				 l_2 = +16; end
		8742: begin l_1 = -1;
				 l_2 = -16; end
		10189: begin l_1 = +1;
				 l_2 = +17; end
		3650: begin l_1 = +1;
				 l_2 = -17; end
		10187: begin l_1 = -1;
				 l_2 = +17; end
		3648: begin l_1 = -1;
				 l_2 = -17; end
		6540: begin l_1 = +1;
				 l_2 = +18; end
		7299: begin l_1 = +1;
				 l_2 = -18; end
		6538: begin l_1 = -1;
				 l_2 = +18; end
		7297: begin l_1 = -1;
				 l_2 = -18; end
		13079: begin l_1 = +1;
				 l_2 = +19; end
		760: begin l_1 = +1;
				 l_2 = -19; end
		13077: begin l_1 = -1;
				 l_2 = +19; end
		758: begin l_1 = -1;
				 l_2 = -19; end
		12320: begin l_1 = +1;
				 l_2 = +20; end
		1519: begin l_1 = +1;
				 l_2 = -20; end
		12318: begin l_1 = -1;
				 l_2 = +20; end
		1517: begin l_1 = -1;
				 l_2 = -20; end
		10802: begin l_1 = +1;
				 l_2 = +21; end
		3037: begin l_1 = +1;
				 l_2 = -21; end
		10800: begin l_1 = -1;
				 l_2 = +21; end
		3035: begin l_1 = -1;
				 l_2 = -21; end
		7766: begin l_1 = +1;
				 l_2 = +22; end
		6073: begin l_1 = +1;
				 l_2 = -22; end
		7764: begin l_1 = -1;
				 l_2 = +22; end
		6071: begin l_1 = -1;
				 l_2 = -22; end
		1694: begin l_1 = +1;
				 l_2 = +23; end
		12145: begin l_1 = +1;
				 l_2 = -23; end
		1692: begin l_1 = -1;
				 l_2 = +23; end
		12143: begin l_1 = -1;
				 l_2 = -23; end
		3387: begin l_1 = +1;
				 l_2 = +24; end
		10452: begin l_1 = +1;
				 l_2 = -24; end
		3385: begin l_1 = -1;
				 l_2 = +24; end
		10450: begin l_1 = -1;
				 l_2 = -24; end
		6773: begin l_1 = +1;
				 l_2 = +25; end
		7066: begin l_1 = +1;
				 l_2 = -25; end
		6771: begin l_1 = -1;
				 l_2 = +25; end
		7064: begin l_1 = -1;
				 l_2 = -25; end
		13545: begin l_1 = +1;
				 l_2 = +26; end
		294: begin l_1 = +1;
				 l_2 = -26; end
		13543: begin l_1 = -1;
				 l_2 = +26; end
		292: begin l_1 = -1;
				 l_2 = -26; end
		13252: begin l_1 = +1;
				 l_2 = +27; end
		587: begin l_1 = +1;
				 l_2 = -27; end
		13250: begin l_1 = -1;
				 l_2 = +27; end
		585: begin l_1 = -1;
				 l_2 = -27; end
		12666: begin l_1 = +1;
				 l_2 = +28; end
		1173: begin l_1 = +1;
				 l_2 = -28; end
		12664: begin l_1 = -1;
				 l_2 = +28; end
		1171: begin l_1 = -1;
				 l_2 = -28; end
		11494: begin l_1 = +1;
				 l_2 = +29; end
		2345: begin l_1 = +1;
				 l_2 = -29; end
		11492: begin l_1 = -1;
				 l_2 = +29; end
		2343: begin l_1 = -1;
				 l_2 = -29; end
		9150: begin l_1 = +1;
				 l_2 = +30; end
		4689: begin l_1 = +1;
				 l_2 = -30; end
		9148: begin l_1 = -1;
				 l_2 = +30; end
		4687: begin l_1 = -1;
				 l_2 = -30; end
		4462: begin l_1 = +1;
				 l_2 = +31; end
		9377: begin l_1 = +1;
				 l_2 = -31; end
		4460: begin l_1 = -1;
				 l_2 = +31; end
		9375: begin l_1 = -1;
				 l_2 = -31; end
		8923: begin l_1 = +1;
				 l_2 = +32; end
		4916: begin l_1 = +1;
				 l_2 = -32; end
		8921: begin l_1 = -1;
				 l_2 = +32; end
		4914: begin l_1 = -1;
				 l_2 = -32; end
		4008: begin l_1 = +1;
				 l_2 = +33; end
		9831: begin l_1 = +1;
				 l_2 = -33; end
		4006: begin l_1 = -1;
				 l_2 = +33; end
		9829: begin l_1 = -1;
				 l_2 = -33; end
		8015: begin l_1 = +1;
				 l_2 = +34; end
		5824: begin l_1 = +1;
				 l_2 = -34; end
		8013: begin l_1 = -1;
				 l_2 = +34; end
		5822: begin l_1 = -1;
				 l_2 = -34; end
		2192: begin l_1 = +1;
				 l_2 = +35; end
		11647: begin l_1 = +1;
				 l_2 = -35; end
		2190: begin l_1 = -1;
				 l_2 = +35; end
		11645: begin l_1 = -1;
				 l_2 = -35; end
		4383: begin l_1 = +1;
				 l_2 = +36; end
		9456: begin l_1 = +1;
				 l_2 = -36; end
		4381: begin l_1 = -1;
				 l_2 = +36; end
		9454: begin l_1 = -1;
				 l_2 = -36; end
		8765: begin l_1 = +1;
				 l_2 = +37; end
		5074: begin l_1 = +1;
				 l_2 = -37; end
		8763: begin l_1 = -1;
				 l_2 = +37; end
		5072: begin l_1 = -1;
				 l_2 = -37; end
		3692: begin l_1 = +1;
				 l_2 = +38; end
		10147: begin l_1 = +1;
				 l_2 = -38; end
		3690: begin l_1 = -1;
				 l_2 = +38; end
		10145: begin l_1 = -1;
				 l_2 = -38; end
		6: begin l_1 = -2;
				 l_2 = +4; end
		13831: begin l_1 = -2;
				 l_2 = -3; end
		10: begin l_1 = +2;
				 l_2 = +4; end
		13827: begin l_1 = -2;
				 l_2 = -4; end
		18: begin l_1 = +2;
				 l_2 = +5; end
		13823: begin l_1 = +2;
				 l_2 = -5; end
		14: begin l_1 = -2;
				 l_2 = +5; end
		13819: begin l_1 = -2;
				 l_2 = -5; end
		34: begin l_1 = +2;
				 l_2 = +6; end
		13807: begin l_1 = +2;
				 l_2 = -6; end
		30: begin l_1 = -2;
				 l_2 = +6; end
		13803: begin l_1 = -2;
				 l_2 = -6; end
		66: begin l_1 = +2;
				 l_2 = +7; end
		13775: begin l_1 = +2;
				 l_2 = -7; end
		62: begin l_1 = -2;
				 l_2 = +7; end
		13771: begin l_1 = -2;
				 l_2 = -7; end
		130: begin l_1 = +2;
				 l_2 = +8; end
		13711: begin l_1 = +2;
				 l_2 = -8; end
		126: begin l_1 = -2;
				 l_2 = +8; end
		13707: begin l_1 = -2;
				 l_2 = -8; end
		258: begin l_1 = +2;
				 l_2 = +9; end
		13583: begin l_1 = +2;
				 l_2 = -9; end
		254: begin l_1 = -2;
				 l_2 = +9; end
		13579: begin l_1 = -2;
				 l_2 = -9; end
		514: begin l_1 = +2;
				 l_2 = +10; end
		13327: begin l_1 = +2;
				 l_2 = -10; end
		510: begin l_1 = -2;
				 l_2 = +10; end
		13323: begin l_1 = -2;
				 l_2 = -10; end
		1026: begin l_1 = +2;
				 l_2 = +11; end
		12815: begin l_1 = +2;
				 l_2 = -11; end
		1022: begin l_1 = -2;
				 l_2 = +11; end
		12811: begin l_1 = -2;
				 l_2 = -11; end
		2050: begin l_1 = +2;
				 l_2 = +12; end
		11791: begin l_1 = +2;
				 l_2 = -12; end
		2046: begin l_1 = -2;
				 l_2 = +12; end
		11787: begin l_1 = -2;
				 l_2 = -12; end
		4098: begin l_1 = +2;
				 l_2 = +13; end
		9743: begin l_1 = +2;
				 l_2 = -13; end
		4094: begin l_1 = -2;
				 l_2 = +13; end
		9739: begin l_1 = -2;
				 l_2 = -13; end
		8194: begin l_1 = +2;
				 l_2 = +14; end
		5647: begin l_1 = +2;
				 l_2 = -14; end
		8190: begin l_1 = -2;
				 l_2 = +14; end
		5643: begin l_1 = -2;
				 l_2 = -14; end
		2549: begin l_1 = +2;
				 l_2 = +15; end
		11292: begin l_1 = +2;
				 l_2 = -15; end
		2545: begin l_1 = -2;
				 l_2 = +15; end
		11288: begin l_1 = -2;
				 l_2 = -15; end
		5096: begin l_1 = +2;
				 l_2 = +16; end
		8745: begin l_1 = +2;
				 l_2 = -16; end
		5092: begin l_1 = -2;
				 l_2 = +16; end
		8741: begin l_1 = -2;
				 l_2 = -16; end
		10190: begin l_1 = +2;
				 l_2 = +17; end
		3651: begin l_1 = +2;
				 l_2 = -17; end
		10186: begin l_1 = -2;
				 l_2 = +17; end
		3647: begin l_1 = -2;
				 l_2 = -17; end
		6541: begin l_1 = +2;
				 l_2 = +18; end
		7300: begin l_1 = +2;
				 l_2 = -18; end
		6537: begin l_1 = -2;
				 l_2 = +18; end
		7296: begin l_1 = -2;
				 l_2 = -18; end
		13080: begin l_1 = +2;
				 l_2 = +19; end
		761: begin l_1 = +2;
				 l_2 = -19; end
		13076: begin l_1 = -2;
				 l_2 = +19; end
		757: begin l_1 = -2;
				 l_2 = -19; end
		12321: begin l_1 = +2;
				 l_2 = +20; end
		1520: begin l_1 = +2;
				 l_2 = -20; end
		12317: begin l_1 = -2;
				 l_2 = +20; end
		1516: begin l_1 = -2;
				 l_2 = -20; end
		10803: begin l_1 = +2;
				 l_2 = +21; end
		3038: begin l_1 = +2;
				 l_2 = -21; end
		10799: begin l_1 = -2;
				 l_2 = +21; end
		3034: begin l_1 = -2;
				 l_2 = -21; end
		7767: begin l_1 = +2;
				 l_2 = +22; end
		6074: begin l_1 = +2;
				 l_2 = -22; end
		7763: begin l_1 = -2;
				 l_2 = +22; end
		6070: begin l_1 = -2;
				 l_2 = -22; end
		1695: begin l_1 = +2;
				 l_2 = +23; end
		12146: begin l_1 = +2;
				 l_2 = -23; end
		1691: begin l_1 = -2;
				 l_2 = +23; end
		12142: begin l_1 = -2;
				 l_2 = -23; end
		3388: begin l_1 = +2;
				 l_2 = +24; end
		10453: begin l_1 = +2;
				 l_2 = -24; end
		3384: begin l_1 = -2;
				 l_2 = +24; end
		10449: begin l_1 = -2;
				 l_2 = -24; end
		6774: begin l_1 = +2;
				 l_2 = +25; end
		7067: begin l_1 = +2;
				 l_2 = -25; end
		6770: begin l_1 = -2;
				 l_2 = +25; end
		7063: begin l_1 = -2;
				 l_2 = -25; end
		13546: begin l_1 = +2;
				 l_2 = +26; end
		295: begin l_1 = +2;
				 l_2 = -26; end
		13542: begin l_1 = -2;
				 l_2 = +26; end
		291: begin l_1 = -2;
				 l_2 = -26; end
		13253: begin l_1 = +2;
				 l_2 = +27; end
		588: begin l_1 = +2;
				 l_2 = -27; end
		13249: begin l_1 = -2;
				 l_2 = +27; end
		584: begin l_1 = -2;
				 l_2 = -27; end
		12667: begin l_1 = +2;
				 l_2 = +28; end
		1174: begin l_1 = +2;
				 l_2 = -28; end
		12663: begin l_1 = -2;
				 l_2 = +28; end
		1170: begin l_1 = -2;
				 l_2 = -28; end
		11495: begin l_1 = +2;
				 l_2 = +29; end
		2346: begin l_1 = +2;
				 l_2 = -29; end
		11491: begin l_1 = -2;
				 l_2 = +29; end
		2342: begin l_1 = -2;
				 l_2 = -29; end
		9151: begin l_1 = +2;
				 l_2 = +30; end
		4690: begin l_1 = +2;
				 l_2 = -30; end
		9147: begin l_1 = -2;
				 l_2 = +30; end
		4686: begin l_1 = -2;
				 l_2 = -30; end
		4463: begin l_1 = +2;
				 l_2 = +31; end
		9378: begin l_1 = +2;
				 l_2 = -31; end
		4459: begin l_1 = -2;
				 l_2 = +31; end
		9374: begin l_1 = -2;
				 l_2 = -31; end
		8924: begin l_1 = +2;
				 l_2 = +32; end
		4917: begin l_1 = +2;
				 l_2 = -32; end
		8920: begin l_1 = -2;
				 l_2 = +32; end
		4913: begin l_1 = -2;
				 l_2 = -32; end
		4009: begin l_1 = +2;
				 l_2 = +33; end
		9832: begin l_1 = +2;
				 l_2 = -33; end
		4005: begin l_1 = -2;
				 l_2 = +33; end
		9828: begin l_1 = -2;
				 l_2 = -33; end
		8016: begin l_1 = +2;
				 l_2 = +34; end
		5825: begin l_1 = +2;
				 l_2 = -34; end
		8012: begin l_1 = -2;
				 l_2 = +34; end
		5821: begin l_1 = -2;
				 l_2 = -34; end
		2193: begin l_1 = +2;
				 l_2 = +35; end
		11648: begin l_1 = +2;
				 l_2 = -35; end
		2189: begin l_1 = -2;
				 l_2 = +35; end
		11644: begin l_1 = -2;
				 l_2 = -35; end
		4384: begin l_1 = +2;
				 l_2 = +36; end
		9457: begin l_1 = +2;
				 l_2 = -36; end
		4380: begin l_1 = -2;
				 l_2 = +36; end
		9453: begin l_1 = -2;
				 l_2 = -36; end
		8766: begin l_1 = +2;
				 l_2 = +37; end
		5075: begin l_1 = +2;
				 l_2 = -37; end
		8762: begin l_1 = -2;
				 l_2 = +37; end
		5071: begin l_1 = -2;
				 l_2 = -37; end
		3693: begin l_1 = +2;
				 l_2 = +38; end
		10148: begin l_1 = +2;
				 l_2 = -38; end
		3689: begin l_1 = -2;
				 l_2 = +38; end
		10144: begin l_1 = -2;
				 l_2 = -38; end
		12: begin l_1 = -3;
				 l_2 = +5; end
		13825: begin l_1 = -3;
				 l_2 = -4; end
		20: begin l_1 = +3;
				 l_2 = +5; end
		13817: begin l_1 = -3;
				 l_2 = -5; end
		36: begin l_1 = +3;
				 l_2 = +6; end
		13809: begin l_1 = +3;
				 l_2 = -6; end
		28: begin l_1 = -3;
				 l_2 = +6; end
		13801: begin l_1 = -3;
				 l_2 = -6; end
		68: begin l_1 = +3;
				 l_2 = +7; end
		13777: begin l_1 = +3;
				 l_2 = -7; end
		60: begin l_1 = -3;
				 l_2 = +7; end
		13769: begin l_1 = -3;
				 l_2 = -7; end
		132: begin l_1 = +3;
				 l_2 = +8; end
		13713: begin l_1 = +3;
				 l_2 = -8; end
		124: begin l_1 = -3;
				 l_2 = +8; end
		13705: begin l_1 = -3;
				 l_2 = -8; end
		260: begin l_1 = +3;
				 l_2 = +9; end
		13585: begin l_1 = +3;
				 l_2 = -9; end
		252: begin l_1 = -3;
				 l_2 = +9; end
		13577: begin l_1 = -3;
				 l_2 = -9; end
		516: begin l_1 = +3;
				 l_2 = +10; end
		13329: begin l_1 = +3;
				 l_2 = -10; end
		508: begin l_1 = -3;
				 l_2 = +10; end
		13321: begin l_1 = -3;
				 l_2 = -10; end
		1028: begin l_1 = +3;
				 l_2 = +11; end
		12817: begin l_1 = +3;
				 l_2 = -11; end
		1020: begin l_1 = -3;
				 l_2 = +11; end
		12809: begin l_1 = -3;
				 l_2 = -11; end
		2052: begin l_1 = +3;
				 l_2 = +12; end
		11793: begin l_1 = +3;
				 l_2 = -12; end
		2044: begin l_1 = -3;
				 l_2 = +12; end
		11785: begin l_1 = -3;
				 l_2 = -12; end
		4100: begin l_1 = +3;
				 l_2 = +13; end
		9745: begin l_1 = +3;
				 l_2 = -13; end
		4092: begin l_1 = -3;
				 l_2 = +13; end
		9737: begin l_1 = -3;
				 l_2 = -13; end
		8196: begin l_1 = +3;
				 l_2 = +14; end
		5649: begin l_1 = +3;
				 l_2 = -14; end
		8188: begin l_1 = -3;
				 l_2 = +14; end
		5641: begin l_1 = -3;
				 l_2 = -14; end
		2551: begin l_1 = +3;
				 l_2 = +15; end
		11294: begin l_1 = +3;
				 l_2 = -15; end
		2543: begin l_1 = -3;
				 l_2 = +15; end
		11286: begin l_1 = -3;
				 l_2 = -15; end
		5098: begin l_1 = +3;
				 l_2 = +16; end
		8747: begin l_1 = +3;
				 l_2 = -16; end
		5090: begin l_1 = -3;
				 l_2 = +16; end
		8739: begin l_1 = -3;
				 l_2 = -16; end
		10192: begin l_1 = +3;
				 l_2 = +17; end
		3653: begin l_1 = +3;
				 l_2 = -17; end
		10184: begin l_1 = -3;
				 l_2 = +17; end
		3645: begin l_1 = -3;
				 l_2 = -17; end
		6543: begin l_1 = +3;
				 l_2 = +18; end
		7302: begin l_1 = +3;
				 l_2 = -18; end
		6535: begin l_1 = -3;
				 l_2 = +18; end
		7294: begin l_1 = -3;
				 l_2 = -18; end
		13082: begin l_1 = +3;
				 l_2 = +19; end
		763: begin l_1 = +3;
				 l_2 = -19; end
		13074: begin l_1 = -3;
				 l_2 = +19; end
		755: begin l_1 = -3;
				 l_2 = -19; end
		12323: begin l_1 = +3;
				 l_2 = +20; end
		1522: begin l_1 = +3;
				 l_2 = -20; end
		12315: begin l_1 = -3;
				 l_2 = +20; end
		1514: begin l_1 = -3;
				 l_2 = -20; end
		10805: begin l_1 = +3;
				 l_2 = +21; end
		3040: begin l_1 = +3;
				 l_2 = -21; end
		10797: begin l_1 = -3;
				 l_2 = +21; end
		3032: begin l_1 = -3;
				 l_2 = -21; end
		7769: begin l_1 = +3;
				 l_2 = +22; end
		6076: begin l_1 = +3;
				 l_2 = -22; end
		7761: begin l_1 = -3;
				 l_2 = +22; end
		6068: begin l_1 = -3;
				 l_2 = -22; end
		1697: begin l_1 = +3;
				 l_2 = +23; end
		12148: begin l_1 = +3;
				 l_2 = -23; end
		1689: begin l_1 = -3;
				 l_2 = +23; end
		12140: begin l_1 = -3;
				 l_2 = -23; end
		3390: begin l_1 = +3;
				 l_2 = +24; end
		10455: begin l_1 = +3;
				 l_2 = -24; end
		3382: begin l_1 = -3;
				 l_2 = +24; end
		10447: begin l_1 = -3;
				 l_2 = -24; end
		6776: begin l_1 = +3;
				 l_2 = +25; end
		7069: begin l_1 = +3;
				 l_2 = -25; end
		6768: begin l_1 = -3;
				 l_2 = +25; end
		7061: begin l_1 = -3;
				 l_2 = -25; end
		13548: begin l_1 = +3;
				 l_2 = +26; end
		297: begin l_1 = +3;
				 l_2 = -26; end
		13540: begin l_1 = -3;
				 l_2 = +26; end
		289: begin l_1 = -3;
				 l_2 = -26; end
		13255: begin l_1 = +3;
				 l_2 = +27; end
		590: begin l_1 = +3;
				 l_2 = -27; end
		13247: begin l_1 = -3;
				 l_2 = +27; end
		582: begin l_1 = -3;
				 l_2 = -27; end
		12669: begin l_1 = +3;
				 l_2 = +28; end
		1176: begin l_1 = +3;
				 l_2 = -28; end
		12661: begin l_1 = -3;
				 l_2 = +28; end
		1168: begin l_1 = -3;
				 l_2 = -28; end
		11497: begin l_1 = +3;
				 l_2 = +29; end
		2348: begin l_1 = +3;
				 l_2 = -29; end
		11489: begin l_1 = -3;
				 l_2 = +29; end
		2340: begin l_1 = -3;
				 l_2 = -29; end
		9153: begin l_1 = +3;
				 l_2 = +30; end
		4692: begin l_1 = +3;
				 l_2 = -30; end
		9145: begin l_1 = -3;
				 l_2 = +30; end
		4684: begin l_1 = -3;
				 l_2 = -30; end
		4465: begin l_1 = +3;
				 l_2 = +31; end
		9380: begin l_1 = +3;
				 l_2 = -31; end
		4457: begin l_1 = -3;
				 l_2 = +31; end
		9372: begin l_1 = -3;
				 l_2 = -31; end
		8926: begin l_1 = +3;
				 l_2 = +32; end
		4919: begin l_1 = +3;
				 l_2 = -32; end
		8918: begin l_1 = -3;
				 l_2 = +32; end
		4911: begin l_1 = -3;
				 l_2 = -32; end
		4011: begin l_1 = +3;
				 l_2 = +33; end
		9834: begin l_1 = +3;
				 l_2 = -33; end
		4003: begin l_1 = -3;
				 l_2 = +33; end
		9826: begin l_1 = -3;
				 l_2 = -33; end
		8018: begin l_1 = +3;
				 l_2 = +34; end
		5827: begin l_1 = +3;
				 l_2 = -34; end
		8010: begin l_1 = -3;
				 l_2 = +34; end
		5819: begin l_1 = -3;
				 l_2 = -34; end
		2195: begin l_1 = +3;
				 l_2 = +35; end
		11650: begin l_1 = +3;
				 l_2 = -35; end
		2187: begin l_1 = -3;
				 l_2 = +35; end
		11642: begin l_1 = -3;
				 l_2 = -35; end
		4386: begin l_1 = +3;
				 l_2 = +36; end
		9459: begin l_1 = +3;
				 l_2 = -36; end
		4378: begin l_1 = -3;
				 l_2 = +36; end
		9451: begin l_1 = -3;
				 l_2 = -36; end
		8768: begin l_1 = +3;
				 l_2 = +37; end
		5077: begin l_1 = +3;
				 l_2 = -37; end
		8760: begin l_1 = -3;
				 l_2 = +37; end
		5069: begin l_1 = -3;
				 l_2 = -37; end
		3695: begin l_1 = +3;
				 l_2 = +38; end
		10150: begin l_1 = +3;
				 l_2 = -38; end
		3687: begin l_1 = -3;
				 l_2 = +38; end
		10142: begin l_1 = -3;
				 l_2 = -38; end
		24: begin l_1 = -4;
				 l_2 = +6; end
		13813: begin l_1 = -4;
				 l_2 = -5; end
		40: begin l_1 = +4;
				 l_2 = +6; end
		13797: begin l_1 = -4;
				 l_2 = -6; end
		72: begin l_1 = +4;
				 l_2 = +7; end
		13781: begin l_1 = +4;
				 l_2 = -7; end
		56: begin l_1 = -4;
				 l_2 = +7; end
		13765: begin l_1 = -4;
				 l_2 = -7; end
		136: begin l_1 = +4;
				 l_2 = +8; end
		13717: begin l_1 = +4;
				 l_2 = -8; end
		120: begin l_1 = -4;
				 l_2 = +8; end
		13701: begin l_1 = -4;
				 l_2 = -8; end
		264: begin l_1 = +4;
				 l_2 = +9; end
		13589: begin l_1 = +4;
				 l_2 = -9; end
		248: begin l_1 = -4;
				 l_2 = +9; end
		13573: begin l_1 = -4;
				 l_2 = -9; end
		520: begin l_1 = +4;
				 l_2 = +10; end
		13333: begin l_1 = +4;
				 l_2 = -10; end
		504: begin l_1 = -4;
				 l_2 = +10; end
		13317: begin l_1 = -4;
				 l_2 = -10; end
		1032: begin l_1 = +4;
				 l_2 = +11; end
		12821: begin l_1 = +4;
				 l_2 = -11; end
		1016: begin l_1 = -4;
				 l_2 = +11; end
		12805: begin l_1 = -4;
				 l_2 = -11; end
		2056: begin l_1 = +4;
				 l_2 = +12; end
		11797: begin l_1 = +4;
				 l_2 = -12; end
		2040: begin l_1 = -4;
				 l_2 = +12; end
		11781: begin l_1 = -4;
				 l_2 = -12; end
		4104: begin l_1 = +4;
				 l_2 = +13; end
		9749: begin l_1 = +4;
				 l_2 = -13; end
		4088: begin l_1 = -4;
				 l_2 = +13; end
		9733: begin l_1 = -4;
				 l_2 = -13; end
		8200: begin l_1 = +4;
				 l_2 = +14; end
		5653: begin l_1 = +4;
				 l_2 = -14; end
		8184: begin l_1 = -4;
				 l_2 = +14; end
		5637: begin l_1 = -4;
				 l_2 = -14; end
		2555: begin l_1 = +4;
				 l_2 = +15; end
		11298: begin l_1 = +4;
				 l_2 = -15; end
		2539: begin l_1 = -4;
				 l_2 = +15; end
		11282: begin l_1 = -4;
				 l_2 = -15; end
		5102: begin l_1 = +4;
				 l_2 = +16; end
		8751: begin l_1 = +4;
				 l_2 = -16; end
		5086: begin l_1 = -4;
				 l_2 = +16; end
		8735: begin l_1 = -4;
				 l_2 = -16; end
		10196: begin l_1 = +4;
				 l_2 = +17; end
		3657: begin l_1 = +4;
				 l_2 = -17; end
		10180: begin l_1 = -4;
				 l_2 = +17; end
		3641: begin l_1 = -4;
				 l_2 = -17; end
		6547: begin l_1 = +4;
				 l_2 = +18; end
		7306: begin l_1 = +4;
				 l_2 = -18; end
		6531: begin l_1 = -4;
				 l_2 = +18; end
		7290: begin l_1 = -4;
				 l_2 = -18; end
		13086: begin l_1 = +4;
				 l_2 = +19; end
		767: begin l_1 = +4;
				 l_2 = -19; end
		13070: begin l_1 = -4;
				 l_2 = +19; end
		751: begin l_1 = -4;
				 l_2 = -19; end
		12327: begin l_1 = +4;
				 l_2 = +20; end
		1526: begin l_1 = +4;
				 l_2 = -20; end
		12311: begin l_1 = -4;
				 l_2 = +20; end
		1510: begin l_1 = -4;
				 l_2 = -20; end
		10809: begin l_1 = +4;
				 l_2 = +21; end
		3044: begin l_1 = +4;
				 l_2 = -21; end
		10793: begin l_1 = -4;
				 l_2 = +21; end
		3028: begin l_1 = -4;
				 l_2 = -21; end
		7773: begin l_1 = +4;
				 l_2 = +22; end
		6080: begin l_1 = +4;
				 l_2 = -22; end
		7757: begin l_1 = -4;
				 l_2 = +22; end
		6064: begin l_1 = -4;
				 l_2 = -22; end
		1701: begin l_1 = +4;
				 l_2 = +23; end
		12152: begin l_1 = +4;
				 l_2 = -23; end
		1685: begin l_1 = -4;
				 l_2 = +23; end
		12136: begin l_1 = -4;
				 l_2 = -23; end
		3394: begin l_1 = +4;
				 l_2 = +24; end
		10459: begin l_1 = +4;
				 l_2 = -24; end
		3378: begin l_1 = -4;
				 l_2 = +24; end
		10443: begin l_1 = -4;
				 l_2 = -24; end
		6780: begin l_1 = +4;
				 l_2 = +25; end
		7073: begin l_1 = +4;
				 l_2 = -25; end
		6764: begin l_1 = -4;
				 l_2 = +25; end
		7057: begin l_1 = -4;
				 l_2 = -25; end
		13552: begin l_1 = +4;
				 l_2 = +26; end
		301: begin l_1 = +4;
				 l_2 = -26; end
		13536: begin l_1 = -4;
				 l_2 = +26; end
		285: begin l_1 = -4;
				 l_2 = -26; end
		13259: begin l_1 = +4;
				 l_2 = +27; end
		594: begin l_1 = +4;
				 l_2 = -27; end
		13243: begin l_1 = -4;
				 l_2 = +27; end
		578: begin l_1 = -4;
				 l_2 = -27; end
		12673: begin l_1 = +4;
				 l_2 = +28; end
		1180: begin l_1 = +4;
				 l_2 = -28; end
		12657: begin l_1 = -4;
				 l_2 = +28; end
		1164: begin l_1 = -4;
				 l_2 = -28; end
		11501: begin l_1 = +4;
				 l_2 = +29; end
		2352: begin l_1 = +4;
				 l_2 = -29; end
		11485: begin l_1 = -4;
				 l_2 = +29; end
		2336: begin l_1 = -4;
				 l_2 = -29; end
		9157: begin l_1 = +4;
				 l_2 = +30; end
		4696: begin l_1 = +4;
				 l_2 = -30; end
		9141: begin l_1 = -4;
				 l_2 = +30; end
		4680: begin l_1 = -4;
				 l_2 = -30; end
		4469: begin l_1 = +4;
				 l_2 = +31; end
		9384: begin l_1 = +4;
				 l_2 = -31; end
		4453: begin l_1 = -4;
				 l_2 = +31; end
		9368: begin l_1 = -4;
				 l_2 = -31; end
		8930: begin l_1 = +4;
				 l_2 = +32; end
		4923: begin l_1 = +4;
				 l_2 = -32; end
		8914: begin l_1 = -4;
				 l_2 = +32; end
		4907: begin l_1 = -4;
				 l_2 = -32; end
		4015: begin l_1 = +4;
				 l_2 = +33; end
		9838: begin l_1 = +4;
				 l_2 = -33; end
		3999: begin l_1 = -4;
				 l_2 = +33; end
		9822: begin l_1 = -4;
				 l_2 = -33; end
		8022: begin l_1 = +4;
				 l_2 = +34; end
		5831: begin l_1 = +4;
				 l_2 = -34; end
		8006: begin l_1 = -4;
				 l_2 = +34; end
		5815: begin l_1 = -4;
				 l_2 = -34; end
		2199: begin l_1 = +4;
				 l_2 = +35; end
		11654: begin l_1 = +4;
				 l_2 = -35; end
		2183: begin l_1 = -4;
				 l_2 = +35; end
		11638: begin l_1 = -4;
				 l_2 = -35; end
		4390: begin l_1 = +4;
				 l_2 = +36; end
		9463: begin l_1 = +4;
				 l_2 = -36; end
		4374: begin l_1 = -4;
				 l_2 = +36; end
		9447: begin l_1 = -4;
				 l_2 = -36; end
		8772: begin l_1 = +4;
				 l_2 = +37; end
		5081: begin l_1 = +4;
				 l_2 = -37; end
		8756: begin l_1 = -4;
				 l_2 = +37; end
		5065: begin l_1 = -4;
				 l_2 = -37; end
		3699: begin l_1 = +4;
				 l_2 = +38; end
		10154: begin l_1 = +4;
				 l_2 = -38; end
		3683: begin l_1 = -4;
				 l_2 = +38; end
		10138: begin l_1 = -4;
				 l_2 = -38; end
		48: begin l_1 = -5;
				 l_2 = +7; end
		13789: begin l_1 = -5;
				 l_2 = -6; end
		80: begin l_1 = +5;
				 l_2 = +7; end
		13757: begin l_1 = -5;
				 l_2 = -7; end
		144: begin l_1 = +5;
				 l_2 = +8; end
		13725: begin l_1 = +5;
				 l_2 = -8; end
		112: begin l_1 = -5;
				 l_2 = +8; end
		13693: begin l_1 = -5;
				 l_2 = -8; end
		272: begin l_1 = +5;
				 l_2 = +9; end
		13597: begin l_1 = +5;
				 l_2 = -9; end
		240: begin l_1 = -5;
				 l_2 = +9; end
		13565: begin l_1 = -5;
				 l_2 = -9; end
		528: begin l_1 = +5;
				 l_2 = +10; end
		13341: begin l_1 = +5;
				 l_2 = -10; end
		496: begin l_1 = -5;
				 l_2 = +10; end
		13309: begin l_1 = -5;
				 l_2 = -10; end
		1040: begin l_1 = +5;
				 l_2 = +11; end
		12829: begin l_1 = +5;
				 l_2 = -11; end
		1008: begin l_1 = -5;
				 l_2 = +11; end
		12797: begin l_1 = -5;
				 l_2 = -11; end
		2064: begin l_1 = +5;
				 l_2 = +12; end
		11805: begin l_1 = +5;
				 l_2 = -12; end
		2032: begin l_1 = -5;
				 l_2 = +12; end
		11773: begin l_1 = -5;
				 l_2 = -12; end
		4112: begin l_1 = +5;
				 l_2 = +13; end
		9757: begin l_1 = +5;
				 l_2 = -13; end
		4080: begin l_1 = -5;
				 l_2 = +13; end
		9725: begin l_1 = -5;
				 l_2 = -13; end
		8208: begin l_1 = +5;
				 l_2 = +14; end
		5661: begin l_1 = +5;
				 l_2 = -14; end
		8176: begin l_1 = -5;
				 l_2 = +14; end
		5629: begin l_1 = -5;
				 l_2 = -14; end
		2563: begin l_1 = +5;
				 l_2 = +15; end
		11306: begin l_1 = +5;
				 l_2 = -15; end
		2531: begin l_1 = -5;
				 l_2 = +15; end
		11274: begin l_1 = -5;
				 l_2 = -15; end
		5110: begin l_1 = +5;
				 l_2 = +16; end
		8759: begin l_1 = +5;
				 l_2 = -16; end
		5078: begin l_1 = -5;
				 l_2 = +16; end
		8727: begin l_1 = -5;
				 l_2 = -16; end
		10204: begin l_1 = +5;
				 l_2 = +17; end
		3665: begin l_1 = +5;
				 l_2 = -17; end
		10172: begin l_1 = -5;
				 l_2 = +17; end
		3633: begin l_1 = -5;
				 l_2 = -17; end
		6555: begin l_1 = +5;
				 l_2 = +18; end
		7314: begin l_1 = +5;
				 l_2 = -18; end
		6523: begin l_1 = -5;
				 l_2 = +18; end
		7282: begin l_1 = -5;
				 l_2 = -18; end
		13094: begin l_1 = +5;
				 l_2 = +19; end
		775: begin l_1 = +5;
				 l_2 = -19; end
		13062: begin l_1 = -5;
				 l_2 = +19; end
		743: begin l_1 = -5;
				 l_2 = -19; end
		12335: begin l_1 = +5;
				 l_2 = +20; end
		1534: begin l_1 = +5;
				 l_2 = -20; end
		12303: begin l_1 = -5;
				 l_2 = +20; end
		1502: begin l_1 = -5;
				 l_2 = -20; end
		10817: begin l_1 = +5;
				 l_2 = +21; end
		3052: begin l_1 = +5;
				 l_2 = -21; end
		10785: begin l_1 = -5;
				 l_2 = +21; end
		3020: begin l_1 = -5;
				 l_2 = -21; end
		7781: begin l_1 = +5;
				 l_2 = +22; end
		6088: begin l_1 = +5;
				 l_2 = -22; end
		7749: begin l_1 = -5;
				 l_2 = +22; end
		6056: begin l_1 = -5;
				 l_2 = -22; end
		1709: begin l_1 = +5;
				 l_2 = +23; end
		12160: begin l_1 = +5;
				 l_2 = -23; end
		1677: begin l_1 = -5;
				 l_2 = +23; end
		12128: begin l_1 = -5;
				 l_2 = -23; end
		3402: begin l_1 = +5;
				 l_2 = +24; end
		10467: begin l_1 = +5;
				 l_2 = -24; end
		3370: begin l_1 = -5;
				 l_2 = +24; end
		10435: begin l_1 = -5;
				 l_2 = -24; end
		6788: begin l_1 = +5;
				 l_2 = +25; end
		7081: begin l_1 = +5;
				 l_2 = -25; end
		6756: begin l_1 = -5;
				 l_2 = +25; end
		7049: begin l_1 = -5;
				 l_2 = -25; end
		13560: begin l_1 = +5;
				 l_2 = +26; end
		309: begin l_1 = +5;
				 l_2 = -26; end
		13528: begin l_1 = -5;
				 l_2 = +26; end
		277: begin l_1 = -5;
				 l_2 = -26; end
		13267: begin l_1 = +5;
				 l_2 = +27; end
		602: begin l_1 = +5;
				 l_2 = -27; end
		13235: begin l_1 = -5;
				 l_2 = +27; end
		570: begin l_1 = -5;
				 l_2 = -27; end
		12681: begin l_1 = +5;
				 l_2 = +28; end
		1188: begin l_1 = +5;
				 l_2 = -28; end
		12649: begin l_1 = -5;
				 l_2 = +28; end
		1156: begin l_1 = -5;
				 l_2 = -28; end
		11509: begin l_1 = +5;
				 l_2 = +29; end
		2360: begin l_1 = +5;
				 l_2 = -29; end
		11477: begin l_1 = -5;
				 l_2 = +29; end
		2328: begin l_1 = -5;
				 l_2 = -29; end
		9165: begin l_1 = +5;
				 l_2 = +30; end
		4704: begin l_1 = +5;
				 l_2 = -30; end
		9133: begin l_1 = -5;
				 l_2 = +30; end
		4672: begin l_1 = -5;
				 l_2 = -30; end
		4477: begin l_1 = +5;
				 l_2 = +31; end
		9392: begin l_1 = +5;
				 l_2 = -31; end
		4445: begin l_1 = -5;
				 l_2 = +31; end
		9360: begin l_1 = -5;
				 l_2 = -31; end
		8938: begin l_1 = +5;
				 l_2 = +32; end
		4931: begin l_1 = +5;
				 l_2 = -32; end
		8906: begin l_1 = -5;
				 l_2 = +32; end
		4899: begin l_1 = -5;
				 l_2 = -32; end
		4023: begin l_1 = +5;
				 l_2 = +33; end
		9846: begin l_1 = +5;
				 l_2 = -33; end
		3991: begin l_1 = -5;
				 l_2 = +33; end
		9814: begin l_1 = -5;
				 l_2 = -33; end
		8030: begin l_1 = +5;
				 l_2 = +34; end
		5839: begin l_1 = +5;
				 l_2 = -34; end
		7998: begin l_1 = -5;
				 l_2 = +34; end
		5807: begin l_1 = -5;
				 l_2 = -34; end
		2207: begin l_1 = +5;
				 l_2 = +35; end
		11662: begin l_1 = +5;
				 l_2 = -35; end
		2175: begin l_1 = -5;
				 l_2 = +35; end
		11630: begin l_1 = -5;
				 l_2 = -35; end
		4398: begin l_1 = +5;
				 l_2 = +36; end
		9471: begin l_1 = +5;
				 l_2 = -36; end
		4366: begin l_1 = -5;
				 l_2 = +36; end
		9439: begin l_1 = -5;
				 l_2 = -36; end
		8780: begin l_1 = +5;
				 l_2 = +37; end
		5089: begin l_1 = +5;
				 l_2 = -37; end
		8748: begin l_1 = -5;
				 l_2 = +37; end
		5057: begin l_1 = -5;
				 l_2 = -37; end
		3707: begin l_1 = +5;
				 l_2 = +38; end
		10162: begin l_1 = +5;
				 l_2 = -38; end
		3675: begin l_1 = -5;
				 l_2 = +38; end
		10130: begin l_1 = -5;
				 l_2 = -38; end
		96: begin l_1 = -6;
				 l_2 = +8; end
		13741: begin l_1 = -6;
				 l_2 = -7; end
		160: begin l_1 = +6;
				 l_2 = +8; end
		13677: begin l_1 = -6;
				 l_2 = -8; end
		288: begin l_1 = +6;
				 l_2 = +9; end
		13613: begin l_1 = +6;
				 l_2 = -9; end
		224: begin l_1 = -6;
				 l_2 = +9; end
		13549: begin l_1 = -6;
				 l_2 = -9; end
		544: begin l_1 = +6;
				 l_2 = +10; end
		13357: begin l_1 = +6;
				 l_2 = -10; end
		480: begin l_1 = -6;
				 l_2 = +10; end
		13293: begin l_1 = -6;
				 l_2 = -10; end
		1056: begin l_1 = +6;
				 l_2 = +11; end
		12845: begin l_1 = +6;
				 l_2 = -11; end
		992: begin l_1 = -6;
				 l_2 = +11; end
		12781: begin l_1 = -6;
				 l_2 = -11; end
		2080: begin l_1 = +6;
				 l_2 = +12; end
		11821: begin l_1 = +6;
				 l_2 = -12; end
		2016: begin l_1 = -6;
				 l_2 = +12; end
		11757: begin l_1 = -6;
				 l_2 = -12; end
		4128: begin l_1 = +6;
				 l_2 = +13; end
		9773: begin l_1 = +6;
				 l_2 = -13; end
		4064: begin l_1 = -6;
				 l_2 = +13; end
		9709: begin l_1 = -6;
				 l_2 = -13; end
		8224: begin l_1 = +6;
				 l_2 = +14; end
		5677: begin l_1 = +6;
				 l_2 = -14; end
		8160: begin l_1 = -6;
				 l_2 = +14; end
		5613: begin l_1 = -6;
				 l_2 = -14; end
		2579: begin l_1 = +6;
				 l_2 = +15; end
		11322: begin l_1 = +6;
				 l_2 = -15; end
		2515: begin l_1 = -6;
				 l_2 = +15; end
		11258: begin l_1 = -6;
				 l_2 = -15; end
		5126: begin l_1 = +6;
				 l_2 = +16; end
		8775: begin l_1 = +6;
				 l_2 = -16; end
		5062: begin l_1 = -6;
				 l_2 = +16; end
		8711: begin l_1 = -6;
				 l_2 = -16; end
		10220: begin l_1 = +6;
				 l_2 = +17; end
		3681: begin l_1 = +6;
				 l_2 = -17; end
		10156: begin l_1 = -6;
				 l_2 = +17; end
		3617: begin l_1 = -6;
				 l_2 = -17; end
		6571: begin l_1 = +6;
				 l_2 = +18; end
		7330: begin l_1 = +6;
				 l_2 = -18; end
		6507: begin l_1 = -6;
				 l_2 = +18; end
		7266: begin l_1 = -6;
				 l_2 = -18; end
		13110: begin l_1 = +6;
				 l_2 = +19; end
		791: begin l_1 = +6;
				 l_2 = -19; end
		13046: begin l_1 = -6;
				 l_2 = +19; end
		727: begin l_1 = -6;
				 l_2 = -19; end
		12351: begin l_1 = +6;
				 l_2 = +20; end
		1550: begin l_1 = +6;
				 l_2 = -20; end
		12287: begin l_1 = -6;
				 l_2 = +20; end
		1486: begin l_1 = -6;
				 l_2 = -20; end
		10833: begin l_1 = +6;
				 l_2 = +21; end
		3068: begin l_1 = +6;
				 l_2 = -21; end
		10769: begin l_1 = -6;
				 l_2 = +21; end
		3004: begin l_1 = -6;
				 l_2 = -21; end
		7797: begin l_1 = +6;
				 l_2 = +22; end
		6104: begin l_1 = +6;
				 l_2 = -22; end
		7733: begin l_1 = -6;
				 l_2 = +22; end
		6040: begin l_1 = -6;
				 l_2 = -22; end
		1725: begin l_1 = +6;
				 l_2 = +23; end
		12176: begin l_1 = +6;
				 l_2 = -23; end
		1661: begin l_1 = -6;
				 l_2 = +23; end
		12112: begin l_1 = -6;
				 l_2 = -23; end
		3418: begin l_1 = +6;
				 l_2 = +24; end
		10483: begin l_1 = +6;
				 l_2 = -24; end
		3354: begin l_1 = -6;
				 l_2 = +24; end
		10419: begin l_1 = -6;
				 l_2 = -24; end
		6804: begin l_1 = +6;
				 l_2 = +25; end
		7097: begin l_1 = +6;
				 l_2 = -25; end
		6740: begin l_1 = -6;
				 l_2 = +25; end
		7033: begin l_1 = -6;
				 l_2 = -25; end
		13576: begin l_1 = +6;
				 l_2 = +26; end
		325: begin l_1 = +6;
				 l_2 = -26; end
		13512: begin l_1 = -6;
				 l_2 = +26; end
		261: begin l_1 = -6;
				 l_2 = -26; end
		13283: begin l_1 = +6;
				 l_2 = +27; end
		618: begin l_1 = +6;
				 l_2 = -27; end
		13219: begin l_1 = -6;
				 l_2 = +27; end
		554: begin l_1 = -6;
				 l_2 = -27; end
		12697: begin l_1 = +6;
				 l_2 = +28; end
		1204: begin l_1 = +6;
				 l_2 = -28; end
		12633: begin l_1 = -6;
				 l_2 = +28; end
		1140: begin l_1 = -6;
				 l_2 = -28; end
		11525: begin l_1 = +6;
				 l_2 = +29; end
		2376: begin l_1 = +6;
				 l_2 = -29; end
		11461: begin l_1 = -6;
				 l_2 = +29; end
		2312: begin l_1 = -6;
				 l_2 = -29; end
		9181: begin l_1 = +6;
				 l_2 = +30; end
		4720: begin l_1 = +6;
				 l_2 = -30; end
		9117: begin l_1 = -6;
				 l_2 = +30; end
		4656: begin l_1 = -6;
				 l_2 = -30; end
		4493: begin l_1 = +6;
				 l_2 = +31; end
		9408: begin l_1 = +6;
				 l_2 = -31; end
		4429: begin l_1 = -6;
				 l_2 = +31; end
		9344: begin l_1 = -6;
				 l_2 = -31; end
		8954: begin l_1 = +6;
				 l_2 = +32; end
		4947: begin l_1 = +6;
				 l_2 = -32; end
		8890: begin l_1 = -6;
				 l_2 = +32; end
		4883: begin l_1 = -6;
				 l_2 = -32; end
		4039: begin l_1 = +6;
				 l_2 = +33; end
		9862: begin l_1 = +6;
				 l_2 = -33; end
		3975: begin l_1 = -6;
				 l_2 = +33; end
		9798: begin l_1 = -6;
				 l_2 = -33; end
		8046: begin l_1 = +6;
				 l_2 = +34; end
		5855: begin l_1 = +6;
				 l_2 = -34; end
		7982: begin l_1 = -6;
				 l_2 = +34; end
		5791: begin l_1 = -6;
				 l_2 = -34; end
		2223: begin l_1 = +6;
				 l_2 = +35; end
		11678: begin l_1 = +6;
				 l_2 = -35; end
		2159: begin l_1 = -6;
				 l_2 = +35; end
		11614: begin l_1 = -6;
				 l_2 = -35; end
		4414: begin l_1 = +6;
				 l_2 = +36; end
		9487: begin l_1 = +6;
				 l_2 = -36; end
		4350: begin l_1 = -6;
				 l_2 = +36; end
		9423: begin l_1 = -6;
				 l_2 = -36; end
		8796: begin l_1 = +6;
				 l_2 = +37; end
		5105: begin l_1 = +6;
				 l_2 = -37; end
		8732: begin l_1 = -6;
				 l_2 = +37; end
		5041: begin l_1 = -6;
				 l_2 = -37; end
		3723: begin l_1 = +6;
				 l_2 = +38; end
		10178: begin l_1 = +6;
				 l_2 = -38; end
		3659: begin l_1 = -6;
				 l_2 = +38; end
		10114: begin l_1 = -6;
				 l_2 = -38; end
		192: begin l_1 = -7;
				 l_2 = +9; end
		13645: begin l_1 = -7;
				 l_2 = -8; end
		320: begin l_1 = +7;
				 l_2 = +9; end
		13517: begin l_1 = -7;
				 l_2 = -9; end
		576: begin l_1 = +7;
				 l_2 = +10; end
		13389: begin l_1 = +7;
				 l_2 = -10; end
		448: begin l_1 = -7;
				 l_2 = +10; end
		13261: begin l_1 = -7;
				 l_2 = -10; end
		1088: begin l_1 = +7;
				 l_2 = +11; end
		12877: begin l_1 = +7;
				 l_2 = -11; end
		960: begin l_1 = -7;
				 l_2 = +11; end
		12749: begin l_1 = -7;
				 l_2 = -11; end
		2112: begin l_1 = +7;
				 l_2 = +12; end
		11853: begin l_1 = +7;
				 l_2 = -12; end
		1984: begin l_1 = -7;
				 l_2 = +12; end
		11725: begin l_1 = -7;
				 l_2 = -12; end
		4160: begin l_1 = +7;
				 l_2 = +13; end
		9805: begin l_1 = +7;
				 l_2 = -13; end
		4032: begin l_1 = -7;
				 l_2 = +13; end
		9677: begin l_1 = -7;
				 l_2 = -13; end
		8256: begin l_1 = +7;
				 l_2 = +14; end
		5709: begin l_1 = +7;
				 l_2 = -14; end
		8128: begin l_1 = -7;
				 l_2 = +14; end
		5581: begin l_1 = -7;
				 l_2 = -14; end
		2611: begin l_1 = +7;
				 l_2 = +15; end
		11354: begin l_1 = +7;
				 l_2 = -15; end
		2483: begin l_1 = -7;
				 l_2 = +15; end
		11226: begin l_1 = -7;
				 l_2 = -15; end
		5158: begin l_1 = +7;
				 l_2 = +16; end
		8807: begin l_1 = +7;
				 l_2 = -16; end
		5030: begin l_1 = -7;
				 l_2 = +16; end
		8679: begin l_1 = -7;
				 l_2 = -16; end
		10252: begin l_1 = +7;
				 l_2 = +17; end
		3713: begin l_1 = +7;
				 l_2 = -17; end
		10124: begin l_1 = -7;
				 l_2 = +17; end
		3585: begin l_1 = -7;
				 l_2 = -17; end
		6603: begin l_1 = +7;
				 l_2 = +18; end
		7362: begin l_1 = +7;
				 l_2 = -18; end
		6475: begin l_1 = -7;
				 l_2 = +18; end
		7234: begin l_1 = -7;
				 l_2 = -18; end
		13142: begin l_1 = +7;
				 l_2 = +19; end
		823: begin l_1 = +7;
				 l_2 = -19; end
		13014: begin l_1 = -7;
				 l_2 = +19; end
		695: begin l_1 = -7;
				 l_2 = -19; end
		12383: begin l_1 = +7;
				 l_2 = +20; end
		1582: begin l_1 = +7;
				 l_2 = -20; end
		12255: begin l_1 = -7;
				 l_2 = +20; end
		1454: begin l_1 = -7;
				 l_2 = -20; end
		10865: begin l_1 = +7;
				 l_2 = +21; end
		3100: begin l_1 = +7;
				 l_2 = -21; end
		10737: begin l_1 = -7;
				 l_2 = +21; end
		2972: begin l_1 = -7;
				 l_2 = -21; end
		7829: begin l_1 = +7;
				 l_2 = +22; end
		6136: begin l_1 = +7;
				 l_2 = -22; end
		7701: begin l_1 = -7;
				 l_2 = +22; end
		6008: begin l_1 = -7;
				 l_2 = -22; end
		1757: begin l_1 = +7;
				 l_2 = +23; end
		12208: begin l_1 = +7;
				 l_2 = -23; end
		1629: begin l_1 = -7;
				 l_2 = +23; end
		12080: begin l_1 = -7;
				 l_2 = -23; end
		3450: begin l_1 = +7;
				 l_2 = +24; end
		10515: begin l_1 = +7;
				 l_2 = -24; end
		3322: begin l_1 = -7;
				 l_2 = +24; end
		10387: begin l_1 = -7;
				 l_2 = -24; end
		6836: begin l_1 = +7;
				 l_2 = +25; end
		7129: begin l_1 = +7;
				 l_2 = -25; end
		6708: begin l_1 = -7;
				 l_2 = +25; end
		7001: begin l_1 = -7;
				 l_2 = -25; end
		13608: begin l_1 = +7;
				 l_2 = +26; end
		357: begin l_1 = +7;
				 l_2 = -26; end
		13480: begin l_1 = -7;
				 l_2 = +26; end
		229: begin l_1 = -7;
				 l_2 = -26; end
		13315: begin l_1 = +7;
				 l_2 = +27; end
		650: begin l_1 = +7;
				 l_2 = -27; end
		13187: begin l_1 = -7;
				 l_2 = +27; end
		522: begin l_1 = -7;
				 l_2 = -27; end
		12729: begin l_1 = +7;
				 l_2 = +28; end
		1236: begin l_1 = +7;
				 l_2 = -28; end
		12601: begin l_1 = -7;
				 l_2 = +28; end
		1108: begin l_1 = -7;
				 l_2 = -28; end
		11557: begin l_1 = +7;
				 l_2 = +29; end
		2408: begin l_1 = +7;
				 l_2 = -29; end
		11429: begin l_1 = -7;
				 l_2 = +29; end
		2280: begin l_1 = -7;
				 l_2 = -29; end
		9213: begin l_1 = +7;
				 l_2 = +30; end
		4752: begin l_1 = +7;
				 l_2 = -30; end
		9085: begin l_1 = -7;
				 l_2 = +30; end
		4624: begin l_1 = -7;
				 l_2 = -30; end
		4525: begin l_1 = +7;
				 l_2 = +31; end
		9440: begin l_1 = +7;
				 l_2 = -31; end
		4397: begin l_1 = -7;
				 l_2 = +31; end
		9312: begin l_1 = -7;
				 l_2 = -31; end
		8986: begin l_1 = +7;
				 l_2 = +32; end
		4979: begin l_1 = +7;
				 l_2 = -32; end
		8858: begin l_1 = -7;
				 l_2 = +32; end
		4851: begin l_1 = -7;
				 l_2 = -32; end
		4071: begin l_1 = +7;
				 l_2 = +33; end
		9894: begin l_1 = +7;
				 l_2 = -33; end
		3943: begin l_1 = -7;
				 l_2 = +33; end
		9766: begin l_1 = -7;
				 l_2 = -33; end
		8078: begin l_1 = +7;
				 l_2 = +34; end
		5887: begin l_1 = +7;
				 l_2 = -34; end
		7950: begin l_1 = -7;
				 l_2 = +34; end
		5759: begin l_1 = -7;
				 l_2 = -34; end
		2255: begin l_1 = +7;
				 l_2 = +35; end
		11710: begin l_1 = +7;
				 l_2 = -35; end
		2127: begin l_1 = -7;
				 l_2 = +35; end
		11582: begin l_1 = -7;
				 l_2 = -35; end
		4446: begin l_1 = +7;
				 l_2 = +36; end
		9519: begin l_1 = +7;
				 l_2 = -36; end
		4318: begin l_1 = -7;
				 l_2 = +36; end
		9391: begin l_1 = -7;
				 l_2 = -36; end
		8828: begin l_1 = +7;
				 l_2 = +37; end
		5137: begin l_1 = +7;
				 l_2 = -37; end
		8700: begin l_1 = -7;
				 l_2 = +37; end
		5009: begin l_1 = -7;
				 l_2 = -37; end
		3755: begin l_1 = +7;
				 l_2 = +38; end
		10210: begin l_1 = +7;
				 l_2 = -38; end
		3627: begin l_1 = -7;
				 l_2 = +38; end
		10082: begin l_1 = -7;
				 l_2 = -38; end
		384: begin l_1 = -8;
				 l_2 = +10; end
		13453: begin l_1 = -8;
				 l_2 = -9; end
		640: begin l_1 = +8;
				 l_2 = +10; end
		13197: begin l_1 = -8;
				 l_2 = -10; end
		1152: begin l_1 = +8;
				 l_2 = +11; end
		12941: begin l_1 = +8;
				 l_2 = -11; end
		896: begin l_1 = -8;
				 l_2 = +11; end
		12685: begin l_1 = -8;
				 l_2 = -11; end
		2176: begin l_1 = +8;
				 l_2 = +12; end
		11917: begin l_1 = +8;
				 l_2 = -12; end
		1920: begin l_1 = -8;
				 l_2 = +12; end
		11661: begin l_1 = -8;
				 l_2 = -12; end
		4224: begin l_1 = +8;
				 l_2 = +13; end
		9869: begin l_1 = +8;
				 l_2 = -13; end
		3968: begin l_1 = -8;
				 l_2 = +13; end
		9613: begin l_1 = -8;
				 l_2 = -13; end
		8320: begin l_1 = +8;
				 l_2 = +14; end
		5773: begin l_1 = +8;
				 l_2 = -14; end
		8064: begin l_1 = -8;
				 l_2 = +14; end
		5517: begin l_1 = -8;
				 l_2 = -14; end
		2675: begin l_1 = +8;
				 l_2 = +15; end
		11418: begin l_1 = +8;
				 l_2 = -15; end
		2419: begin l_1 = -8;
				 l_2 = +15; end
		11162: begin l_1 = -8;
				 l_2 = -15; end
		5222: begin l_1 = +8;
				 l_2 = +16; end
		8871: begin l_1 = +8;
				 l_2 = -16; end
		4966: begin l_1 = -8;
				 l_2 = +16; end
		8615: begin l_1 = -8;
				 l_2 = -16; end
		10316: begin l_1 = +8;
				 l_2 = +17; end
		3777: begin l_1 = +8;
				 l_2 = -17; end
		10060: begin l_1 = -8;
				 l_2 = +17; end
		3521: begin l_1 = -8;
				 l_2 = -17; end
		6667: begin l_1 = +8;
				 l_2 = +18; end
		7426: begin l_1 = +8;
				 l_2 = -18; end
		6411: begin l_1 = -8;
				 l_2 = +18; end
		7170: begin l_1 = -8;
				 l_2 = -18; end
		13206: begin l_1 = +8;
				 l_2 = +19; end
		887: begin l_1 = +8;
				 l_2 = -19; end
		12950: begin l_1 = -8;
				 l_2 = +19; end
		631: begin l_1 = -8;
				 l_2 = -19; end
		12447: begin l_1 = +8;
				 l_2 = +20; end
		1646: begin l_1 = +8;
				 l_2 = -20; end
		12191: begin l_1 = -8;
				 l_2 = +20; end
		1390: begin l_1 = -8;
				 l_2 = -20; end
		10929: begin l_1 = +8;
				 l_2 = +21; end
		3164: begin l_1 = +8;
				 l_2 = -21; end
		10673: begin l_1 = -8;
				 l_2 = +21; end
		2908: begin l_1 = -8;
				 l_2 = -21; end
		7893: begin l_1 = +8;
				 l_2 = +22; end
		6200: begin l_1 = +8;
				 l_2 = -22; end
		7637: begin l_1 = -8;
				 l_2 = +22; end
		5944: begin l_1 = -8;
				 l_2 = -22; end
		1821: begin l_1 = +8;
				 l_2 = +23; end
		12272: begin l_1 = +8;
				 l_2 = -23; end
		1565: begin l_1 = -8;
				 l_2 = +23; end
		12016: begin l_1 = -8;
				 l_2 = -23; end
		3514: begin l_1 = +8;
				 l_2 = +24; end
		10579: begin l_1 = +8;
				 l_2 = -24; end
		3258: begin l_1 = -8;
				 l_2 = +24; end
		10323: begin l_1 = -8;
				 l_2 = -24; end
		6900: begin l_1 = +8;
				 l_2 = +25; end
		7193: begin l_1 = +8;
				 l_2 = -25; end
		6644: begin l_1 = -8;
				 l_2 = +25; end
		6937: begin l_1 = -8;
				 l_2 = -25; end
		13672: begin l_1 = +8;
				 l_2 = +26; end
		421: begin l_1 = +8;
				 l_2 = -26; end
		13416: begin l_1 = -8;
				 l_2 = +26; end
		165: begin l_1 = -8;
				 l_2 = -26; end
		13379: begin l_1 = +8;
				 l_2 = +27; end
		714: begin l_1 = +8;
				 l_2 = -27; end
		13123: begin l_1 = -8;
				 l_2 = +27; end
		458: begin l_1 = -8;
				 l_2 = -27; end
		12793: begin l_1 = +8;
				 l_2 = +28; end
		1300: begin l_1 = +8;
				 l_2 = -28; end
		12537: begin l_1 = -8;
				 l_2 = +28; end
		1044: begin l_1 = -8;
				 l_2 = -28; end
		11621: begin l_1 = +8;
				 l_2 = +29; end
		2472: begin l_1 = +8;
				 l_2 = -29; end
		11365: begin l_1 = -8;
				 l_2 = +29; end
		2216: begin l_1 = -8;
				 l_2 = -29; end
		9277: begin l_1 = +8;
				 l_2 = +30; end
		4816: begin l_1 = +8;
				 l_2 = -30; end
		9021: begin l_1 = -8;
				 l_2 = +30; end
		4560: begin l_1 = -8;
				 l_2 = -30; end
		4589: begin l_1 = +8;
				 l_2 = +31; end
		9504: begin l_1 = +8;
				 l_2 = -31; end
		4333: begin l_1 = -8;
				 l_2 = +31; end
		9248: begin l_1 = -8;
				 l_2 = -31; end
		9050: begin l_1 = +8;
				 l_2 = +32; end
		5043: begin l_1 = +8;
				 l_2 = -32; end
		8794: begin l_1 = -8;
				 l_2 = +32; end
		4787: begin l_1 = -8;
				 l_2 = -32; end
		4135: begin l_1 = +8;
				 l_2 = +33; end
		9958: begin l_1 = +8;
				 l_2 = -33; end
		3879: begin l_1 = -8;
				 l_2 = +33; end
		9702: begin l_1 = -8;
				 l_2 = -33; end
		8142: begin l_1 = +8;
				 l_2 = +34; end
		5951: begin l_1 = +8;
				 l_2 = -34; end
		7886: begin l_1 = -8;
				 l_2 = +34; end
		5695: begin l_1 = -8;
				 l_2 = -34; end
		2319: begin l_1 = +8;
				 l_2 = +35; end
		11774: begin l_1 = +8;
				 l_2 = -35; end
		2063: begin l_1 = -8;
				 l_2 = +35; end
		11518: begin l_1 = -8;
				 l_2 = -35; end
		4510: begin l_1 = +8;
				 l_2 = +36; end
		9583: begin l_1 = +8;
				 l_2 = -36; end
		4254: begin l_1 = -8;
				 l_2 = +36; end
		9327: begin l_1 = -8;
				 l_2 = -36; end
		8892: begin l_1 = +8;
				 l_2 = +37; end
		5201: begin l_1 = +8;
				 l_2 = -37; end
		8636: begin l_1 = -8;
				 l_2 = +37; end
		4945: begin l_1 = -8;
				 l_2 = -37; end
		3819: begin l_1 = +8;
				 l_2 = +38; end
		10274: begin l_1 = +8;
				 l_2 = -38; end
		3563: begin l_1 = -8;
				 l_2 = +38; end
		10018: begin l_1 = -8;
				 l_2 = -38; end
		768: begin l_1 = -9;
				 l_2 = +11; end
		13069: begin l_1 = -9;
				 l_2 = -10; end
		1280: begin l_1 = +9;
				 l_2 = +11; end
		12557: begin l_1 = -9;
				 l_2 = -11; end
		2304: begin l_1 = +9;
				 l_2 = +12; end
		12045: begin l_1 = +9;
				 l_2 = -12; end
		1792: begin l_1 = -9;
				 l_2 = +12; end
		11533: begin l_1 = -9;
				 l_2 = -12; end
		4352: begin l_1 = +9;
				 l_2 = +13; end
		9997: begin l_1 = +9;
				 l_2 = -13; end
		3840: begin l_1 = -9;
				 l_2 = +13; end
		9485: begin l_1 = -9;
				 l_2 = -13; end
		8448: begin l_1 = +9;
				 l_2 = +14; end
		5901: begin l_1 = +9;
				 l_2 = -14; end
		7936: begin l_1 = -9;
				 l_2 = +14; end
		5389: begin l_1 = -9;
				 l_2 = -14; end
		2803: begin l_1 = +9;
				 l_2 = +15; end
		11546: begin l_1 = +9;
				 l_2 = -15; end
		2291: begin l_1 = -9;
				 l_2 = +15; end
		11034: begin l_1 = -9;
				 l_2 = -15; end
		5350: begin l_1 = +9;
				 l_2 = +16; end
		8999: begin l_1 = +9;
				 l_2 = -16; end
		4838: begin l_1 = -9;
				 l_2 = +16; end
		8487: begin l_1 = -9;
				 l_2 = -16; end
		10444: begin l_1 = +9;
				 l_2 = +17; end
		3905: begin l_1 = +9;
				 l_2 = -17; end
		9932: begin l_1 = -9;
				 l_2 = +17; end
		3393: begin l_1 = -9;
				 l_2 = -17; end
		6795: begin l_1 = +9;
				 l_2 = +18; end
		7554: begin l_1 = +9;
				 l_2 = -18; end
		6283: begin l_1 = -9;
				 l_2 = +18; end
		7042: begin l_1 = -9;
				 l_2 = -18; end
		13334: begin l_1 = +9;
				 l_2 = +19; end
		1015: begin l_1 = +9;
				 l_2 = -19; end
		12822: begin l_1 = -9;
				 l_2 = +19; end
		503: begin l_1 = -9;
				 l_2 = -19; end
		12575: begin l_1 = +9;
				 l_2 = +20; end
		1774: begin l_1 = +9;
				 l_2 = -20; end
		12063: begin l_1 = -9;
				 l_2 = +20; end
		1262: begin l_1 = -9;
				 l_2 = -20; end
		11057: begin l_1 = +9;
				 l_2 = +21; end
		3292: begin l_1 = +9;
				 l_2 = -21; end
		10545: begin l_1 = -9;
				 l_2 = +21; end
		2780: begin l_1 = -9;
				 l_2 = -21; end
		8021: begin l_1 = +9;
				 l_2 = +22; end
		6328: begin l_1 = +9;
				 l_2 = -22; end
		7509: begin l_1 = -9;
				 l_2 = +22; end
		5816: begin l_1 = -9;
				 l_2 = -22; end
		1949: begin l_1 = +9;
				 l_2 = +23; end
		12400: begin l_1 = +9;
				 l_2 = -23; end
		1437: begin l_1 = -9;
				 l_2 = +23; end
		11888: begin l_1 = -9;
				 l_2 = -23; end
		3642: begin l_1 = +9;
				 l_2 = +24; end
		10707: begin l_1 = +9;
				 l_2 = -24; end
		3130: begin l_1 = -9;
				 l_2 = +24; end
		10195: begin l_1 = -9;
				 l_2 = -24; end
		7028: begin l_1 = +9;
				 l_2 = +25; end
		7321: begin l_1 = +9;
				 l_2 = -25; end
		6516: begin l_1 = -9;
				 l_2 = +25; end
		6809: begin l_1 = -9;
				 l_2 = -25; end
		13800: begin l_1 = +9;
				 l_2 = +26; end
		549: begin l_1 = +9;
				 l_2 = -26; end
		13288: begin l_1 = -9;
				 l_2 = +26; end
		37: begin l_1 = -9;
				 l_2 = -26; end
		13507: begin l_1 = +9;
				 l_2 = +27; end
		842: begin l_1 = +9;
				 l_2 = -27; end
		12995: begin l_1 = -9;
				 l_2 = +27; end
		330: begin l_1 = -9;
				 l_2 = -27; end
		12921: begin l_1 = +9;
				 l_2 = +28; end
		1428: begin l_1 = +9;
				 l_2 = -28; end
		12409: begin l_1 = -9;
				 l_2 = +28; end
		916: begin l_1 = -9;
				 l_2 = -28; end
		11749: begin l_1 = +9;
				 l_2 = +29; end
		2600: begin l_1 = +9;
				 l_2 = -29; end
		11237: begin l_1 = -9;
				 l_2 = +29; end
		2088: begin l_1 = -9;
				 l_2 = -29; end
		9405: begin l_1 = +9;
				 l_2 = +30; end
		4944: begin l_1 = +9;
				 l_2 = -30; end
		8893: begin l_1 = -9;
				 l_2 = +30; end
		4432: begin l_1 = -9;
				 l_2 = -30; end
		4717: begin l_1 = +9;
				 l_2 = +31; end
		9632: begin l_1 = +9;
				 l_2 = -31; end
		4205: begin l_1 = -9;
				 l_2 = +31; end
		9120: begin l_1 = -9;
				 l_2 = -31; end
		9178: begin l_1 = +9;
				 l_2 = +32; end
		5171: begin l_1 = +9;
				 l_2 = -32; end
		8666: begin l_1 = -9;
				 l_2 = +32; end
		4659: begin l_1 = -9;
				 l_2 = -32; end
		4263: begin l_1 = +9;
				 l_2 = +33; end
		10086: begin l_1 = +9;
				 l_2 = -33; end
		3751: begin l_1 = -9;
				 l_2 = +33; end
		9574: begin l_1 = -9;
				 l_2 = -33; end
		8270: begin l_1 = +9;
				 l_2 = +34; end
		6079: begin l_1 = +9;
				 l_2 = -34; end
		7758: begin l_1 = -9;
				 l_2 = +34; end
		5567: begin l_1 = -9;
				 l_2 = -34; end
		2447: begin l_1 = +9;
				 l_2 = +35; end
		11902: begin l_1 = +9;
				 l_2 = -35; end
		1935: begin l_1 = -9;
				 l_2 = +35; end
		11390: begin l_1 = -9;
				 l_2 = -35; end
		4638: begin l_1 = +9;
				 l_2 = +36; end
		9711: begin l_1 = +9;
				 l_2 = -36; end
		4126: begin l_1 = -9;
				 l_2 = +36; end
		9199: begin l_1 = -9;
				 l_2 = -36; end
		9020: begin l_1 = +9;
				 l_2 = +37; end
		5329: begin l_1 = +9;
				 l_2 = -37; end
		8508: begin l_1 = -9;
				 l_2 = +37; end
		4817: begin l_1 = -9;
				 l_2 = -37; end
		3947: begin l_1 = +9;
				 l_2 = +38; end
		10402: begin l_1 = +9;
				 l_2 = -38; end
		3435: begin l_1 = -9;
				 l_2 = +38; end
		9890: begin l_1 = -9;
				 l_2 = -38; end
		1536: begin l_1 = -10;
				 l_2 = +12; end
		12301: begin l_1 = -10;
				 l_2 = -11; end
		2560: begin l_1 = +10;
				 l_2 = +12; end
		11277: begin l_1 = -10;
				 l_2 = -12; end
		4608: begin l_1 = +10;
				 l_2 = +13; end
		10253: begin l_1 = +10;
				 l_2 = -13; end
		3584: begin l_1 = -10;
				 l_2 = +13; end
		9229: begin l_1 = -10;
				 l_2 = -13; end
		8704: begin l_1 = +10;
				 l_2 = +14; end
		6157: begin l_1 = +10;
				 l_2 = -14; end
		7680: begin l_1 = -10;
				 l_2 = +14; end
		5133: begin l_1 = -10;
				 l_2 = -14; end
		3059: begin l_1 = +10;
				 l_2 = +15; end
		11802: begin l_1 = +10;
				 l_2 = -15; end
		2035: begin l_1 = -10;
				 l_2 = +15; end
		10778: begin l_1 = -10;
				 l_2 = -15; end
		5606: begin l_1 = +10;
				 l_2 = +16; end
		9255: begin l_1 = +10;
				 l_2 = -16; end
		4582: begin l_1 = -10;
				 l_2 = +16; end
		8231: begin l_1 = -10;
				 l_2 = -16; end
		10700: begin l_1 = +10;
				 l_2 = +17; end
		4161: begin l_1 = +10;
				 l_2 = -17; end
		9676: begin l_1 = -10;
				 l_2 = +17; end
		3137: begin l_1 = -10;
				 l_2 = -17; end
		7051: begin l_1 = +10;
				 l_2 = +18; end
		7810: begin l_1 = +10;
				 l_2 = -18; end
		6027: begin l_1 = -10;
				 l_2 = +18; end
		6786: begin l_1 = -10;
				 l_2 = -18; end
		13590: begin l_1 = +10;
				 l_2 = +19; end
		1271: begin l_1 = +10;
				 l_2 = -19; end
		12566: begin l_1 = -10;
				 l_2 = +19; end
		247: begin l_1 = -10;
				 l_2 = -19; end
		12831: begin l_1 = +10;
				 l_2 = +20; end
		2030: begin l_1 = +10;
				 l_2 = -20; end
		11807: begin l_1 = -10;
				 l_2 = +20; end
		1006: begin l_1 = -10;
				 l_2 = -20; end
		11313: begin l_1 = +10;
				 l_2 = +21; end
		3548: begin l_1 = +10;
				 l_2 = -21; end
		10289: begin l_1 = -10;
				 l_2 = +21; end
		2524: begin l_1 = -10;
				 l_2 = -21; end
		8277: begin l_1 = +10;
				 l_2 = +22; end
		6584: begin l_1 = +10;
				 l_2 = -22; end
		7253: begin l_1 = -10;
				 l_2 = +22; end
		5560: begin l_1 = -10;
				 l_2 = -22; end
		2205: begin l_1 = +10;
				 l_2 = +23; end
		12656: begin l_1 = +10;
				 l_2 = -23; end
		1181: begin l_1 = -10;
				 l_2 = +23; end
		11632: begin l_1 = -10;
				 l_2 = -23; end
		3898: begin l_1 = +10;
				 l_2 = +24; end
		10963: begin l_1 = +10;
				 l_2 = -24; end
		2874: begin l_1 = -10;
				 l_2 = +24; end
		9939: begin l_1 = -10;
				 l_2 = -24; end
		7284: begin l_1 = +10;
				 l_2 = +25; end
		7577: begin l_1 = +10;
				 l_2 = -25; end
		6260: begin l_1 = -10;
				 l_2 = +25; end
		6553: begin l_1 = -10;
				 l_2 = -25; end
		219: begin l_1 = +10;
				 l_2 = +26; end
		805: begin l_1 = +10;
				 l_2 = -26; end
		13032: begin l_1 = -10;
				 l_2 = +26; end
		13618: begin l_1 = -10;
				 l_2 = -26; end
		13763: begin l_1 = +10;
				 l_2 = +27; end
		1098: begin l_1 = +10;
				 l_2 = -27; end
		12739: begin l_1 = -10;
				 l_2 = +27; end
		74: begin l_1 = -10;
				 l_2 = -27; end
		13177: begin l_1 = +10;
				 l_2 = +28; end
		1684: begin l_1 = +10;
				 l_2 = -28; end
		12153: begin l_1 = -10;
				 l_2 = +28; end
		660: begin l_1 = -10;
				 l_2 = -28; end
		12005: begin l_1 = +10;
				 l_2 = +29; end
		2856: begin l_1 = +10;
				 l_2 = -29; end
		10981: begin l_1 = -10;
				 l_2 = +29; end
		1832: begin l_1 = -10;
				 l_2 = -29; end
		9661: begin l_1 = +10;
				 l_2 = +30; end
		5200: begin l_1 = +10;
				 l_2 = -30; end
		8637: begin l_1 = -10;
				 l_2 = +30; end
		4176: begin l_1 = -10;
				 l_2 = -30; end
		4973: begin l_1 = +10;
				 l_2 = +31; end
		9888: begin l_1 = +10;
				 l_2 = -31; end
		3949: begin l_1 = -10;
				 l_2 = +31; end
		8864: begin l_1 = -10;
				 l_2 = -31; end
		9434: begin l_1 = +10;
				 l_2 = +32; end
		5427: begin l_1 = +10;
				 l_2 = -32; end
		8410: begin l_1 = -10;
				 l_2 = +32; end
		4403: begin l_1 = -10;
				 l_2 = -32; end
		4519: begin l_1 = +10;
				 l_2 = +33; end
		10342: begin l_1 = +10;
				 l_2 = -33; end
		3495: begin l_1 = -10;
				 l_2 = +33; end
		9318: begin l_1 = -10;
				 l_2 = -33; end
		8526: begin l_1 = +10;
				 l_2 = +34; end
		6335: begin l_1 = +10;
				 l_2 = -34; end
		7502: begin l_1 = -10;
				 l_2 = +34; end
		5311: begin l_1 = -10;
				 l_2 = -34; end
		2703: begin l_1 = +10;
				 l_2 = +35; end
		12158: begin l_1 = +10;
				 l_2 = -35; end
		1679: begin l_1 = -10;
				 l_2 = +35; end
		11134: begin l_1 = -10;
				 l_2 = -35; end
		4894: begin l_1 = +10;
				 l_2 = +36; end
		9967: begin l_1 = +10;
				 l_2 = -36; end
		3870: begin l_1 = -10;
				 l_2 = +36; end
		8943: begin l_1 = -10;
				 l_2 = -36; end
		9276: begin l_1 = +10;
				 l_2 = +37; end
		5585: begin l_1 = +10;
				 l_2 = -37; end
		8252: begin l_1 = -10;
				 l_2 = +37; end
		4561: begin l_1 = -10;
				 l_2 = -37; end
		4203: begin l_1 = +10;
				 l_2 = +38; end
		10658: begin l_1 = +10;
				 l_2 = -38; end
		3179: begin l_1 = -10;
				 l_2 = +38; end
		9634: begin l_1 = -10;
				 l_2 = -38; end
		3072: begin l_1 = -11;
				 l_2 = +13; end
		10765: begin l_1 = -11;
				 l_2 = -12; end
		5120: begin l_1 = +11;
				 l_2 = +13; end
		8717: begin l_1 = -11;
				 l_2 = -13; end
		9216: begin l_1 = +11;
				 l_2 = +14; end
		6669: begin l_1 = +11;
				 l_2 = -14; end
		7168: begin l_1 = -11;
				 l_2 = +14; end
		4621: begin l_1 = -11;
				 l_2 = -14; end
		3571: begin l_1 = +11;
				 l_2 = +15; end
		12314: begin l_1 = +11;
				 l_2 = -15; end
		1523: begin l_1 = -11;
				 l_2 = +15; end
		10266: begin l_1 = -11;
				 l_2 = -15; end
		6118: begin l_1 = +11;
				 l_2 = +16; end
		9767: begin l_1 = +11;
				 l_2 = -16; end
		4070: begin l_1 = -11;
				 l_2 = +16; end
		7719: begin l_1 = -11;
				 l_2 = -16; end
		11212: begin l_1 = +11;
				 l_2 = +17; end
		4673: begin l_1 = +11;
				 l_2 = -17; end
		9164: begin l_1 = -11;
				 l_2 = +17; end
		2625: begin l_1 = -11;
				 l_2 = -17; end
		7563: begin l_1 = +11;
				 l_2 = +18; end
		8322: begin l_1 = +11;
				 l_2 = -18; end
		5515: begin l_1 = -11;
				 l_2 = +18; end
		6274: begin l_1 = -11;
				 l_2 = -18; end
		265: begin l_1 = +11;
				 l_2 = +19; end
		1783: begin l_1 = +11;
				 l_2 = -19; end
		12054: begin l_1 = -11;
				 l_2 = +19; end
		13572: begin l_1 = -11;
				 l_2 = -19; end
		13343: begin l_1 = +11;
				 l_2 = +20; end
		2542: begin l_1 = +11;
				 l_2 = -20; end
		11295: begin l_1 = -11;
				 l_2 = +20; end
		494: begin l_1 = -11;
				 l_2 = -20; end
		11825: begin l_1 = +11;
				 l_2 = +21; end
		4060: begin l_1 = +11;
				 l_2 = -21; end
		9777: begin l_1 = -11;
				 l_2 = +21; end
		2012: begin l_1 = -11;
				 l_2 = -21; end
		8789: begin l_1 = +11;
				 l_2 = +22; end
		7096: begin l_1 = +11;
				 l_2 = -22; end
		6741: begin l_1 = -11;
				 l_2 = +22; end
		5048: begin l_1 = -11;
				 l_2 = -22; end
		2717: begin l_1 = +11;
				 l_2 = +23; end
		13168: begin l_1 = +11;
				 l_2 = -23; end
		669: begin l_1 = -11;
				 l_2 = +23; end
		11120: begin l_1 = -11;
				 l_2 = -23; end
		4410: begin l_1 = +11;
				 l_2 = +24; end
		11475: begin l_1 = +11;
				 l_2 = -24; end
		2362: begin l_1 = -11;
				 l_2 = +24; end
		9427: begin l_1 = -11;
				 l_2 = -24; end
		7796: begin l_1 = +11;
				 l_2 = +25; end
		8089: begin l_1 = +11;
				 l_2 = -25; end
		5748: begin l_1 = -11;
				 l_2 = +25; end
		6041: begin l_1 = -11;
				 l_2 = -25; end
		731: begin l_1 = +11;
				 l_2 = +26; end
		1317: begin l_1 = +11;
				 l_2 = -26; end
		12520: begin l_1 = -11;
				 l_2 = +26; end
		13106: begin l_1 = -11;
				 l_2 = -26; end
		438: begin l_1 = +11;
				 l_2 = +27; end
		1610: begin l_1 = +11;
				 l_2 = -27; end
		12227: begin l_1 = -11;
				 l_2 = +27; end
		13399: begin l_1 = -11;
				 l_2 = -27; end
		13689: begin l_1 = +11;
				 l_2 = +28; end
		2196: begin l_1 = +11;
				 l_2 = -28; end
		11641: begin l_1 = -11;
				 l_2 = +28; end
		148: begin l_1 = -11;
				 l_2 = -28; end
		12517: begin l_1 = +11;
				 l_2 = +29; end
		3368: begin l_1 = +11;
				 l_2 = -29; end
		10469: begin l_1 = -11;
				 l_2 = +29; end
		1320: begin l_1 = -11;
				 l_2 = -29; end
		10173: begin l_1 = +11;
				 l_2 = +30; end
		5712: begin l_1 = +11;
				 l_2 = -30; end
		8125: begin l_1 = -11;
				 l_2 = +30; end
		3664: begin l_1 = -11;
				 l_2 = -30; end
		5485: begin l_1 = +11;
				 l_2 = +31; end
		10400: begin l_1 = +11;
				 l_2 = -31; end
		3437: begin l_1 = -11;
				 l_2 = +31; end
		8352: begin l_1 = -11;
				 l_2 = -31; end
		9946: begin l_1 = +11;
				 l_2 = +32; end
		5939: begin l_1 = +11;
				 l_2 = -32; end
		7898: begin l_1 = -11;
				 l_2 = +32; end
		3891: begin l_1 = -11;
				 l_2 = -32; end
		5031: begin l_1 = +11;
				 l_2 = +33; end
		10854: begin l_1 = +11;
				 l_2 = -33; end
		2983: begin l_1 = -11;
				 l_2 = +33; end
		8806: begin l_1 = -11;
				 l_2 = -33; end
		9038: begin l_1 = +11;
				 l_2 = +34; end
		6847: begin l_1 = +11;
				 l_2 = -34; end
		6990: begin l_1 = -11;
				 l_2 = +34; end
		4799: begin l_1 = -11;
				 l_2 = -34; end
		3215: begin l_1 = +11;
				 l_2 = +35; end
		12670: begin l_1 = +11;
				 l_2 = -35; end
		1167: begin l_1 = -11;
				 l_2 = +35; end
		10622: begin l_1 = -11;
				 l_2 = -35; end
		5406: begin l_1 = +11;
				 l_2 = +36; end
		10479: begin l_1 = +11;
				 l_2 = -36; end
		3358: begin l_1 = -11;
				 l_2 = +36; end
		8431: begin l_1 = -11;
				 l_2 = -36; end
		9788: begin l_1 = +11;
				 l_2 = +37; end
		6097: begin l_1 = +11;
				 l_2 = -37; end
		7740: begin l_1 = -11;
				 l_2 = +37; end
		4049: begin l_1 = -11;
				 l_2 = -37; end
		4715: begin l_1 = +11;
				 l_2 = +38; end
		11170: begin l_1 = +11;
				 l_2 = -38; end
		2667: begin l_1 = -11;
				 l_2 = +38; end
		9122: begin l_1 = -11;
				 l_2 = -38; end
		6144: begin l_1 = -12;
				 l_2 = +14; end
		7693: begin l_1 = -12;
				 l_2 = -13; end
		10240: begin l_1 = +12;
				 l_2 = +14; end
		3597: begin l_1 = -12;
				 l_2 = -14; end
		4595: begin l_1 = +12;
				 l_2 = +15; end
		13338: begin l_1 = +12;
				 l_2 = -15; end
		499: begin l_1 = -12;
				 l_2 = +15; end
		9242: begin l_1 = -12;
				 l_2 = -15; end
		7142: begin l_1 = +12;
				 l_2 = +16; end
		10791: begin l_1 = +12;
				 l_2 = -16; end
		3046: begin l_1 = -12;
				 l_2 = +16; end
		6695: begin l_1 = -12;
				 l_2 = -16; end
		12236: begin l_1 = +12;
				 l_2 = +17; end
		5697: begin l_1 = +12;
				 l_2 = -17; end
		8140: begin l_1 = -12;
				 l_2 = +17; end
		1601: begin l_1 = -12;
				 l_2 = -17; end
		8587: begin l_1 = +12;
				 l_2 = +18; end
		9346: begin l_1 = +12;
				 l_2 = -18; end
		4491: begin l_1 = -12;
				 l_2 = +18; end
		5250: begin l_1 = -12;
				 l_2 = -18; end
		1289: begin l_1 = +12;
				 l_2 = +19; end
		2807: begin l_1 = +12;
				 l_2 = -19; end
		11030: begin l_1 = -12;
				 l_2 = +19; end
		12548: begin l_1 = -12;
				 l_2 = -19; end
		530: begin l_1 = +12;
				 l_2 = +20; end
		3566: begin l_1 = +12;
				 l_2 = -20; end
		10271: begin l_1 = -12;
				 l_2 = +20; end
		13307: begin l_1 = -12;
				 l_2 = -20; end
		12849: begin l_1 = +12;
				 l_2 = +21; end
		5084: begin l_1 = +12;
				 l_2 = -21; end
		8753: begin l_1 = -12;
				 l_2 = +21; end
		988: begin l_1 = -12;
				 l_2 = -21; end
		9813: begin l_1 = +12;
				 l_2 = +22; end
		8120: begin l_1 = +12;
				 l_2 = -22; end
		5717: begin l_1 = -12;
				 l_2 = +22; end
		4024: begin l_1 = -12;
				 l_2 = -22; end
		3741: begin l_1 = +12;
				 l_2 = +23; end
		355: begin l_1 = +12;
				 l_2 = -23; end
		13482: begin l_1 = -12;
				 l_2 = +23; end
		10096: begin l_1 = -12;
				 l_2 = -23; end
		5434: begin l_1 = +12;
				 l_2 = +24; end
		12499: begin l_1 = +12;
				 l_2 = -24; end
		1338: begin l_1 = -12;
				 l_2 = +24; end
		8403: begin l_1 = -12;
				 l_2 = -24; end
		8820: begin l_1 = +12;
				 l_2 = +25; end
		9113: begin l_1 = +12;
				 l_2 = -25; end
		4724: begin l_1 = -12;
				 l_2 = +25; end
		5017: begin l_1 = -12;
				 l_2 = -25; end
		1755: begin l_1 = +12;
				 l_2 = +26; end
		2341: begin l_1 = +12;
				 l_2 = -26; end
		11496: begin l_1 = -12;
				 l_2 = +26; end
		12082: begin l_1 = -12;
				 l_2 = -26; end
		1462: begin l_1 = +12;
				 l_2 = +27; end
		2634: begin l_1 = +12;
				 l_2 = -27; end
		11203: begin l_1 = -12;
				 l_2 = +27; end
		12375: begin l_1 = -12;
				 l_2 = -27; end
		876: begin l_1 = +12;
				 l_2 = +28; end
		3220: begin l_1 = +12;
				 l_2 = -28; end
		10617: begin l_1 = -12;
				 l_2 = +28; end
		12961: begin l_1 = -12;
				 l_2 = -28; end
		13541: begin l_1 = +12;
				 l_2 = +29; end
		4392: begin l_1 = +12;
				 l_2 = -29; end
		9445: begin l_1 = -12;
				 l_2 = +29; end
		296: begin l_1 = -12;
				 l_2 = -29; end
		11197: begin l_1 = +12;
				 l_2 = +30; end
		6736: begin l_1 = +12;
				 l_2 = -30; end
		7101: begin l_1 = -12;
				 l_2 = +30; end
		2640: begin l_1 = -12;
				 l_2 = -30; end
		6509: begin l_1 = +12;
				 l_2 = +31; end
		11424: begin l_1 = +12;
				 l_2 = -31; end
		2413: begin l_1 = -12;
				 l_2 = +31; end
		7328: begin l_1 = -12;
				 l_2 = -31; end
		10970: begin l_1 = +12;
				 l_2 = +32; end
		6963: begin l_1 = +12;
				 l_2 = -32; end
		6874: begin l_1 = -12;
				 l_2 = +32; end
		2867: begin l_1 = -12;
				 l_2 = -32; end
		6055: begin l_1 = +12;
				 l_2 = +33; end
		11878: begin l_1 = +12;
				 l_2 = -33; end
		1959: begin l_1 = -12;
				 l_2 = +33; end
		7782: begin l_1 = -12;
				 l_2 = -33; end
		10062: begin l_1 = +12;
				 l_2 = +34; end
		7871: begin l_1 = +12;
				 l_2 = -34; end
		5966: begin l_1 = -12;
				 l_2 = +34; end
		3775: begin l_1 = -12;
				 l_2 = -34; end
		4239: begin l_1 = +12;
				 l_2 = +35; end
		13694: begin l_1 = +12;
				 l_2 = -35; end
		143: begin l_1 = -12;
				 l_2 = +35; end
		9598: begin l_1 = -12;
				 l_2 = -35; end
		6430: begin l_1 = +12;
				 l_2 = +36; end
		11503: begin l_1 = +12;
				 l_2 = -36; end
		2334: begin l_1 = -12;
				 l_2 = +36; end
		7407: begin l_1 = -12;
				 l_2 = -36; end
		10812: begin l_1 = +12;
				 l_2 = +37; end
		7121: begin l_1 = +12;
				 l_2 = -37; end
		6716: begin l_1 = -12;
				 l_2 = +37; end
		3025: begin l_1 = -12;
				 l_2 = -37; end
		5739: begin l_1 = +12;
				 l_2 = +38; end
		12194: begin l_1 = +12;
				 l_2 = -38; end
		1643: begin l_1 = -12;
				 l_2 = +38; end
		8098: begin l_1 = -12;
				 l_2 = -38; end
		12288: begin l_1 = -13;
				 l_2 = +15; end
		1549: begin l_1 = -13;
				 l_2 = -14; end
		6643: begin l_1 = +13;
				 l_2 = +15; end
		7194: begin l_1 = -13;
				 l_2 = -15; end
		9190: begin l_1 = +13;
				 l_2 = +16; end
		12839: begin l_1 = +13;
				 l_2 = -16; end
		998: begin l_1 = -13;
				 l_2 = +16; end
		4647: begin l_1 = -13;
				 l_2 = -16; end
		447: begin l_1 = +13;
				 l_2 = +17; end
		7745: begin l_1 = +13;
				 l_2 = -17; end
		6092: begin l_1 = -13;
				 l_2 = +17; end
		13390: begin l_1 = -13;
				 l_2 = -17; end
		10635: begin l_1 = +13;
				 l_2 = +18; end
		11394: begin l_1 = +13;
				 l_2 = -18; end
		2443: begin l_1 = -13;
				 l_2 = +18; end
		3202: begin l_1 = -13;
				 l_2 = -18; end
		3337: begin l_1 = +13;
				 l_2 = +19; end
		4855: begin l_1 = +13;
				 l_2 = -19; end
		8982: begin l_1 = -13;
				 l_2 = +19; end
		10500: begin l_1 = -13;
				 l_2 = -19; end
		2578: begin l_1 = +13;
				 l_2 = +20; end
		5614: begin l_1 = +13;
				 l_2 = -20; end
		8223: begin l_1 = -13;
				 l_2 = +20; end
		11259: begin l_1 = -13;
				 l_2 = -20; end
		1060: begin l_1 = +13;
				 l_2 = +21; end
		7132: begin l_1 = +13;
				 l_2 = -21; end
		6705: begin l_1 = -13;
				 l_2 = +21; end
		12777: begin l_1 = -13;
				 l_2 = -21; end
		11861: begin l_1 = +13;
				 l_2 = +22; end
		10168: begin l_1 = +13;
				 l_2 = -22; end
		3669: begin l_1 = -13;
				 l_2 = +22; end
		1976: begin l_1 = -13;
				 l_2 = -22; end
		5789: begin l_1 = +13;
				 l_2 = +23; end
		2403: begin l_1 = +13;
				 l_2 = -23; end
		11434: begin l_1 = -13;
				 l_2 = +23; end
		8048: begin l_1 = -13;
				 l_2 = -23; end
		7482: begin l_1 = +13;
				 l_2 = +24; end
		710: begin l_1 = +13;
				 l_2 = -24; end
		13127: begin l_1 = -13;
				 l_2 = +24; end
		6355: begin l_1 = -13;
				 l_2 = -24; end
		10868: begin l_1 = +13;
				 l_2 = +25; end
		11161: begin l_1 = +13;
				 l_2 = -25; end
		2676: begin l_1 = -13;
				 l_2 = +25; end
		2969: begin l_1 = -13;
				 l_2 = -25; end
		3803: begin l_1 = +13;
				 l_2 = +26; end
		4389: begin l_1 = +13;
				 l_2 = -26; end
		9448: begin l_1 = -13;
				 l_2 = +26; end
		10034: begin l_1 = -13;
				 l_2 = -26; end
		3510: begin l_1 = +13;
				 l_2 = +27; end
		4682: begin l_1 = +13;
				 l_2 = -27; end
		9155: begin l_1 = -13;
				 l_2 = +27; end
		10327: begin l_1 = -13;
				 l_2 = -27; end
		2924: begin l_1 = +13;
				 l_2 = +28; end
		5268: begin l_1 = +13;
				 l_2 = -28; end
		8569: begin l_1 = -13;
				 l_2 = +28; end
		10913: begin l_1 = -13;
				 l_2 = -28; end
		1752: begin l_1 = +13;
				 l_2 = +29; end
		6440: begin l_1 = +13;
				 l_2 = -29; end
		7397: begin l_1 = -13;
				 l_2 = +29; end
		12085: begin l_1 = -13;
				 l_2 = -29; end
		13245: begin l_1 = +13;
				 l_2 = +30; end
		8784: begin l_1 = +13;
				 l_2 = -30; end
		5053: begin l_1 = -13;
				 l_2 = +30; end
		592: begin l_1 = -13;
				 l_2 = -30; end
		8557: begin l_1 = +13;
				 l_2 = +31; end
		13472: begin l_1 = +13;
				 l_2 = -31; end
		365: begin l_1 = -13;
				 l_2 = +31; end
		5280: begin l_1 = -13;
				 l_2 = -31; end
		13018: begin l_1 = +13;
				 l_2 = +32; end
		9011: begin l_1 = +13;
				 l_2 = -32; end
		4826: begin l_1 = -13;
				 l_2 = +32; end
		819: begin l_1 = -13;
				 l_2 = -32; end
		8103: begin l_1 = +13;
				 l_2 = +33; end
		89: begin l_1 = +13;
				 l_2 = -33; end
		13748: begin l_1 = -13;
				 l_2 = +33; end
		5734: begin l_1 = -13;
				 l_2 = -33; end
		12110: begin l_1 = +13;
				 l_2 = +34; end
		9919: begin l_1 = +13;
				 l_2 = -34; end
		3918: begin l_1 = -13;
				 l_2 = +34; end
		1727: begin l_1 = -13;
				 l_2 = -34; end
		6287: begin l_1 = +13;
				 l_2 = +35; end
		1905: begin l_1 = +13;
				 l_2 = -35; end
		11932: begin l_1 = -13;
				 l_2 = +35; end
		7550: begin l_1 = -13;
				 l_2 = -35; end
		8478: begin l_1 = +13;
				 l_2 = +36; end
		13551: begin l_1 = +13;
				 l_2 = -36; end
		286: begin l_1 = -13;
				 l_2 = +36; end
		5359: begin l_1 = -13;
				 l_2 = -36; end
		12860: begin l_1 = +13;
				 l_2 = +37; end
		9169: begin l_1 = +13;
				 l_2 = -37; end
		4668: begin l_1 = -13;
				 l_2 = +37; end
		977: begin l_1 = -13;
				 l_2 = -37; end
		7787: begin l_1 = +13;
				 l_2 = +38; end
		405: begin l_1 = +13;
				 l_2 = -38; end
		13432: begin l_1 = -13;
				 l_2 = +38; end
		6050: begin l_1 = -13;
				 l_2 = -38; end
		10739: begin l_1 = -14;
				 l_2 = +16; end
		3098: begin l_1 = -14;
				 l_2 = -15; end
		13286: begin l_1 = +14;
				 l_2 = +16; end
		551: begin l_1 = -14;
				 l_2 = -16; end
		4543: begin l_1 = +14;
				 l_2 = +17; end
		11841: begin l_1 = +14;
				 l_2 = -17; end
		1996: begin l_1 = -14;
				 l_2 = +17; end
		9294: begin l_1 = -14;
				 l_2 = -17; end
		894: begin l_1 = +14;
				 l_2 = +18; end
		1653: begin l_1 = +14;
				 l_2 = -18; end
		12184: begin l_1 = -14;
				 l_2 = +18; end
		12943: begin l_1 = -14;
				 l_2 = -18; end
		7433: begin l_1 = +14;
				 l_2 = +19; end
		8951: begin l_1 = +14;
				 l_2 = -19; end
		4886: begin l_1 = -14;
				 l_2 = +19; end
		6404: begin l_1 = -14;
				 l_2 = -19; end
		6674: begin l_1 = +14;
				 l_2 = +20; end
		9710: begin l_1 = +14;
				 l_2 = -20; end
		4127: begin l_1 = -14;
				 l_2 = +20; end
		7163: begin l_1 = -14;
				 l_2 = -20; end
		5156: begin l_1 = +14;
				 l_2 = +21; end
		11228: begin l_1 = +14;
				 l_2 = -21; end
		2609: begin l_1 = -14;
				 l_2 = +21; end
		8681: begin l_1 = -14;
				 l_2 = -21; end
		2120: begin l_1 = +14;
				 l_2 = +22; end
		427: begin l_1 = +14;
				 l_2 = -22; end
		13410: begin l_1 = -14;
				 l_2 = +22; end
		11717: begin l_1 = -14;
				 l_2 = -22; end
		9885: begin l_1 = +14;
				 l_2 = +23; end
		6499: begin l_1 = +14;
				 l_2 = -23; end
		7338: begin l_1 = -14;
				 l_2 = +23; end
		3952: begin l_1 = -14;
				 l_2 = -23; end
		11578: begin l_1 = +14;
				 l_2 = +24; end
		4806: begin l_1 = +14;
				 l_2 = -24; end
		9031: begin l_1 = -14;
				 l_2 = +24; end
		2259: begin l_1 = -14;
				 l_2 = -24; end
		1127: begin l_1 = +14;
				 l_2 = +25; end
		1420: begin l_1 = +14;
				 l_2 = -25; end
		12417: begin l_1 = -14;
				 l_2 = +25; end
		12710: begin l_1 = -14;
				 l_2 = -25; end
		7899: begin l_1 = +14;
				 l_2 = +26; end
		8485: begin l_1 = +14;
				 l_2 = -26; end
		5352: begin l_1 = -14;
				 l_2 = +26; end
		5938: begin l_1 = -14;
				 l_2 = -26; end
		7606: begin l_1 = +14;
				 l_2 = +27; end
		8778: begin l_1 = +14;
				 l_2 = -27; end
		5059: begin l_1 = -14;
				 l_2 = +27; end
		6231: begin l_1 = -14;
				 l_2 = -27; end
		7020: begin l_1 = +14;
				 l_2 = +28; end
		9364: begin l_1 = +14;
				 l_2 = -28; end
		4473: begin l_1 = -14;
				 l_2 = +28; end
		6817: begin l_1 = -14;
				 l_2 = -28; end
		5848: begin l_1 = +14;
				 l_2 = +29; end
		10536: begin l_1 = +14;
				 l_2 = -29; end
		3301: begin l_1 = -14;
				 l_2 = +29; end
		7989: begin l_1 = -14;
				 l_2 = -29; end
		3504: begin l_1 = +14;
				 l_2 = +30; end
		12880: begin l_1 = +14;
				 l_2 = -30; end
		957: begin l_1 = -14;
				 l_2 = +30; end
		10333: begin l_1 = -14;
				 l_2 = -30; end
		12653: begin l_1 = +14;
				 l_2 = +31; end
		3731: begin l_1 = +14;
				 l_2 = -31; end
		10106: begin l_1 = -14;
				 l_2 = +31; end
		1184: begin l_1 = -14;
				 l_2 = -31; end
		3277: begin l_1 = +14;
				 l_2 = +32; end
		13107: begin l_1 = +14;
				 l_2 = -32; end
		730: begin l_1 = -14;
				 l_2 = +32; end
		10560: begin l_1 = -14;
				 l_2 = -32; end
		12199: begin l_1 = +14;
				 l_2 = +33; end
		4185: begin l_1 = +14;
				 l_2 = -33; end
		9652: begin l_1 = -14;
				 l_2 = +33; end
		1638: begin l_1 = -14;
				 l_2 = -33; end
		2369: begin l_1 = +14;
				 l_2 = +34; end
		178: begin l_1 = +14;
				 l_2 = -34; end
		13659: begin l_1 = -14;
				 l_2 = +34; end
		11468: begin l_1 = -14;
				 l_2 = -34; end
		10383: begin l_1 = +14;
				 l_2 = +35; end
		6001: begin l_1 = +14;
				 l_2 = -35; end
		7836: begin l_1 = -14;
				 l_2 = +35; end
		3454: begin l_1 = -14;
				 l_2 = -35; end
		12574: begin l_1 = +14;
				 l_2 = +36; end
		3810: begin l_1 = +14;
				 l_2 = -36; end
		10027: begin l_1 = -14;
				 l_2 = +36; end
		1263: begin l_1 = -14;
				 l_2 = -36; end
		3119: begin l_1 = +14;
				 l_2 = +37; end
		13265: begin l_1 = +14;
				 l_2 = -37; end
		572: begin l_1 = -14;
				 l_2 = +37; end
		10718: begin l_1 = -14;
				 l_2 = -37; end
		11883: begin l_1 = +14;
				 l_2 = +38; end
		4501: begin l_1 = +14;
				 l_2 = -38; end
		9336: begin l_1 = -14;
				 l_2 = +38; end
		1954: begin l_1 = -14;
				 l_2 = -38; end
		7641: begin l_1 = -15;
				 l_2 = +17; end
		6196: begin l_1 = -15;
				 l_2 = -16; end
		12735: begin l_1 = +15;
				 l_2 = +17; end
		1102: begin l_1 = -15;
				 l_2 = -17; end
		9086: begin l_1 = +15;
				 l_2 = +18; end
		9845: begin l_1 = +15;
				 l_2 = -18; end
		3992: begin l_1 = -15;
				 l_2 = +18; end
		4751: begin l_1 = -15;
				 l_2 = -18; end
		1788: begin l_1 = +15;
				 l_2 = +19; end
		3306: begin l_1 = +15;
				 l_2 = -19; end
		10531: begin l_1 = -15;
				 l_2 = +19; end
		12049: begin l_1 = -15;
				 l_2 = -19; end
		1029: begin l_1 = +15;
				 l_2 = +20; end
		4065: begin l_1 = +15;
				 l_2 = -20; end
		9772: begin l_1 = -15;
				 l_2 = +20; end
		12808: begin l_1 = -15;
				 l_2 = -20; end
		13348: begin l_1 = +15;
				 l_2 = +21; end
		5583: begin l_1 = +15;
				 l_2 = -21; end
		8254: begin l_1 = -15;
				 l_2 = +21; end
		489: begin l_1 = -15;
				 l_2 = -21; end
		10312: begin l_1 = +15;
				 l_2 = +22; end
		8619: begin l_1 = +15;
				 l_2 = -22; end
		5218: begin l_1 = -15;
				 l_2 = +22; end
		3525: begin l_1 = -15;
				 l_2 = -22; end
		4240: begin l_1 = +15;
				 l_2 = +23; end
		854: begin l_1 = +15;
				 l_2 = -23; end
		12983: begin l_1 = -15;
				 l_2 = +23; end
		9597: begin l_1 = -15;
				 l_2 = -23; end
		5933: begin l_1 = +15;
				 l_2 = +24; end
		12998: begin l_1 = +15;
				 l_2 = -24; end
		839: begin l_1 = -15;
				 l_2 = +24; end
		7904: begin l_1 = -15;
				 l_2 = -24; end
		9319: begin l_1 = +15;
				 l_2 = +25; end
		9612: begin l_1 = +15;
				 l_2 = -25; end
		4225: begin l_1 = -15;
				 l_2 = +25; end
		4518: begin l_1 = -15;
				 l_2 = -25; end
		2254: begin l_1 = +15;
				 l_2 = +26; end
		2840: begin l_1 = +15;
				 l_2 = -26; end
		10997: begin l_1 = -15;
				 l_2 = +26; end
		11583: begin l_1 = -15;
				 l_2 = -26; end
		1961: begin l_1 = +15;
				 l_2 = +27; end
		3133: begin l_1 = +15;
				 l_2 = -27; end
		10704: begin l_1 = -15;
				 l_2 = +27; end
		11876: begin l_1 = -15;
				 l_2 = -27; end
		1375: begin l_1 = +15;
				 l_2 = +28; end
		3719: begin l_1 = +15;
				 l_2 = -28; end
		10118: begin l_1 = -15;
				 l_2 = +28; end
		12462: begin l_1 = -15;
				 l_2 = -28; end
		203: begin l_1 = +15;
				 l_2 = +29; end
		4891: begin l_1 = +15;
				 l_2 = -29; end
		8946: begin l_1 = -15;
				 l_2 = +29; end
		13634: begin l_1 = -15;
				 l_2 = -29; end
		11696: begin l_1 = +15;
				 l_2 = +30; end
		7235: begin l_1 = +15;
				 l_2 = -30; end
		6602: begin l_1 = -15;
				 l_2 = +30; end
		2141: begin l_1 = -15;
				 l_2 = -30; end
		7008: begin l_1 = +15;
				 l_2 = +31; end
		11923: begin l_1 = +15;
				 l_2 = -31; end
		1914: begin l_1 = -15;
				 l_2 = +31; end
		6829: begin l_1 = -15;
				 l_2 = -31; end
		11469: begin l_1 = +15;
				 l_2 = +32; end
		7462: begin l_1 = +15;
				 l_2 = -32; end
		6375: begin l_1 = -15;
				 l_2 = +32; end
		2368: begin l_1 = -15;
				 l_2 = -32; end
		6554: begin l_1 = +15;
				 l_2 = +33; end
		12377: begin l_1 = +15;
				 l_2 = -33; end
		1460: begin l_1 = -15;
				 l_2 = +33; end
		7283: begin l_1 = -15;
				 l_2 = -33; end
		10561: begin l_1 = +15;
				 l_2 = +34; end
		8370: begin l_1 = +15;
				 l_2 = -34; end
		5467: begin l_1 = -15;
				 l_2 = +34; end
		3276: begin l_1 = -15;
				 l_2 = -34; end
		4738: begin l_1 = +15;
				 l_2 = +35; end
		356: begin l_1 = +15;
				 l_2 = -35; end
		13481: begin l_1 = -15;
				 l_2 = +35; end
		9099: begin l_1 = -15;
				 l_2 = -35; end
		6929: begin l_1 = +15;
				 l_2 = +36; end
		12002: begin l_1 = +15;
				 l_2 = -36; end
		1835: begin l_1 = -15;
				 l_2 = +36; end
		6908: begin l_1 = -15;
				 l_2 = -36; end
		11311: begin l_1 = +15;
				 l_2 = +37; end
		7620: begin l_1 = +15;
				 l_2 = -37; end
		6217: begin l_1 = -15;
				 l_2 = +37; end
		2526: begin l_1 = -15;
				 l_2 = -37; end
		6238: begin l_1 = +15;
				 l_2 = +38; end
		12693: begin l_1 = +15;
				 l_2 = -38; end
		1144: begin l_1 = -15;
				 l_2 = +38; end
		7599: begin l_1 = -15;
				 l_2 = -38; end
		1445: begin l_1 = -16;
				 l_2 = +18; end
		12392: begin l_1 = -16;
				 l_2 = -17; end
		11633: begin l_1 = +16;
				 l_2 = +18; end
		2204: begin l_1 = -16;
				 l_2 = -18; end
		4335: begin l_1 = +16;
				 l_2 = +19; end
		5853: begin l_1 = +16;
				 l_2 = -19; end
		7984: begin l_1 = -16;
				 l_2 = +19; end
		9502: begin l_1 = -16;
				 l_2 = -19; end
		3576: begin l_1 = +16;
				 l_2 = +20; end
		6612: begin l_1 = +16;
				 l_2 = -20; end
		7225: begin l_1 = -16;
				 l_2 = +20; end
		10261: begin l_1 = -16;
				 l_2 = -20; end
		2058: begin l_1 = +16;
				 l_2 = +21; end
		8130: begin l_1 = +16;
				 l_2 = -21; end
		5707: begin l_1 = -16;
				 l_2 = +21; end
		11779: begin l_1 = -16;
				 l_2 = -21; end
		12859: begin l_1 = +16;
				 l_2 = +22; end
		11166: begin l_1 = +16;
				 l_2 = -22; end
		2671: begin l_1 = -16;
				 l_2 = +22; end
		978: begin l_1 = -16;
				 l_2 = -22; end
		6787: begin l_1 = +16;
				 l_2 = +23; end
		3401: begin l_1 = +16;
				 l_2 = -23; end
		10436: begin l_1 = -16;
				 l_2 = +23; end
		7050: begin l_1 = -16;
				 l_2 = -23; end
		8480: begin l_1 = +16;
				 l_2 = +24; end
		1708: begin l_1 = +16;
				 l_2 = -24; end
		12129: begin l_1 = -16;
				 l_2 = +24; end
		5357: begin l_1 = -16;
				 l_2 = -24; end
		11866: begin l_1 = +16;
				 l_2 = +25; end
		12159: begin l_1 = +16;
				 l_2 = -25; end
		1678: begin l_1 = -16;
				 l_2 = +25; end
		1971: begin l_1 = -16;
				 l_2 = -25; end
		4801: begin l_1 = +16;
				 l_2 = +26; end
		5387: begin l_1 = +16;
				 l_2 = -26; end
		8450: begin l_1 = -16;
				 l_2 = +26; end
		9036: begin l_1 = -16;
				 l_2 = -26; end
		4508: begin l_1 = +16;
				 l_2 = +27; end
		5680: begin l_1 = +16;
				 l_2 = -27; end
		8157: begin l_1 = -16;
				 l_2 = +27; end
		9329: begin l_1 = -16;
				 l_2 = -27; end
		3922: begin l_1 = +16;
				 l_2 = +28; end
		6266: begin l_1 = +16;
				 l_2 = -28; end
		7571: begin l_1 = -16;
				 l_2 = +28; end
		9915: begin l_1 = -16;
				 l_2 = -28; end
		2750: begin l_1 = +16;
				 l_2 = +29; end
		7438: begin l_1 = +16;
				 l_2 = -29; end
		6399: begin l_1 = -16;
				 l_2 = +29; end
		11087: begin l_1 = -16;
				 l_2 = -29; end
		406: begin l_1 = +16;
				 l_2 = +30; end
		9782: begin l_1 = +16;
				 l_2 = -30; end
		4055: begin l_1 = -16;
				 l_2 = +30; end
		13431: begin l_1 = -16;
				 l_2 = -30; end
		9555: begin l_1 = +16;
				 l_2 = +31; end
		633: begin l_1 = +16;
				 l_2 = -31; end
		13204: begin l_1 = -16;
				 l_2 = +31; end
		4282: begin l_1 = -16;
				 l_2 = -31; end
		179: begin l_1 = +16;
				 l_2 = +32; end
		10009: begin l_1 = +16;
				 l_2 = -32; end
		3828: begin l_1 = -16;
				 l_2 = +32; end
		13658: begin l_1 = -16;
				 l_2 = -32; end
		9101: begin l_1 = +16;
				 l_2 = +33; end
		1087: begin l_1 = +16;
				 l_2 = -33; end
		12750: begin l_1 = -16;
				 l_2 = +33; end
		4736: begin l_1 = -16;
				 l_2 = -33; end
		13108: begin l_1 = +16;
				 l_2 = +34; end
		10917: begin l_1 = +16;
				 l_2 = -34; end
		2920: begin l_1 = -16;
				 l_2 = +34; end
		729: begin l_1 = -16;
				 l_2 = -34; end
		7285: begin l_1 = +16;
				 l_2 = +35; end
		2903: begin l_1 = +16;
				 l_2 = -35; end
		10934: begin l_1 = -16;
				 l_2 = +35; end
		6552: begin l_1 = -16;
				 l_2 = -35; end
		9476: begin l_1 = +16;
				 l_2 = +36; end
		712: begin l_1 = +16;
				 l_2 = -36; end
		13125: begin l_1 = -16;
				 l_2 = +36; end
		4361: begin l_1 = -16;
				 l_2 = -36; end
		21: begin l_1 = +16;
				 l_2 = +37; end
		10167: begin l_1 = +16;
				 l_2 = -37; end
		3670: begin l_1 = -16;
				 l_2 = +37; end
		13816: begin l_1 = -16;
				 l_2 = -37; end
		8785: begin l_1 = +16;
				 l_2 = +38; end
		1403: begin l_1 = +16;
				 l_2 = -38; end
		12434: begin l_1 = -16;
				 l_2 = +38; end
		5052: begin l_1 = -16;
				 l_2 = -38; end
		2890: begin l_1 = -17;
				 l_2 = +19; end
		10947: begin l_1 = -17;
				 l_2 = -18; end
		9429: begin l_1 = +17;
				 l_2 = +19; end
		4408: begin l_1 = -17;
				 l_2 = -19; end
		8670: begin l_1 = +17;
				 l_2 = +20; end
		11706: begin l_1 = +17;
				 l_2 = -20; end
		2131: begin l_1 = -17;
				 l_2 = +20; end
		5167: begin l_1 = -17;
				 l_2 = -20; end
		7152: begin l_1 = +17;
				 l_2 = +21; end
		13224: begin l_1 = +17;
				 l_2 = -21; end
		613: begin l_1 = -17;
				 l_2 = +21; end
		6685: begin l_1 = -17;
				 l_2 = -21; end
		4116: begin l_1 = +17;
				 l_2 = +22; end
		2423: begin l_1 = +17;
				 l_2 = -22; end
		11414: begin l_1 = -17;
				 l_2 = +22; end
		9721: begin l_1 = -17;
				 l_2 = -22; end
		11881: begin l_1 = +17;
				 l_2 = +23; end
		8495: begin l_1 = +17;
				 l_2 = -23; end
		5342: begin l_1 = -17;
				 l_2 = +23; end
		1956: begin l_1 = -17;
				 l_2 = -23; end
		13574: begin l_1 = +17;
				 l_2 = +24; end
		6802: begin l_1 = +17;
				 l_2 = -24; end
		7035: begin l_1 = -17;
				 l_2 = +24; end
		263: begin l_1 = -17;
				 l_2 = -24; end
		3123: begin l_1 = +17;
				 l_2 = +25; end
		3416: begin l_1 = +17;
				 l_2 = -25; end
		10421: begin l_1 = -17;
				 l_2 = +25; end
		10714: begin l_1 = -17;
				 l_2 = -25; end
		9895: begin l_1 = +17;
				 l_2 = +26; end
		10481: begin l_1 = +17;
				 l_2 = -26; end
		3356: begin l_1 = -17;
				 l_2 = +26; end
		3942: begin l_1 = -17;
				 l_2 = -26; end
		9602: begin l_1 = +17;
				 l_2 = +27; end
		10774: begin l_1 = +17;
				 l_2 = -27; end
		3063: begin l_1 = -17;
				 l_2 = +27; end
		4235: begin l_1 = -17;
				 l_2 = -27; end
		9016: begin l_1 = +17;
				 l_2 = +28; end
		11360: begin l_1 = +17;
				 l_2 = -28; end
		2477: begin l_1 = -17;
				 l_2 = +28; end
		4821: begin l_1 = -17;
				 l_2 = -28; end
		7844: begin l_1 = +17;
				 l_2 = +29; end
		12532: begin l_1 = +17;
				 l_2 = -29; end
		1305: begin l_1 = -17;
				 l_2 = +29; end
		5993: begin l_1 = -17;
				 l_2 = -29; end
		5500: begin l_1 = +17;
				 l_2 = +30; end
		1039: begin l_1 = +17;
				 l_2 = -30; end
		12798: begin l_1 = -17;
				 l_2 = +30; end
		8337: begin l_1 = -17;
				 l_2 = -30; end
		812: begin l_1 = +17;
				 l_2 = +31; end
		5727: begin l_1 = +17;
				 l_2 = -31; end
		8110: begin l_1 = -17;
				 l_2 = +31; end
		13025: begin l_1 = -17;
				 l_2 = -31; end
		5273: begin l_1 = +17;
				 l_2 = +32; end
		1266: begin l_1 = +17;
				 l_2 = -32; end
		12571: begin l_1 = -17;
				 l_2 = +32; end
		8564: begin l_1 = -17;
				 l_2 = -32; end
		358: begin l_1 = +17;
				 l_2 = +33; end
		6181: begin l_1 = +17;
				 l_2 = -33; end
		7656: begin l_1 = -17;
				 l_2 = +33; end
		13479: begin l_1 = -17;
				 l_2 = -33; end
		4365: begin l_1 = +17;
				 l_2 = +34; end
		2174: begin l_1 = +17;
				 l_2 = -34; end
		11663: begin l_1 = -17;
				 l_2 = +34; end
		9472: begin l_1 = -17;
				 l_2 = -34; end
		12379: begin l_1 = +17;
				 l_2 = +35; end
		7997: begin l_1 = +17;
				 l_2 = -35; end
		5840: begin l_1 = -17;
				 l_2 = +35; end
		1458: begin l_1 = -17;
				 l_2 = -35; end
		733: begin l_1 = +17;
				 l_2 = +36; end
		5806: begin l_1 = +17;
				 l_2 = -36; end
		8031: begin l_1 = -17;
				 l_2 = +36; end
		13104: begin l_1 = -17;
				 l_2 = -36; end
		5115: begin l_1 = +17;
				 l_2 = +37; end
		1424: begin l_1 = +17;
				 l_2 = -37; end
		12413: begin l_1 = -17;
				 l_2 = +37; end
		8722: begin l_1 = -17;
				 l_2 = -37; end
		42: begin l_1 = +17;
				 l_2 = +38; end
		6497: begin l_1 = +17;
				 l_2 = -38; end
		7340: begin l_1 = -17;
				 l_2 = +38; end
		13795: begin l_1 = -17;
				 l_2 = -38; end
		5780: begin l_1 = -18;
				 l_2 = +20; end
		8057: begin l_1 = -18;
				 l_2 = -19; end
		5021: begin l_1 = +18;
				 l_2 = +20; end
		8816: begin l_1 = -18;
				 l_2 = -20; end
		3503: begin l_1 = +18;
				 l_2 = +21; end
		9575: begin l_1 = +18;
				 l_2 = -21; end
		4262: begin l_1 = -18;
				 l_2 = +21; end
		10334: begin l_1 = -18;
				 l_2 = -21; end
		467: begin l_1 = +18;
				 l_2 = +22; end
		12611: begin l_1 = +18;
				 l_2 = -22; end
		1226: begin l_1 = -18;
				 l_2 = +22; end
		13370: begin l_1 = -18;
				 l_2 = -22; end
		8232: begin l_1 = +18;
				 l_2 = +23; end
		4846: begin l_1 = +18;
				 l_2 = -23; end
		8991: begin l_1 = -18;
				 l_2 = +23; end
		5605: begin l_1 = -18;
				 l_2 = -23; end
		9925: begin l_1 = +18;
				 l_2 = +24; end
		3153: begin l_1 = +18;
				 l_2 = -24; end
		10684: begin l_1 = -18;
				 l_2 = +24; end
		3912: begin l_1 = -18;
				 l_2 = -24; end
		13311: begin l_1 = +18;
				 l_2 = +25; end
		13604: begin l_1 = +18;
				 l_2 = -25; end
		233: begin l_1 = -18;
				 l_2 = +25; end
		526: begin l_1 = -18;
				 l_2 = -25; end
		6246: begin l_1 = +18;
				 l_2 = +26; end
		6832: begin l_1 = +18;
				 l_2 = -26; end
		7005: begin l_1 = -18;
				 l_2 = +26; end
		7591: begin l_1 = -18;
				 l_2 = -26; end
		5953: begin l_1 = +18;
				 l_2 = +27; end
		7125: begin l_1 = +18;
				 l_2 = -27; end
		6712: begin l_1 = -18;
				 l_2 = +27; end
		7884: begin l_1 = -18;
				 l_2 = -27; end
		5367: begin l_1 = +18;
				 l_2 = +28; end
		7711: begin l_1 = +18;
				 l_2 = -28; end
		6126: begin l_1 = -18;
				 l_2 = +28; end
		8470: begin l_1 = -18;
				 l_2 = -28; end
		4195: begin l_1 = +18;
				 l_2 = +29; end
		8883: begin l_1 = +18;
				 l_2 = -29; end
		4954: begin l_1 = -18;
				 l_2 = +29; end
		9642: begin l_1 = -18;
				 l_2 = -29; end
		1851: begin l_1 = +18;
				 l_2 = +30; end
		11227: begin l_1 = +18;
				 l_2 = -30; end
		2610: begin l_1 = -18;
				 l_2 = +30; end
		11986: begin l_1 = -18;
				 l_2 = -30; end
		11000: begin l_1 = +18;
				 l_2 = +31; end
		2078: begin l_1 = +18;
				 l_2 = -31; end
		11759: begin l_1 = -18;
				 l_2 = +31; end
		2837: begin l_1 = -18;
				 l_2 = -31; end
		1624: begin l_1 = +18;
				 l_2 = +32; end
		11454: begin l_1 = +18;
				 l_2 = -32; end
		2383: begin l_1 = -18;
				 l_2 = +32; end
		12213: begin l_1 = -18;
				 l_2 = -32; end
		10546: begin l_1 = +18;
				 l_2 = +33; end
		2532: begin l_1 = +18;
				 l_2 = -33; end
		11305: begin l_1 = -18;
				 l_2 = +33; end
		3291: begin l_1 = -18;
				 l_2 = -33; end
		716: begin l_1 = +18;
				 l_2 = +34; end
		12362: begin l_1 = +18;
				 l_2 = -34; end
		1475: begin l_1 = -18;
				 l_2 = +34; end
		13121: begin l_1 = -18;
				 l_2 = -34; end
		8730: begin l_1 = +18;
				 l_2 = +35; end
		4348: begin l_1 = +18;
				 l_2 = -35; end
		9489: begin l_1 = -18;
				 l_2 = +35; end
		5107: begin l_1 = -18;
				 l_2 = -35; end
		10921: begin l_1 = +18;
				 l_2 = +36; end
		2157: begin l_1 = +18;
				 l_2 = -36; end
		11680: begin l_1 = -18;
				 l_2 = +36; end
		2916: begin l_1 = -18;
				 l_2 = -36; end
		1466: begin l_1 = +18;
				 l_2 = +37; end
		11612: begin l_1 = +18;
				 l_2 = -37; end
		2225: begin l_1 = -18;
				 l_2 = +37; end
		12371: begin l_1 = -18;
				 l_2 = -37; end
		10230: begin l_1 = +18;
				 l_2 = +38; end
		2848: begin l_1 = +18;
				 l_2 = -38; end
		10989: begin l_1 = -18;
				 l_2 = +38; end
		3607: begin l_1 = -18;
				 l_2 = -38; end
		11560: begin l_1 = -19;
				 l_2 = +21; end
		2277: begin l_1 = -19;
				 l_2 = -20; end
		10042: begin l_1 = +19;
				 l_2 = +21; end
		3795: begin l_1 = -19;
				 l_2 = -21; end
		7006: begin l_1 = +19;
				 l_2 = +22; end
		5313: begin l_1 = +19;
				 l_2 = -22; end
		8524: begin l_1 = -19;
				 l_2 = +22; end
		6831: begin l_1 = -19;
				 l_2 = -22; end
		934: begin l_1 = +19;
				 l_2 = +23; end
		11385: begin l_1 = +19;
				 l_2 = -23; end
		2452: begin l_1 = -19;
				 l_2 = +23; end
		12903: begin l_1 = -19;
				 l_2 = -23; end
		2627: begin l_1 = +19;
				 l_2 = +24; end
		9692: begin l_1 = +19;
				 l_2 = -24; end
		4145: begin l_1 = -19;
				 l_2 = +24; end
		11210: begin l_1 = -19;
				 l_2 = -24; end
		6013: begin l_1 = +19;
				 l_2 = +25; end
		6306: begin l_1 = +19;
				 l_2 = -25; end
		7531: begin l_1 = -19;
				 l_2 = +25; end
		7824: begin l_1 = -19;
				 l_2 = -25; end
		12785: begin l_1 = +19;
				 l_2 = +26; end
		13371: begin l_1 = +19;
				 l_2 = -26; end
		466: begin l_1 = -19;
				 l_2 = +26; end
		1052: begin l_1 = -19;
				 l_2 = -26; end
		12492: begin l_1 = +19;
				 l_2 = +27; end
		13664: begin l_1 = +19;
				 l_2 = -27; end
		173: begin l_1 = -19;
				 l_2 = +27; end
		1345: begin l_1 = -19;
				 l_2 = -27; end
		11906: begin l_1 = +19;
				 l_2 = +28; end
		413: begin l_1 = +19;
				 l_2 = -28; end
		13424: begin l_1 = -19;
				 l_2 = +28; end
		1931: begin l_1 = -19;
				 l_2 = -28; end
		10734: begin l_1 = +19;
				 l_2 = +29; end
		1585: begin l_1 = +19;
				 l_2 = -29; end
		12252: begin l_1 = -19;
				 l_2 = +29; end
		3103: begin l_1 = -19;
				 l_2 = -29; end
		8390: begin l_1 = +19;
				 l_2 = +30; end
		3929: begin l_1 = +19;
				 l_2 = -30; end
		9908: begin l_1 = -19;
				 l_2 = +30; end
		5447: begin l_1 = -19;
				 l_2 = -30; end
		3702: begin l_1 = +19;
				 l_2 = +31; end
		8617: begin l_1 = +19;
				 l_2 = -31; end
		5220: begin l_1 = -19;
				 l_2 = +31; end
		10135: begin l_1 = -19;
				 l_2 = -31; end
		8163: begin l_1 = +19;
				 l_2 = +32; end
		4156: begin l_1 = +19;
				 l_2 = -32; end
		9681: begin l_1 = -19;
				 l_2 = +32; end
		5674: begin l_1 = -19;
				 l_2 = -32; end
		3248: begin l_1 = +19;
				 l_2 = +33; end
		9071: begin l_1 = +19;
				 l_2 = -33; end
		4766: begin l_1 = -19;
				 l_2 = +33; end
		10589: begin l_1 = -19;
				 l_2 = -33; end
		7255: begin l_1 = +19;
				 l_2 = +34; end
		5064: begin l_1 = +19;
				 l_2 = -34; end
		8773: begin l_1 = -19;
				 l_2 = +34; end
		6582: begin l_1 = -19;
				 l_2 = -34; end
		1432: begin l_1 = +19;
				 l_2 = +35; end
		10887: begin l_1 = +19;
				 l_2 = -35; end
		2950: begin l_1 = -19;
				 l_2 = +35; end
		12405: begin l_1 = -19;
				 l_2 = -35; end
		3623: begin l_1 = +19;
				 l_2 = +36; end
		8696: begin l_1 = +19;
				 l_2 = -36; end
		5141: begin l_1 = -19;
				 l_2 = +36; end
		10214: begin l_1 = -19;
				 l_2 = -36; end
		8005: begin l_1 = +19;
				 l_2 = +37; end
		4314: begin l_1 = +19;
				 l_2 = -37; end
		9523: begin l_1 = -19;
				 l_2 = +37; end
		5832: begin l_1 = -19;
				 l_2 = -37; end
		2932: begin l_1 = +19;
				 l_2 = +38; end
		9387: begin l_1 = +19;
				 l_2 = -38; end
		4450: begin l_1 = -19;
				 l_2 = +38; end
		10905: begin l_1 = -19;
				 l_2 = -38; end
		9283: begin l_1 = -20;
				 l_2 = +22; end
		4554: begin l_1 = -20;
				 l_2 = -21; end
		6247: begin l_1 = +20;
				 l_2 = +22; end
		7590: begin l_1 = -20;
				 l_2 = -22; end
		175: begin l_1 = +20;
				 l_2 = +23; end
		10626: begin l_1 = +20;
				 l_2 = -23; end
		3211: begin l_1 = -20;
				 l_2 = +23; end
		13662: begin l_1 = -20;
				 l_2 = -23; end
		1868: begin l_1 = +20;
				 l_2 = +24; end
		8933: begin l_1 = +20;
				 l_2 = -24; end
		4904: begin l_1 = -20;
				 l_2 = +24; end
		11969: begin l_1 = -20;
				 l_2 = -24; end
		5254: begin l_1 = +20;
				 l_2 = +25; end
		5547: begin l_1 = +20;
				 l_2 = -25; end
		8290: begin l_1 = -20;
				 l_2 = +25; end
		8583: begin l_1 = -20;
				 l_2 = -25; end
		12026: begin l_1 = +20;
				 l_2 = +26; end
		12612: begin l_1 = +20;
				 l_2 = -26; end
		1225: begin l_1 = -20;
				 l_2 = +26; end
		1811: begin l_1 = -20;
				 l_2 = -26; end
		11733: begin l_1 = +20;
				 l_2 = +27; end
		12905: begin l_1 = +20;
				 l_2 = -27; end
		932: begin l_1 = -20;
				 l_2 = +27; end
		2104: begin l_1 = -20;
				 l_2 = -27; end
		11147: begin l_1 = +20;
				 l_2 = +28; end
		13491: begin l_1 = +20;
				 l_2 = -28; end
		346: begin l_1 = -20;
				 l_2 = +28; end
		2690: begin l_1 = -20;
				 l_2 = -28; end
		9975: begin l_1 = +20;
				 l_2 = +29; end
		826: begin l_1 = +20;
				 l_2 = -29; end
		13011: begin l_1 = -20;
				 l_2 = +29; end
		3862: begin l_1 = -20;
				 l_2 = -29; end
		7631: begin l_1 = +20;
				 l_2 = +30; end
		3170: begin l_1 = +20;
				 l_2 = -30; end
		10667: begin l_1 = -20;
				 l_2 = +30; end
		6206: begin l_1 = -20;
				 l_2 = -30; end
		2943: begin l_1 = +20;
				 l_2 = +31; end
		7858: begin l_1 = +20;
				 l_2 = -31; end
		5979: begin l_1 = -20;
				 l_2 = +31; end
		10894: begin l_1 = -20;
				 l_2 = -31; end
		7404: begin l_1 = +20;
				 l_2 = +32; end
		3397: begin l_1 = +20;
				 l_2 = -32; end
		10440: begin l_1 = -20;
				 l_2 = +32; end
		6433: begin l_1 = -20;
				 l_2 = -32; end
		2489: begin l_1 = +20;
				 l_2 = +33; end
		8312: begin l_1 = +20;
				 l_2 = -33; end
		5525: begin l_1 = -20;
				 l_2 = +33; end
		11348: begin l_1 = -20;
				 l_2 = -33; end
		6496: begin l_1 = +20;
				 l_2 = +34; end
		4305: begin l_1 = +20;
				 l_2 = -34; end
		9532: begin l_1 = -20;
				 l_2 = +34; end
		7341: begin l_1 = -20;
				 l_2 = -34; end
		673: begin l_1 = +20;
				 l_2 = +35; end
		10128: begin l_1 = +20;
				 l_2 = -35; end
		3709: begin l_1 = -20;
				 l_2 = +35; end
		13164: begin l_1 = -20;
				 l_2 = -35; end
		2864: begin l_1 = +20;
				 l_2 = +36; end
		7937: begin l_1 = +20;
				 l_2 = -36; end
		5900: begin l_1 = -20;
				 l_2 = +36; end
		10973: begin l_1 = -20;
				 l_2 = -36; end
		7246: begin l_1 = +20;
				 l_2 = +37; end
		3555: begin l_1 = +20;
				 l_2 = -37; end
		10282: begin l_1 = -20;
				 l_2 = +37; end
		6591: begin l_1 = -20;
				 l_2 = -37; end
		2173: begin l_1 = +20;
				 l_2 = +38; end
		8628: begin l_1 = +20;
				 l_2 = -38; end
		5209: begin l_1 = -20;
				 l_2 = +38; end
		11664: begin l_1 = -20;
				 l_2 = -38; end
		4729: begin l_1 = -21;
				 l_2 = +23; end
		9108: begin l_1 = -21;
				 l_2 = -22; end
		12494: begin l_1 = +21;
				 l_2 = +23; end
		1343: begin l_1 = -21;
				 l_2 = -23; end
		350: begin l_1 = +21;
				 l_2 = +24; end
		7415: begin l_1 = +21;
				 l_2 = -24; end
		6422: begin l_1 = -21;
				 l_2 = +24; end
		13487: begin l_1 = -21;
				 l_2 = -24; end
		3736: begin l_1 = +21;
				 l_2 = +25; end
		4029: begin l_1 = +21;
				 l_2 = -25; end
		9808: begin l_1 = -21;
				 l_2 = +25; end
		10101: begin l_1 = -21;
				 l_2 = -25; end
		10508: begin l_1 = +21;
				 l_2 = +26; end
		11094: begin l_1 = +21;
				 l_2 = -26; end
		2743: begin l_1 = -21;
				 l_2 = +26; end
		3329: begin l_1 = -21;
				 l_2 = -26; end
		10215: begin l_1 = +21;
				 l_2 = +27; end
		11387: begin l_1 = +21;
				 l_2 = -27; end
		2450: begin l_1 = -21;
				 l_2 = +27; end
		3622: begin l_1 = -21;
				 l_2 = -27; end
		9629: begin l_1 = +21;
				 l_2 = +28; end
		11973: begin l_1 = +21;
				 l_2 = -28; end
		1864: begin l_1 = -21;
				 l_2 = +28; end
		4208: begin l_1 = -21;
				 l_2 = -28; end
		8457: begin l_1 = +21;
				 l_2 = +29; end
		13145: begin l_1 = +21;
				 l_2 = -29; end
		692: begin l_1 = -21;
				 l_2 = +29; end
		5380: begin l_1 = -21;
				 l_2 = -29; end
		6113: begin l_1 = +21;
				 l_2 = +30; end
		1652: begin l_1 = +21;
				 l_2 = -30; end
		12185: begin l_1 = -21;
				 l_2 = +30; end
		7724: begin l_1 = -21;
				 l_2 = -30; end
		1425: begin l_1 = +21;
				 l_2 = +31; end
		6340: begin l_1 = +21;
				 l_2 = -31; end
		7497: begin l_1 = -21;
				 l_2 = +31; end
		12412: begin l_1 = -21;
				 l_2 = -31; end
		5886: begin l_1 = +21;
				 l_2 = +32; end
		1879: begin l_1 = +21;
				 l_2 = -32; end
		11958: begin l_1 = -21;
				 l_2 = +32; end
		7951: begin l_1 = -21;
				 l_2 = -32; end
		971: begin l_1 = +21;
				 l_2 = +33; end
		6794: begin l_1 = +21;
				 l_2 = -33; end
		7043: begin l_1 = -21;
				 l_2 = +33; end
		12866: begin l_1 = -21;
				 l_2 = -33; end
		4978: begin l_1 = +21;
				 l_2 = +34; end
		2787: begin l_1 = +21;
				 l_2 = -34; end
		11050: begin l_1 = -21;
				 l_2 = +34; end
		8859: begin l_1 = -21;
				 l_2 = -34; end
		12992: begin l_1 = +21;
				 l_2 = +35; end
		8610: begin l_1 = +21;
				 l_2 = -35; end
		5227: begin l_1 = -21;
				 l_2 = +35; end
		845: begin l_1 = -21;
				 l_2 = -35; end
		1346: begin l_1 = +21;
				 l_2 = +36; end
		6419: begin l_1 = +21;
				 l_2 = -36; end
		7418: begin l_1 = -21;
				 l_2 = +36; end
		12491: begin l_1 = -21;
				 l_2 = -36; end
		5728: begin l_1 = +21;
				 l_2 = +37; end
		2037: begin l_1 = +21;
				 l_2 = -37; end
		11800: begin l_1 = -21;
				 l_2 = +37; end
		8109: begin l_1 = -21;
				 l_2 = -37; end
		655: begin l_1 = +21;
				 l_2 = +38; end
		7110: begin l_1 = +21;
				 l_2 = -38; end
		6727: begin l_1 = -21;
				 l_2 = +38; end
		13182: begin l_1 = -21;
				 l_2 = -38; end
		9458: begin l_1 = -22;
				 l_2 = +24; end
		4379: begin l_1 = -22;
				 l_2 = -23; end
		11151: begin l_1 = +22;
				 l_2 = +24; end
		2686: begin l_1 = -22;
				 l_2 = -24; end
		700: begin l_1 = +22;
				 l_2 = +25; end
		993: begin l_1 = +22;
				 l_2 = -25; end
		12844: begin l_1 = -22;
				 l_2 = +25; end
		13137: begin l_1 = -22;
				 l_2 = -25; end
		7472: begin l_1 = +22;
				 l_2 = +26; end
		8058: begin l_1 = +22;
				 l_2 = -26; end
		5779: begin l_1 = -22;
				 l_2 = +26; end
		6365: begin l_1 = -22;
				 l_2 = -26; end
		7179: begin l_1 = +22;
				 l_2 = +27; end
		8351: begin l_1 = +22;
				 l_2 = -27; end
		5486: begin l_1 = -22;
				 l_2 = +27; end
		6658: begin l_1 = -22;
				 l_2 = -27; end
		6593: begin l_1 = +22;
				 l_2 = +28; end
		8937: begin l_1 = +22;
				 l_2 = -28; end
		4900: begin l_1 = -22;
				 l_2 = +28; end
		7244: begin l_1 = -22;
				 l_2 = -28; end
		5421: begin l_1 = +22;
				 l_2 = +29; end
		10109: begin l_1 = +22;
				 l_2 = -29; end
		3728: begin l_1 = -22;
				 l_2 = +29; end
		8416: begin l_1 = -22;
				 l_2 = -29; end
		3077: begin l_1 = +22;
				 l_2 = +30; end
		12453: begin l_1 = +22;
				 l_2 = -30; end
		1384: begin l_1 = -22;
				 l_2 = +30; end
		10760: begin l_1 = -22;
				 l_2 = -30; end
		12226: begin l_1 = +22;
				 l_2 = +31; end
		3304: begin l_1 = +22;
				 l_2 = -31; end
		10533: begin l_1 = -22;
				 l_2 = +31; end
		1611: begin l_1 = -22;
				 l_2 = -31; end
		2850: begin l_1 = +22;
				 l_2 = +32; end
		12680: begin l_1 = +22;
				 l_2 = -32; end
		1157: begin l_1 = -22;
				 l_2 = +32; end
		10987: begin l_1 = -22;
				 l_2 = -32; end
		11772: begin l_1 = +22;
				 l_2 = +33; end
		3758: begin l_1 = +22;
				 l_2 = -33; end
		10079: begin l_1 = -22;
				 l_2 = +33; end
		2065: begin l_1 = -22;
				 l_2 = -33; end
		1942: begin l_1 = +22;
				 l_2 = +34; end
		13588: begin l_1 = +22;
				 l_2 = -34; end
		249: begin l_1 = -22;
				 l_2 = +34; end
		11895: begin l_1 = -22;
				 l_2 = -34; end
		9956: begin l_1 = +22;
				 l_2 = +35; end
		5574: begin l_1 = +22;
				 l_2 = -35; end
		8263: begin l_1 = -22;
				 l_2 = +35; end
		3881: begin l_1 = -22;
				 l_2 = -35; end
		12147: begin l_1 = +22;
				 l_2 = +36; end
		3383: begin l_1 = +22;
				 l_2 = -36; end
		10454: begin l_1 = -22;
				 l_2 = +36; end
		1690: begin l_1 = -22;
				 l_2 = -36; end
		2692: begin l_1 = +22;
				 l_2 = +37; end
		12838: begin l_1 = +22;
				 l_2 = -37; end
		999: begin l_1 = -22;
				 l_2 = +37; end
		11145: begin l_1 = -22;
				 l_2 = -37; end
		11456: begin l_1 = +22;
				 l_2 = +38; end
		4074: begin l_1 = +22;
				 l_2 = -38; end
		9763: begin l_1 = -22;
				 l_2 = +38; end
		2381: begin l_1 = -22;
				 l_2 = -38; end
		5079: begin l_1 = -23;
				 l_2 = +25; end
		8758: begin l_1 = -23;
				 l_2 = -24; end
		8465: begin l_1 = +23;
				 l_2 = +25; end
		5372: begin l_1 = -23;
				 l_2 = -25; end
		1400: begin l_1 = +23;
				 l_2 = +26; end
		1986: begin l_1 = +23;
				 l_2 = -26; end
		11851: begin l_1 = -23;
				 l_2 = +26; end
		12437: begin l_1 = -23;
				 l_2 = -26; end
		1107: begin l_1 = +23;
				 l_2 = +27; end
		2279: begin l_1 = +23;
				 l_2 = -27; end
		11558: begin l_1 = -23;
				 l_2 = +27; end
		12730: begin l_1 = -23;
				 l_2 = -27; end
		521: begin l_1 = +23;
				 l_2 = +28; end
		2865: begin l_1 = +23;
				 l_2 = -28; end
		10972: begin l_1 = -23;
				 l_2 = +28; end
		13316: begin l_1 = -23;
				 l_2 = -28; end
		13186: begin l_1 = +23;
				 l_2 = +29; end
		4037: begin l_1 = +23;
				 l_2 = -29; end
		9800: begin l_1 = -23;
				 l_2 = +29; end
		651: begin l_1 = -23;
				 l_2 = -29; end
		10842: begin l_1 = +23;
				 l_2 = +30; end
		6381: begin l_1 = +23;
				 l_2 = -30; end
		7456: begin l_1 = -23;
				 l_2 = +30; end
		2995: begin l_1 = -23;
				 l_2 = -30; end
		6154: begin l_1 = +23;
				 l_2 = +31; end
		11069: begin l_1 = +23;
				 l_2 = -31; end
		2768: begin l_1 = -23;
				 l_2 = +31; end
		7683: begin l_1 = -23;
				 l_2 = -31; end
		10615: begin l_1 = +23;
				 l_2 = +32; end
		6608: begin l_1 = +23;
				 l_2 = -32; end
		7229: begin l_1 = -23;
				 l_2 = +32; end
		3222: begin l_1 = -23;
				 l_2 = -32; end
		5700: begin l_1 = +23;
				 l_2 = +33; end
		11523: begin l_1 = +23;
				 l_2 = -33; end
		2314: begin l_1 = -23;
				 l_2 = +33; end
		8137: begin l_1 = -23;
				 l_2 = -33; end
		9707: begin l_1 = +23;
				 l_2 = +34; end
		7516: begin l_1 = +23;
				 l_2 = -34; end
		6321: begin l_1 = -23;
				 l_2 = +34; end
		4130: begin l_1 = -23;
				 l_2 = -34; end
		3884: begin l_1 = +23;
				 l_2 = +35; end
		13339: begin l_1 = +23;
				 l_2 = -35; end
		498: begin l_1 = -23;
				 l_2 = +35; end
		9953: begin l_1 = -23;
				 l_2 = -35; end
		6075: begin l_1 = +23;
				 l_2 = +36; end
		11148: begin l_1 = +23;
				 l_2 = -36; end
		2689: begin l_1 = -23;
				 l_2 = +36; end
		7762: begin l_1 = -23;
				 l_2 = -36; end
		10457: begin l_1 = +23;
				 l_2 = +37; end
		6766: begin l_1 = +23;
				 l_2 = -37; end
		7071: begin l_1 = -23;
				 l_2 = +37; end
		3380: begin l_1 = -23;
				 l_2 = -37; end
		5384: begin l_1 = +23;
				 l_2 = +38; end
		11839: begin l_1 = +23;
				 l_2 = -38; end
		1998: begin l_1 = -23;
				 l_2 = +38; end
		8453: begin l_1 = -23;
				 l_2 = -38; end
		10158: begin l_1 = -24;
				 l_2 = +26; end
		3679: begin l_1 = -24;
				 l_2 = -25; end
		3093: begin l_1 = +24;
				 l_2 = +26; end
		10744: begin l_1 = -24;
				 l_2 = -26; end
		2800: begin l_1 = +24;
				 l_2 = +27; end
		3972: begin l_1 = +24;
				 l_2 = -27; end
		9865: begin l_1 = -24;
				 l_2 = +27; end
		11037: begin l_1 = -24;
				 l_2 = -27; end
		2214: begin l_1 = +24;
				 l_2 = +28; end
		4558: begin l_1 = +24;
				 l_2 = -28; end
		9279: begin l_1 = -24;
				 l_2 = +28; end
		11623: begin l_1 = -24;
				 l_2 = -28; end
		1042: begin l_1 = +24;
				 l_2 = +29; end
		5730: begin l_1 = +24;
				 l_2 = -29; end
		8107: begin l_1 = -24;
				 l_2 = +29; end
		12795: begin l_1 = -24;
				 l_2 = -29; end
		12535: begin l_1 = +24;
				 l_2 = +30; end
		8074: begin l_1 = +24;
				 l_2 = -30; end
		5763: begin l_1 = -24;
				 l_2 = +30; end
		1302: begin l_1 = -24;
				 l_2 = -30; end
		7847: begin l_1 = +24;
				 l_2 = +31; end
		12762: begin l_1 = +24;
				 l_2 = -31; end
		1075: begin l_1 = -24;
				 l_2 = +31; end
		5990: begin l_1 = -24;
				 l_2 = -31; end
		12308: begin l_1 = +24;
				 l_2 = +32; end
		8301: begin l_1 = +24;
				 l_2 = -32; end
		5536: begin l_1 = -24;
				 l_2 = +32; end
		1529: begin l_1 = -24;
				 l_2 = -32; end
		7393: begin l_1 = +24;
				 l_2 = +33; end
		13216: begin l_1 = +24;
				 l_2 = -33; end
		621: begin l_1 = -24;
				 l_2 = +33; end
		6444: begin l_1 = -24;
				 l_2 = -33; end
		11400: begin l_1 = +24;
				 l_2 = +34; end
		9209: begin l_1 = +24;
				 l_2 = -34; end
		4628: begin l_1 = -24;
				 l_2 = +34; end
		2437: begin l_1 = -24;
				 l_2 = -34; end
		5577: begin l_1 = +24;
				 l_2 = +35; end
		1195: begin l_1 = +24;
				 l_2 = -35; end
		12642: begin l_1 = -24;
				 l_2 = +35; end
		8260: begin l_1 = -24;
				 l_2 = -35; end
		7768: begin l_1 = +24;
				 l_2 = +36; end
		12841: begin l_1 = +24;
				 l_2 = -36; end
		996: begin l_1 = -24;
				 l_2 = +36; end
		6069: begin l_1 = -24;
				 l_2 = -36; end
		12150: begin l_1 = +24;
				 l_2 = +37; end
		8459: begin l_1 = +24;
				 l_2 = -37; end
		5378: begin l_1 = -24;
				 l_2 = +37; end
		1687: begin l_1 = -24;
				 l_2 = -37; end
		7077: begin l_1 = +24;
				 l_2 = +38; end
		13532: begin l_1 = +24;
				 l_2 = -38; end
		305: begin l_1 = -24;
				 l_2 = +38; end
		6760: begin l_1 = -24;
				 l_2 = -38; end
		6479: begin l_1 = -25;
				 l_2 = +27; end
		7358: begin l_1 = -25;
				 l_2 = -26; end
		6186: begin l_1 = +25;
				 l_2 = +27; end
		7651: begin l_1 = -25;
				 l_2 = -27; end
		5600: begin l_1 = +25;
				 l_2 = +28; end
		7944: begin l_1 = +25;
				 l_2 = -28; end
		5893: begin l_1 = -25;
				 l_2 = +28; end
		8237: begin l_1 = -25;
				 l_2 = -28; end
		4428: begin l_1 = +25;
				 l_2 = +29; end
		9116: begin l_1 = +25;
				 l_2 = -29; end
		4721: begin l_1 = -25;
				 l_2 = +29; end
		9409: begin l_1 = -25;
				 l_2 = -29; end
		2084: begin l_1 = +25;
				 l_2 = +30; end
		11460: begin l_1 = +25;
				 l_2 = -30; end
		2377: begin l_1 = -25;
				 l_2 = +30; end
		11753: begin l_1 = -25;
				 l_2 = -30; end
		11233: begin l_1 = +25;
				 l_2 = +31; end
		2311: begin l_1 = +25;
				 l_2 = -31; end
		11526: begin l_1 = -25;
				 l_2 = +31; end
		2604: begin l_1 = -25;
				 l_2 = -31; end
		1857: begin l_1 = +25;
				 l_2 = +32; end
		11687: begin l_1 = +25;
				 l_2 = -32; end
		2150: begin l_1 = -25;
				 l_2 = +32; end
		11980: begin l_1 = -25;
				 l_2 = -32; end
		10779: begin l_1 = +25;
				 l_2 = +33; end
		2765: begin l_1 = +25;
				 l_2 = -33; end
		11072: begin l_1 = -25;
				 l_2 = +33; end
		3058: begin l_1 = -25;
				 l_2 = -33; end
		949: begin l_1 = +25;
				 l_2 = +34; end
		12595: begin l_1 = +25;
				 l_2 = -34; end
		1242: begin l_1 = -25;
				 l_2 = +34; end
		12888: begin l_1 = -25;
				 l_2 = -34; end
		8963: begin l_1 = +25;
				 l_2 = +35; end
		4581: begin l_1 = +25;
				 l_2 = -35; end
		9256: begin l_1 = -25;
				 l_2 = +35; end
		4874: begin l_1 = -25;
				 l_2 = -35; end
		11154: begin l_1 = +25;
				 l_2 = +36; end
		2390: begin l_1 = +25;
				 l_2 = -36; end
		11447: begin l_1 = -25;
				 l_2 = +36; end
		2683: begin l_1 = -25;
				 l_2 = -36; end
		1699: begin l_1 = +25;
				 l_2 = +37; end
		11845: begin l_1 = +25;
				 l_2 = -37; end
		1992: begin l_1 = -25;
				 l_2 = +37; end
		12138: begin l_1 = -25;
				 l_2 = -37; end
		10463: begin l_1 = +25;
				 l_2 = +38; end
		3081: begin l_1 = +25;
				 l_2 = -38; end
		10756: begin l_1 = -25;
				 l_2 = +38; end
		3374: begin l_1 = -25;
				 l_2 = -38; end
		12958: begin l_1 = -26;
				 l_2 = +28; end
		879: begin l_1 = -26;
				 l_2 = -27; end
		12372: begin l_1 = +26;
				 l_2 = +28; end
		1465: begin l_1 = -26;
				 l_2 = -28; end
		11200: begin l_1 = +26;
				 l_2 = +29; end
		2051: begin l_1 = +26;
				 l_2 = -29; end
		11786: begin l_1 = -26;
				 l_2 = +29; end
		2637: begin l_1 = -26;
				 l_2 = -29; end
		8856: begin l_1 = +26;
				 l_2 = +30; end
		4395: begin l_1 = +26;
				 l_2 = -30; end
		9442: begin l_1 = -26;
				 l_2 = +30; end
		4981: begin l_1 = -26;
				 l_2 = -30; end
		4168: begin l_1 = +26;
				 l_2 = +31; end
		9083: begin l_1 = +26;
				 l_2 = -31; end
		4754: begin l_1 = -26;
				 l_2 = +31; end
		9669: begin l_1 = -26;
				 l_2 = -31; end
		8629: begin l_1 = +26;
				 l_2 = +32; end
		4622: begin l_1 = +26;
				 l_2 = -32; end
		9215: begin l_1 = -26;
				 l_2 = +32; end
		5208: begin l_1 = -26;
				 l_2 = -32; end
		3714: begin l_1 = +26;
				 l_2 = +33; end
		9537: begin l_1 = +26;
				 l_2 = -33; end
		4300: begin l_1 = -26;
				 l_2 = +33; end
		10123: begin l_1 = -26;
				 l_2 = -33; end
		7721: begin l_1 = +26;
				 l_2 = +34; end
		5530: begin l_1 = +26;
				 l_2 = -34; end
		8307: begin l_1 = -26;
				 l_2 = +34; end
		6116: begin l_1 = -26;
				 l_2 = -34; end
		1898: begin l_1 = +26;
				 l_2 = +35; end
		11353: begin l_1 = +26;
				 l_2 = -35; end
		2484: begin l_1 = -26;
				 l_2 = +35; end
		11939: begin l_1 = -26;
				 l_2 = -35; end
		4089: begin l_1 = +26;
				 l_2 = +36; end
		9162: begin l_1 = +26;
				 l_2 = -36; end
		4675: begin l_1 = -26;
				 l_2 = +36; end
		9748: begin l_1 = -26;
				 l_2 = -36; end
		8471: begin l_1 = +26;
				 l_2 = +37; end
		4780: begin l_1 = +26;
				 l_2 = -37; end
		9057: begin l_1 = -26;
				 l_2 = +37; end
		5366: begin l_1 = -26;
				 l_2 = -37; end
		3398: begin l_1 = +26;
				 l_2 = +38; end
		9853: begin l_1 = +26;
				 l_2 = -38; end
		3984: begin l_1 = -26;
				 l_2 = +38; end
		10439: begin l_1 = -26;
				 l_2 = -38; end
		12079: begin l_1 = -27;
				 l_2 = +29; end
		1758: begin l_1 = -27;
				 l_2 = -28; end
		10907: begin l_1 = +27;
				 l_2 = +29; end
		2930: begin l_1 = -27;
				 l_2 = -29; end
		8563: begin l_1 = +27;
				 l_2 = +30; end
		4102: begin l_1 = +27;
				 l_2 = -30; end
		9735: begin l_1 = -27;
				 l_2 = +30; end
		5274: begin l_1 = -27;
				 l_2 = -30; end
		3875: begin l_1 = +27;
				 l_2 = +31; end
		8790: begin l_1 = +27;
				 l_2 = -31; end
		5047: begin l_1 = -27;
				 l_2 = +31; end
		9962: begin l_1 = -27;
				 l_2 = -31; end
		8336: begin l_1 = +27;
				 l_2 = +32; end
		4329: begin l_1 = +27;
				 l_2 = -32; end
		9508: begin l_1 = -27;
				 l_2 = +32; end
		5501: begin l_1 = -27;
				 l_2 = -32; end
		3421: begin l_1 = +27;
				 l_2 = +33; end
		9244: begin l_1 = +27;
				 l_2 = -33; end
		4593: begin l_1 = -27;
				 l_2 = +33; end
		10416: begin l_1 = -27;
				 l_2 = -33; end
		7428: begin l_1 = +27;
				 l_2 = +34; end
		5237: begin l_1 = +27;
				 l_2 = -34; end
		8600: begin l_1 = -27;
				 l_2 = +34; end
		6409: begin l_1 = -27;
				 l_2 = -34; end
		1605: begin l_1 = +27;
				 l_2 = +35; end
		11060: begin l_1 = +27;
				 l_2 = -35; end
		2777: begin l_1 = -27;
				 l_2 = +35; end
		12232: begin l_1 = -27;
				 l_2 = -35; end
		3796: begin l_1 = +27;
				 l_2 = +36; end
		8869: begin l_1 = +27;
				 l_2 = -36; end
		4968: begin l_1 = -27;
				 l_2 = +36; end
		10041: begin l_1 = -27;
				 l_2 = -36; end
		8178: begin l_1 = +27;
				 l_2 = +37; end
		4487: begin l_1 = +27;
				 l_2 = -37; end
		9350: begin l_1 = -27;
				 l_2 = +37; end
		5659: begin l_1 = -27;
				 l_2 = -37; end
		3105: begin l_1 = +27;
				 l_2 = +38; end
		9560: begin l_1 = +27;
				 l_2 = -38; end
		4277: begin l_1 = -27;
				 l_2 = +38; end
		10732: begin l_1 = -27;
				 l_2 = -38; end
		10321: begin l_1 = -28;
				 l_2 = +30; end
		3516: begin l_1 = -28;
				 l_2 = -29; end
		7977: begin l_1 = +28;
				 l_2 = +30; end
		5860: begin l_1 = -28;
				 l_2 = -30; end
		3289: begin l_1 = +28;
				 l_2 = +31; end
		8204: begin l_1 = +28;
				 l_2 = -31; end
		5633: begin l_1 = -28;
				 l_2 = +31; end
		10548: begin l_1 = -28;
				 l_2 = -31; end
		7750: begin l_1 = +28;
				 l_2 = +32; end
		3743: begin l_1 = +28;
				 l_2 = -32; end
		10094: begin l_1 = -28;
				 l_2 = +32; end
		6087: begin l_1 = -28;
				 l_2 = -32; end
		2835: begin l_1 = +28;
				 l_2 = +33; end
		8658: begin l_1 = +28;
				 l_2 = -33; end
		5179: begin l_1 = -28;
				 l_2 = +33; end
		11002: begin l_1 = -28;
				 l_2 = -33; end
		6842: begin l_1 = +28;
				 l_2 = +34; end
		4651: begin l_1 = +28;
				 l_2 = -34; end
		9186: begin l_1 = -28;
				 l_2 = +34; end
		6995: begin l_1 = -28;
				 l_2 = -34; end
		1019: begin l_1 = +28;
				 l_2 = +35; end
		10474: begin l_1 = +28;
				 l_2 = -35; end
		3363: begin l_1 = -28;
				 l_2 = +35; end
		12818: begin l_1 = -28;
				 l_2 = -35; end
		3210: begin l_1 = +28;
				 l_2 = +36; end
		8283: begin l_1 = +28;
				 l_2 = -36; end
		5554: begin l_1 = -28;
				 l_2 = +36; end
		10627: begin l_1 = -28;
				 l_2 = -36; end
		7592: begin l_1 = +28;
				 l_2 = +37; end
		3901: begin l_1 = +28;
				 l_2 = -37; end
		9936: begin l_1 = -28;
				 l_2 = +37; end
		6245: begin l_1 = -28;
				 l_2 = -37; end
		2519: begin l_1 = +28;
				 l_2 = +38; end
		8974: begin l_1 = +28;
				 l_2 = -38; end
		4863: begin l_1 = -28;
				 l_2 = +38; end
		11318: begin l_1 = -28;
				 l_2 = -38; end
		6805: begin l_1 = -29;
				 l_2 = +31; end
		7032: begin l_1 = -29;
				 l_2 = -30; end
		2117: begin l_1 = +29;
				 l_2 = +31; end
		11720: begin l_1 = -29;
				 l_2 = -31; end
		6578: begin l_1 = +29;
				 l_2 = +32; end
		2571: begin l_1 = +29;
				 l_2 = -32; end
		11266: begin l_1 = -29;
				 l_2 = +32; end
		7259: begin l_1 = -29;
				 l_2 = -32; end
		1663: begin l_1 = +29;
				 l_2 = +33; end
		7486: begin l_1 = +29;
				 l_2 = -33; end
		6351: begin l_1 = -29;
				 l_2 = +33; end
		12174: begin l_1 = -29;
				 l_2 = -33; end
		5670: begin l_1 = +29;
				 l_2 = +34; end
		3479: begin l_1 = +29;
				 l_2 = -34; end
		10358: begin l_1 = -29;
				 l_2 = +34; end
		8167: begin l_1 = -29;
				 l_2 = -34; end
		13684: begin l_1 = +29;
				 l_2 = +35; end
		9302: begin l_1 = +29;
				 l_2 = -35; end
		4535: begin l_1 = -29;
				 l_2 = +35; end
		153: begin l_1 = -29;
				 l_2 = -35; end
		2038: begin l_1 = +29;
				 l_2 = +36; end
		7111: begin l_1 = +29;
				 l_2 = -36; end
		6726: begin l_1 = -29;
				 l_2 = +36; end
		11799: begin l_1 = -29;
				 l_2 = -36; end
		6420: begin l_1 = +29;
				 l_2 = +37; end
		2729: begin l_1 = +29;
				 l_2 = -37; end
		11108: begin l_1 = -29;
				 l_2 = +37; end
		7417: begin l_1 = -29;
				 l_2 = -37; end
		1347: begin l_1 = +29;
				 l_2 = +38; end
		7802: begin l_1 = +29;
				 l_2 = -38; end
		6035: begin l_1 = -29;
				 l_2 = +38; end
		12490: begin l_1 = -29;
				 l_2 = -38; end
		13610: begin l_1 = -30;
				 l_2 = +32; end
		227: begin l_1 = -30;
				 l_2 = -31; end
		4234: begin l_1 = +30;
				 l_2 = +32; end
		9603: begin l_1 = -30;
				 l_2 = -32; end
		13156: begin l_1 = +30;
				 l_2 = +33; end
		5142: begin l_1 = +30;
				 l_2 = -33; end
		8695: begin l_1 = -30;
				 l_2 = +33; end
		681: begin l_1 = -30;
				 l_2 = -33; end
		3326: begin l_1 = +30;
				 l_2 = +34; end
		1135: begin l_1 = +30;
				 l_2 = -34; end
		12702: begin l_1 = -30;
				 l_2 = +34; end
		10511: begin l_1 = -30;
				 l_2 = -34; end
		11340: begin l_1 = +30;
				 l_2 = +35; end
		6958: begin l_1 = +30;
				 l_2 = -35; end
		6879: begin l_1 = -30;
				 l_2 = +35; end
		2497: begin l_1 = -30;
				 l_2 = -35; end
		13531: begin l_1 = +30;
				 l_2 = +36; end
		4767: begin l_1 = +30;
				 l_2 = -36; end
		9070: begin l_1 = -30;
				 l_2 = +36; end
		306: begin l_1 = -30;
				 l_2 = -36; end
		4076: begin l_1 = +30;
				 l_2 = +37; end
		385: begin l_1 = +30;
				 l_2 = -37; end
		13452: begin l_1 = -30;
				 l_2 = +37; end
		9761: begin l_1 = -30;
				 l_2 = -37; end
		12840: begin l_1 = +30;
				 l_2 = +38; end
		5458: begin l_1 = +30;
				 l_2 = -38; end
		8379: begin l_1 = -30;
				 l_2 = +38; end
		997: begin l_1 = -30;
				 l_2 = -38; end
		13383: begin l_1 = -31;
				 l_2 = +33; end
		454: begin l_1 = -31;
				 l_2 = -32; end
		8468: begin l_1 = +31;
				 l_2 = +33; end
		5369: begin l_1 = -31;
				 l_2 = -33; end
		12475: begin l_1 = +31;
				 l_2 = +34; end
		10284: begin l_1 = +31;
				 l_2 = -34; end
		3553: begin l_1 = -31;
				 l_2 = +34; end
		1362: begin l_1 = -31;
				 l_2 = -34; end
		6652: begin l_1 = +31;
				 l_2 = +35; end
		2270: begin l_1 = +31;
				 l_2 = -35; end
		11567: begin l_1 = -31;
				 l_2 = +35; end
		7185: begin l_1 = -31;
				 l_2 = -35; end
		8843: begin l_1 = +31;
				 l_2 = +36; end
		79: begin l_1 = +31;
				 l_2 = -36; end
		13758: begin l_1 = -31;
				 l_2 = +36; end
		4994: begin l_1 = -31;
				 l_2 = -36; end
		13225: begin l_1 = +31;
				 l_2 = +37; end
		9534: begin l_1 = +31;
				 l_2 = -37; end
		4303: begin l_1 = -31;
				 l_2 = +37; end
		612: begin l_1 = -31;
				 l_2 = -37; end
		8152: begin l_1 = +31;
				 l_2 = +38; end
		770: begin l_1 = +31;
				 l_2 = -38; end
		13067: begin l_1 = -31;
				 l_2 = +38; end
		5685: begin l_1 = -31;
				 l_2 = -38; end
		12929: begin l_1 = -32;
				 l_2 = +34; end
		908: begin l_1 = -32;
				 l_2 = -33; end
		3099: begin l_1 = +32;
				 l_2 = +34; end
		10738: begin l_1 = -32;
				 l_2 = -34; end
		11113: begin l_1 = +32;
				 l_2 = +35; end
		6731: begin l_1 = +32;
				 l_2 = -35; end
		7106: begin l_1 = -32;
				 l_2 = +35; end
		2724: begin l_1 = -32;
				 l_2 = -35; end
		13304: begin l_1 = +32;
				 l_2 = +36; end
		4540: begin l_1 = +32;
				 l_2 = -36; end
		9297: begin l_1 = -32;
				 l_2 = +36; end
		533: begin l_1 = -32;
				 l_2 = -36; end
		3849: begin l_1 = +32;
				 l_2 = +37; end
		158: begin l_1 = +32;
				 l_2 = -37; end
		13679: begin l_1 = -32;
				 l_2 = +37; end
		9988: begin l_1 = -32;
				 l_2 = -37; end
		12613: begin l_1 = +32;
				 l_2 = +38; end
		5231: begin l_1 = +32;
				 l_2 = -38; end
		8606: begin l_1 = -32;
				 l_2 = +38; end
		1224: begin l_1 = -32;
				 l_2 = -38; end
		12021: begin l_1 = -33;
				 l_2 = +35; end
		1816: begin l_1 = -33;
				 l_2 = -34; end
		6198: begin l_1 = +33;
				 l_2 = +35; end
		7639: begin l_1 = -33;
				 l_2 = -35; end
		8389: begin l_1 = +33;
				 l_2 = +36; end
		13462: begin l_1 = +33;
				 l_2 = -36; end
		375: begin l_1 = -33;
				 l_2 = +36; end
		5448: begin l_1 = -33;
				 l_2 = -36; end
		12771: begin l_1 = +33;
				 l_2 = +37; end
		9080: begin l_1 = +33;
				 l_2 = -37; end
		4757: begin l_1 = -33;
				 l_2 = +37; end
		1066: begin l_1 = -33;
				 l_2 = -37; end
		7698: begin l_1 = +33;
				 l_2 = +38; end
		316: begin l_1 = +33;
				 l_2 = -38; end
		13521: begin l_1 = -33;
				 l_2 = +38; end
		6139: begin l_1 = -33;
				 l_2 = -38; end
		10205: begin l_1 = -34;
				 l_2 = +36; end
		3632: begin l_1 = -34;
				 l_2 = -35; end
		12396: begin l_1 = +34;
				 l_2 = +36; end
		1441: begin l_1 = -34;
				 l_2 = -36; end
		2941: begin l_1 = +34;
				 l_2 = +37; end
		13087: begin l_1 = +34;
				 l_2 = -37; end
		750: begin l_1 = -34;
				 l_2 = +37; end
		10896: begin l_1 = -34;
				 l_2 = -37; end
		11705: begin l_1 = +34;
				 l_2 = +38; end
		4323: begin l_1 = +34;
				 l_2 = -38; end
		9514: begin l_1 = -34;
				 l_2 = +38; end
		2132: begin l_1 = -34;
				 l_2 = -38; end
		6573: begin l_1 = -35;
				 l_2 = +37; end
		7264: begin l_1 = -35;
				 l_2 = -36; end
		10955: begin l_1 = +35;
				 l_2 = +37; end
		2882: begin l_1 = -35;
				 l_2 = -37; end
		5882: begin l_1 = +35;
				 l_2 = +38; end
		12337: begin l_1 = +35;
				 l_2 = -38; end
		1500: begin l_1 = -35;
				 l_2 = +38; end
		7955: begin l_1 = -35;
				 l_2 = -38; end
		13146: begin l_1 = -36;
				 l_2 = +38; end
		691: begin l_1 = -36;
				 l_2 = -37; end
		8073: begin l_1 = +36;
				 l_2 = +38; end
		5764: begin l_1 = -36;
				 l_2 = -38; end
		12455: begin l_1 = +37;
				 l_2 = +38; end
		1382: begin l_1 = -37;
				 l_2 = -38; end
		default: begin l_1 = 0;
					   l_2 = 0; end
	endcase
end

endmodule

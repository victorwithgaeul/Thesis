// Product (AN) Code SEC r-LUT
// SEC_rLUT20bits.v
// Received remainder r, output single error location.
module SEC_rLUT20bits(r, l);
input 	[12:0]	r;
output	reg	signed	[6:0]	l;
always@(*) begin
	case(r)
		1: l = +1;
		6310: l = -1;
		2: l = +2;
		6309: l = -2;
		4: l = +3;
		6307: l = -3;
		8: l = +4;
		6303: l = -4;
		16: l = +5;
		6295: l = -5;
		32: l = +6;
		6279: l = -6;
		64: l = +7;
		6247: l = -7;
		128: l = +8;
		6183: l = -8;
		256: l = +9;
		6055: l = -9;
		512: l = +10;
		5799: l = -10;
		1024: l = +11;
		5287: l = -11;
		2048: l = +12;
		4263: l = -12;
		4096: l = +13;
		2215: l = -13;
		1881: l = +14;
		4430: l = -14;
		3762: l = +15;
		2549: l = -15;
		1213: l = +16;
		5098: l = -16;
		2426: l = +17;
		3885: l = -17;
		4852: l = +18;
		1459: l = -18;
		3393: l = +19;
		2918: l = -19;
		475: l = +20;
		5836: l = -20;
		950: l = +21;
		5361: l = -21;
		1900: l = +22;
		4411: l = -22;
		3800: l = +23;
		2511: l = -23;
		1289: l = +24;
		5022: l = -24;
		2578: l = +25;
		3733: l = -25;
		5156: l = +26;
		1155: l = -26;
		4001: l = +27;
		2310: l = -27;
		1691: l = +28;
		4620: l = -28;
		3382: l = +29;
		2929: l = -29;
		453: l = +30;
		5858: l = -30;
		906: l = +31;
		5405: l = -31;
		1812: l = +32;
		4499: l = -32;
		3624: l = +33;
		2687: l = -33;
		default: l = 0;
	endcase
end

endmodule

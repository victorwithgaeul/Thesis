// Product (AN) Code SEC r-LUT
// SEC_rLUT16bits.v
// Received remainder r, output single error location.
module SEC_rLUT16bits(r, l);
input 	[12:0]	r;
output	reg	signed	[5:0]	l;
always@(*) begin
	case(r)
		1: l = +1;
		4546: l = -1;
		2: l = +2;
		4545: l = -2;
		4: l = +3;
		4543: l = -3;
		8: l = +4;
		4539: l = -4;
		16: l = +5;
		4531: l = -5;
		32: l = +6;
		4515: l = -6;
		64: l = +7;
		4483: l = -7;
		128: l = +8;
		4419: l = -8;
		256: l = +9;
		4291: l = -9;
		512: l = +10;
		4035: l = -10;
		1024: l = +11;
		3523: l = -11;
		2048: l = +12;
		2499: l = -12;
		4096: l = +13;
		451: l = -13;
		3645: l = +14;
		902: l = -14;
		2743: l = +15;
		1804: l = -15;
		939: l = +16;
		3608: l = -16;
		1878: l = +17;
		2669: l = -17;
		3756: l = +18;
		791: l = -18;
		2965: l = +19;
		1582: l = -19;
		1383: l = +20;
		3164: l = -20;
		2766: l = +21;
		1781: l = -21;
		985: l = +22;
		3562: l = -22;
		1970: l = +23;
		2577: l = -23;
		3940: l = +24;
		607: l = -24;
		3333: l = +25;
		1214: l = -25;
		2119: l = +26;
		2428: l = -26;
		4238: l = +27;
		309: l = -27;
		3929: l = +28;
		618: l = -28;
		3311: l = +29;
		1236: l = -29;
		default: l = 0;
	endcase
end

endmodule

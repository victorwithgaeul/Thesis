// Product (AN) Code DEC r-LUT
// DEC_rLUT52bits.v
// Used to do DEC, but corrected errors by locations, not AWE
// Received remainder r, output two error locations.
module DEC_rLUT52bits(r, l_1, l_2);
input 	[15:0]	r;
output	reg	signed	[7:0]	l_1;
output	reg	signed	[7:0]	l_2;
always@(*) begin
	case(r)
		1: begin l_1 = -1;
				 l_2 = +2; end
		50860: begin l_1 = +1;
				 l_2 = -2; end
		2: begin l_1 = +1;
				 l_2 = +1; end
		50859: begin l_1 = -1;
				 l_2 = -1; end
		4: begin l_1 = +2;
				 l_2 = +2; end
		50857: begin l_1 = -2;
				 l_2 = -2; end
		8: begin l_1 = +3;
				 l_2 = +3; end
		50853: begin l_1 = -3;
				 l_2 = -3; end
		16: begin l_1 = +4;
				 l_2 = +4; end
		50845: begin l_1 = -4;
				 l_2 = -4; end
		32: begin l_1 = +5;
				 l_2 = +5; end
		50829: begin l_1 = -5;
				 l_2 = -5; end
		64: begin l_1 = +6;
				 l_2 = +6; end
		50797: begin l_1 = -6;
				 l_2 = -6; end
		128: begin l_1 = +7;
				 l_2 = +7; end
		50733: begin l_1 = -7;
				 l_2 = -7; end
		256: begin l_1 = +8;
				 l_2 = +8; end
		50605: begin l_1 = -8;
				 l_2 = -8; end
		512: begin l_1 = +9;
				 l_2 = +9; end
		50349: begin l_1 = -9;
				 l_2 = -9; end
		1024: begin l_1 = +10;
				 l_2 = +10; end
		49837: begin l_1 = -10;
				 l_2 = -10; end
		2048: begin l_1 = +11;
				 l_2 = +11; end
		48813: begin l_1 = -11;
				 l_2 = -11; end
		4096: begin l_1 = +12;
				 l_2 = +12; end
		46765: begin l_1 = -12;
				 l_2 = -12; end
		8192: begin l_1 = +13;
				 l_2 = +13; end
		42669: begin l_1 = -13;
				 l_2 = -13; end
		16384: begin l_1 = +14;
				 l_2 = +14; end
		34477: begin l_1 = -14;
				 l_2 = -14; end
		32768: begin l_1 = +15;
				 l_2 = +15; end
		18093: begin l_1 = -15;
				 l_2 = -15; end
		14675: begin l_1 = +16;
				 l_2 = +16; end
		36186: begin l_1 = -16;
				 l_2 = -16; end
		29350: begin l_1 = +17;
				 l_2 = +17; end
		21511: begin l_1 = -17;
				 l_2 = -17; end
		7839: begin l_1 = +18;
				 l_2 = +18; end
		43022: begin l_1 = -18;
				 l_2 = -18; end
		15678: begin l_1 = +19;
				 l_2 = +19; end
		35183: begin l_1 = -19;
				 l_2 = -19; end
		31356: begin l_1 = +20;
				 l_2 = +20; end
		19505: begin l_1 = -20;
				 l_2 = -20; end
		11851: begin l_1 = +21;
				 l_2 = +21; end
		39010: begin l_1 = -21;
				 l_2 = -21; end
		23702: begin l_1 = +22;
				 l_2 = +22; end
		27159: begin l_1 = -22;
				 l_2 = -22; end
		47404: begin l_1 = +23;
				 l_2 = +23; end
		3457: begin l_1 = -23;
				 l_2 = -23; end
		43947: begin l_1 = +24;
				 l_2 = +24; end
		6914: begin l_1 = -24;
				 l_2 = -24; end
		37033: begin l_1 = +25;
				 l_2 = +25; end
		13828: begin l_1 = -25;
				 l_2 = -25; end
		23205: begin l_1 = +26;
				 l_2 = +26; end
		27656: begin l_1 = -26;
				 l_2 = -26; end
		46410: begin l_1 = +27;
				 l_2 = +27; end
		4451: begin l_1 = -27;
				 l_2 = -27; end
		41959: begin l_1 = +28;
				 l_2 = +28; end
		8902: begin l_1 = -28;
				 l_2 = -28; end
		33057: begin l_1 = +29;
				 l_2 = +29; end
		17804: begin l_1 = -29;
				 l_2 = -29; end
		15253: begin l_1 = +30;
				 l_2 = +30; end
		35608: begin l_1 = -30;
				 l_2 = -30; end
		30506: begin l_1 = +31;
				 l_2 = +31; end
		20355: begin l_1 = -31;
				 l_2 = -31; end
		10151: begin l_1 = +32;
				 l_2 = +32; end
		40710: begin l_1 = -32;
				 l_2 = -32; end
		20302: begin l_1 = +33;
				 l_2 = +33; end
		30559: begin l_1 = -33;
				 l_2 = -33; end
		40604: begin l_1 = +34;
				 l_2 = +34; end
		10257: begin l_1 = -34;
				 l_2 = -34; end
		30347: begin l_1 = +35;
				 l_2 = +35; end
		20514: begin l_1 = -35;
				 l_2 = -35; end
		9833: begin l_1 = +36;
				 l_2 = +36; end
		41028: begin l_1 = -36;
				 l_2 = -36; end
		19666: begin l_1 = +37;
				 l_2 = +37; end
		31195: begin l_1 = -37;
				 l_2 = -37; end
		39332: begin l_1 = +38;
				 l_2 = +38; end
		11529: begin l_1 = -38;
				 l_2 = -38; end
		27803: begin l_1 = +39;
				 l_2 = +39; end
		23058: begin l_1 = -39;
				 l_2 = -39; end
		4745: begin l_1 = +40;
				 l_2 = +40; end
		46116: begin l_1 = -40;
				 l_2 = -40; end
		9490: begin l_1 = +41;
				 l_2 = +41; end
		41371: begin l_1 = -41;
				 l_2 = -41; end
		18980: begin l_1 = +42;
				 l_2 = +42; end
		31881: begin l_1 = -42;
				 l_2 = -42; end
		37960: begin l_1 = +43;
				 l_2 = +43; end
		12901: begin l_1 = -43;
				 l_2 = -43; end
		25059: begin l_1 = +44;
				 l_2 = +44; end
		25802: begin l_1 = -44;
				 l_2 = -44; end
		50118: begin l_1 = +45;
				 l_2 = +45; end
		743: begin l_1 = -45;
				 l_2 = -45; end
		49375: begin l_1 = +46;
				 l_2 = +46; end
		1486: begin l_1 = -46;
				 l_2 = -46; end
		47889: begin l_1 = +47;
				 l_2 = +47; end
		2972: begin l_1 = -47;
				 l_2 = -47; end
		44917: begin l_1 = +48;
				 l_2 = +48; end
		5944: begin l_1 = -48;
				 l_2 = -48; end
		38973: begin l_1 = +49;
				 l_2 = +49; end
		11888: begin l_1 = -49;
				 l_2 = -49; end
		27085: begin l_1 = +50;
				 l_2 = +50; end
		23776: begin l_1 = -50;
				 l_2 = -50; end
		3309: begin l_1 = +51;
				 l_2 = +51; end
		47552: begin l_1 = -51;
				 l_2 = -51; end
		6618: begin l_1 = +52;
				 l_2 = +52; end
		44243: begin l_1 = -52;
				 l_2 = -52; end
		13236: begin l_1 = +53;
				 l_2 = +53; end
		37625: begin l_1 = -53;
				 l_2 = -53; end
		26472: begin l_1 = +54;
				 l_2 = +54; end
		24389: begin l_1 = -54;
				 l_2 = -54; end
		2083: begin l_1 = +55;
				 l_2 = +55; end
		48778: begin l_1 = -55;
				 l_2 = -55; end
		4166: begin l_1 = +56;
				 l_2 = +56; end
		46695: begin l_1 = -56;
				 l_2 = -56; end
		8332: begin l_1 = +57;
				 l_2 = +57; end
		42529: begin l_1 = -57;
				 l_2 = -57; end
		16664: begin l_1 = +58;
				 l_2 = +58; end
		34197: begin l_1 = -58;
				 l_2 = -58; end
		33328: begin l_1 = +59;
				 l_2 = +59; end
		17533: begin l_1 = -59;
				 l_2 = -59; end
		15795: begin l_1 = +60;
				 l_2 = +60; end
		35066: begin l_1 = -60;
				 l_2 = -60; end
		31590: begin l_1 = +61;
				 l_2 = +61; end
		19271: begin l_1 = -61;
				 l_2 = -61; end
		12319: begin l_1 = +62;
				 l_2 = +62; end
		38542: begin l_1 = -62;
				 l_2 = -62; end
		24638: begin l_1 = +63;
				 l_2 = +63; end
		26223: begin l_1 = -63;
				 l_2 = -63; end
		49276: begin l_1 = +64;
				 l_2 = +64; end
		1585: begin l_1 = -64;
				 l_2 = -64; end
		47691: begin l_1 = +65;
				 l_2 = +65; end
		3170: begin l_1 = -65;
				 l_2 = -65; end
		44521: begin l_1 = +66;
				 l_2 = +66; end
		6340: begin l_1 = -66;
				 l_2 = -66; end
		38181: begin l_1 = +67;
				 l_2 = +67; end
		12680: begin l_1 = -67;
				 l_2 = -67; end
		3: begin l_1 = -1;
				 l_2 = +3; end
		50858: begin l_1 = -1;
				 l_2 = -2; end
		5: begin l_1 = +1;
				 l_2 = +3; end
		50856: begin l_1 = -1;
				 l_2 = -3; end
		9: begin l_1 = +1;
				 l_2 = +4; end
		50854: begin l_1 = +1;
				 l_2 = -4; end
		7: begin l_1 = -1;
				 l_2 = +4; end
		50852: begin l_1 = -1;
				 l_2 = -4; end
		17: begin l_1 = +1;
				 l_2 = +5; end
		50846: begin l_1 = +1;
				 l_2 = -5; end
		15: begin l_1 = -1;
				 l_2 = +5; end
		50844: begin l_1 = -1;
				 l_2 = -5; end
		33: begin l_1 = +1;
				 l_2 = +6; end
		50830: begin l_1 = +1;
				 l_2 = -6; end
		31: begin l_1 = -1;
				 l_2 = +6; end
		50828: begin l_1 = -1;
				 l_2 = -6; end
		65: begin l_1 = +1;
				 l_2 = +7; end
		50798: begin l_1 = +1;
				 l_2 = -7; end
		63: begin l_1 = -1;
				 l_2 = +7; end
		50796: begin l_1 = -1;
				 l_2 = -7; end
		129: begin l_1 = +1;
				 l_2 = +8; end
		50734: begin l_1 = +1;
				 l_2 = -8; end
		127: begin l_1 = -1;
				 l_2 = +8; end
		50732: begin l_1 = -1;
				 l_2 = -8; end
		257: begin l_1 = +1;
				 l_2 = +9; end
		50606: begin l_1 = +1;
				 l_2 = -9; end
		255: begin l_1 = -1;
				 l_2 = +9; end
		50604: begin l_1 = -1;
				 l_2 = -9; end
		513: begin l_1 = +1;
				 l_2 = +10; end
		50350: begin l_1 = +1;
				 l_2 = -10; end
		511: begin l_1 = -1;
				 l_2 = +10; end
		50348: begin l_1 = -1;
				 l_2 = -10; end
		1025: begin l_1 = +1;
				 l_2 = +11; end
		49838: begin l_1 = +1;
				 l_2 = -11; end
		1023: begin l_1 = -1;
				 l_2 = +11; end
		49836: begin l_1 = -1;
				 l_2 = -11; end
		2049: begin l_1 = +1;
				 l_2 = +12; end
		48814: begin l_1 = +1;
				 l_2 = -12; end
		2047: begin l_1 = -1;
				 l_2 = +12; end
		48812: begin l_1 = -1;
				 l_2 = -12; end
		4097: begin l_1 = +1;
				 l_2 = +13; end
		46766: begin l_1 = +1;
				 l_2 = -13; end
		4095: begin l_1 = -1;
				 l_2 = +13; end
		46764: begin l_1 = -1;
				 l_2 = -13; end
		8193: begin l_1 = +1;
				 l_2 = +14; end
		42670: begin l_1 = +1;
				 l_2 = -14; end
		8191: begin l_1 = -1;
				 l_2 = +14; end
		42668: begin l_1 = -1;
				 l_2 = -14; end
		16385: begin l_1 = +1;
				 l_2 = +15; end
		34478: begin l_1 = +1;
				 l_2 = -15; end
		16383: begin l_1 = -1;
				 l_2 = +15; end
		34476: begin l_1 = -1;
				 l_2 = -15; end
		32769: begin l_1 = +1;
				 l_2 = +16; end
		18094: begin l_1 = +1;
				 l_2 = -16; end
		32767: begin l_1 = -1;
				 l_2 = +16; end
		18092: begin l_1 = -1;
				 l_2 = -16; end
		14676: begin l_1 = +1;
				 l_2 = +17; end
		36187: begin l_1 = +1;
				 l_2 = -17; end
		14674: begin l_1 = -1;
				 l_2 = +17; end
		36185: begin l_1 = -1;
				 l_2 = -17; end
		29351: begin l_1 = +1;
				 l_2 = +18; end
		21512: begin l_1 = +1;
				 l_2 = -18; end
		29349: begin l_1 = -1;
				 l_2 = +18; end
		21510: begin l_1 = -1;
				 l_2 = -18; end
		7840: begin l_1 = +1;
				 l_2 = +19; end
		43023: begin l_1 = +1;
				 l_2 = -19; end
		7838: begin l_1 = -1;
				 l_2 = +19; end
		43021: begin l_1 = -1;
				 l_2 = -19; end
		15679: begin l_1 = +1;
				 l_2 = +20; end
		35184: begin l_1 = +1;
				 l_2 = -20; end
		15677: begin l_1 = -1;
				 l_2 = +20; end
		35182: begin l_1 = -1;
				 l_2 = -20; end
		31357: begin l_1 = +1;
				 l_2 = +21; end
		19506: begin l_1 = +1;
				 l_2 = -21; end
		31355: begin l_1 = -1;
				 l_2 = +21; end
		19504: begin l_1 = -1;
				 l_2 = -21; end
		11852: begin l_1 = +1;
				 l_2 = +22; end
		39011: begin l_1 = +1;
				 l_2 = -22; end
		11850: begin l_1 = -1;
				 l_2 = +22; end
		39009: begin l_1 = -1;
				 l_2 = -22; end
		23703: begin l_1 = +1;
				 l_2 = +23; end
		27160: begin l_1 = +1;
				 l_2 = -23; end
		23701: begin l_1 = -1;
				 l_2 = +23; end
		27158: begin l_1 = -1;
				 l_2 = -23; end
		47405: begin l_1 = +1;
				 l_2 = +24; end
		3458: begin l_1 = +1;
				 l_2 = -24; end
		47403: begin l_1 = -1;
				 l_2 = +24; end
		3456: begin l_1 = -1;
				 l_2 = -24; end
		43948: begin l_1 = +1;
				 l_2 = +25; end
		6915: begin l_1 = +1;
				 l_2 = -25; end
		43946: begin l_1 = -1;
				 l_2 = +25; end
		6913: begin l_1 = -1;
				 l_2 = -25; end
		37034: begin l_1 = +1;
				 l_2 = +26; end
		13829: begin l_1 = +1;
				 l_2 = -26; end
		37032: begin l_1 = -1;
				 l_2 = +26; end
		13827: begin l_1 = -1;
				 l_2 = -26; end
		23206: begin l_1 = +1;
				 l_2 = +27; end
		27657: begin l_1 = +1;
				 l_2 = -27; end
		23204: begin l_1 = -1;
				 l_2 = +27; end
		27655: begin l_1 = -1;
				 l_2 = -27; end
		46411: begin l_1 = +1;
				 l_2 = +28; end
		4452: begin l_1 = +1;
				 l_2 = -28; end
		46409: begin l_1 = -1;
				 l_2 = +28; end
		4450: begin l_1 = -1;
				 l_2 = -28; end
		41960: begin l_1 = +1;
				 l_2 = +29; end
		8903: begin l_1 = +1;
				 l_2 = -29; end
		41958: begin l_1 = -1;
				 l_2 = +29; end
		8901: begin l_1 = -1;
				 l_2 = -29; end
		33058: begin l_1 = +1;
				 l_2 = +30; end
		17805: begin l_1 = +1;
				 l_2 = -30; end
		33056: begin l_1 = -1;
				 l_2 = +30; end
		17803: begin l_1 = -1;
				 l_2 = -30; end
		15254: begin l_1 = +1;
				 l_2 = +31; end
		35609: begin l_1 = +1;
				 l_2 = -31; end
		15252: begin l_1 = -1;
				 l_2 = +31; end
		35607: begin l_1 = -1;
				 l_2 = -31; end
		30507: begin l_1 = +1;
				 l_2 = +32; end
		20356: begin l_1 = +1;
				 l_2 = -32; end
		30505: begin l_1 = -1;
				 l_2 = +32; end
		20354: begin l_1 = -1;
				 l_2 = -32; end
		10152: begin l_1 = +1;
				 l_2 = +33; end
		40711: begin l_1 = +1;
				 l_2 = -33; end
		10150: begin l_1 = -1;
				 l_2 = +33; end
		40709: begin l_1 = -1;
				 l_2 = -33; end
		20303: begin l_1 = +1;
				 l_2 = +34; end
		30560: begin l_1 = +1;
				 l_2 = -34; end
		20301: begin l_1 = -1;
				 l_2 = +34; end
		30558: begin l_1 = -1;
				 l_2 = -34; end
		40605: begin l_1 = +1;
				 l_2 = +35; end
		10258: begin l_1 = +1;
				 l_2 = -35; end
		40603: begin l_1 = -1;
				 l_2 = +35; end
		10256: begin l_1 = -1;
				 l_2 = -35; end
		30348: begin l_1 = +1;
				 l_2 = +36; end
		20515: begin l_1 = +1;
				 l_2 = -36; end
		30346: begin l_1 = -1;
				 l_2 = +36; end
		20513: begin l_1 = -1;
				 l_2 = -36; end
		9834: begin l_1 = +1;
				 l_2 = +37; end
		41029: begin l_1 = +1;
				 l_2 = -37; end
		9832: begin l_1 = -1;
				 l_2 = +37; end
		41027: begin l_1 = -1;
				 l_2 = -37; end
		19667: begin l_1 = +1;
				 l_2 = +38; end
		31196: begin l_1 = +1;
				 l_2 = -38; end
		19665: begin l_1 = -1;
				 l_2 = +38; end
		31194: begin l_1 = -1;
				 l_2 = -38; end
		39333: begin l_1 = +1;
				 l_2 = +39; end
		11530: begin l_1 = +1;
				 l_2 = -39; end
		39331: begin l_1 = -1;
				 l_2 = +39; end
		11528: begin l_1 = -1;
				 l_2 = -39; end
		27804: begin l_1 = +1;
				 l_2 = +40; end
		23059: begin l_1 = +1;
				 l_2 = -40; end
		27802: begin l_1 = -1;
				 l_2 = +40; end
		23057: begin l_1 = -1;
				 l_2 = -40; end
		4746: begin l_1 = +1;
				 l_2 = +41; end
		46117: begin l_1 = +1;
				 l_2 = -41; end
		4744: begin l_1 = -1;
				 l_2 = +41; end
		46115: begin l_1 = -1;
				 l_2 = -41; end
		9491: begin l_1 = +1;
				 l_2 = +42; end
		41372: begin l_1 = +1;
				 l_2 = -42; end
		9489: begin l_1 = -1;
				 l_2 = +42; end
		41370: begin l_1 = -1;
				 l_2 = -42; end
		18981: begin l_1 = +1;
				 l_2 = +43; end
		31882: begin l_1 = +1;
				 l_2 = -43; end
		18979: begin l_1 = -1;
				 l_2 = +43; end
		31880: begin l_1 = -1;
				 l_2 = -43; end
		37961: begin l_1 = +1;
				 l_2 = +44; end
		12902: begin l_1 = +1;
				 l_2 = -44; end
		37959: begin l_1 = -1;
				 l_2 = +44; end
		12900: begin l_1 = -1;
				 l_2 = -44; end
		25060: begin l_1 = +1;
				 l_2 = +45; end
		25803: begin l_1 = +1;
				 l_2 = -45; end
		25058: begin l_1 = -1;
				 l_2 = +45; end
		25801: begin l_1 = -1;
				 l_2 = -45; end
		50119: begin l_1 = +1;
				 l_2 = +46; end
		744: begin l_1 = +1;
				 l_2 = -46; end
		50117: begin l_1 = -1;
				 l_2 = +46; end
		742: begin l_1 = -1;
				 l_2 = -46; end
		49376: begin l_1 = +1;
				 l_2 = +47; end
		1487: begin l_1 = +1;
				 l_2 = -47; end
		49374: begin l_1 = -1;
				 l_2 = +47; end
		1485: begin l_1 = -1;
				 l_2 = -47; end
		47890: begin l_1 = +1;
				 l_2 = +48; end
		2973: begin l_1 = +1;
				 l_2 = -48; end
		47888: begin l_1 = -1;
				 l_2 = +48; end
		2971: begin l_1 = -1;
				 l_2 = -48; end
		44918: begin l_1 = +1;
				 l_2 = +49; end
		5945: begin l_1 = +1;
				 l_2 = -49; end
		44916: begin l_1 = -1;
				 l_2 = +49; end
		5943: begin l_1 = -1;
				 l_2 = -49; end
		38974: begin l_1 = +1;
				 l_2 = +50; end
		11889: begin l_1 = +1;
				 l_2 = -50; end
		38972: begin l_1 = -1;
				 l_2 = +50; end
		11887: begin l_1 = -1;
				 l_2 = -50; end
		27086: begin l_1 = +1;
				 l_2 = +51; end
		23777: begin l_1 = +1;
				 l_2 = -51; end
		27084: begin l_1 = -1;
				 l_2 = +51; end
		23775: begin l_1 = -1;
				 l_2 = -51; end
		3310: begin l_1 = +1;
				 l_2 = +52; end
		47553: begin l_1 = +1;
				 l_2 = -52; end
		3308: begin l_1 = -1;
				 l_2 = +52; end
		47551: begin l_1 = -1;
				 l_2 = -52; end
		6619: begin l_1 = +1;
				 l_2 = +53; end
		44244: begin l_1 = +1;
				 l_2 = -53; end
		6617: begin l_1 = -1;
				 l_2 = +53; end
		44242: begin l_1 = -1;
				 l_2 = -53; end
		13237: begin l_1 = +1;
				 l_2 = +54; end
		37626: begin l_1 = +1;
				 l_2 = -54; end
		13235: begin l_1 = -1;
				 l_2 = +54; end
		37624: begin l_1 = -1;
				 l_2 = -54; end
		26473: begin l_1 = +1;
				 l_2 = +55; end
		24390: begin l_1 = +1;
				 l_2 = -55; end
		26471: begin l_1 = -1;
				 l_2 = +55; end
		24388: begin l_1 = -1;
				 l_2 = -55; end
		2084: begin l_1 = +1;
				 l_2 = +56; end
		48779: begin l_1 = +1;
				 l_2 = -56; end
		2082: begin l_1 = -1;
				 l_2 = +56; end
		48777: begin l_1 = -1;
				 l_2 = -56; end
		4167: begin l_1 = +1;
				 l_2 = +57; end
		46696: begin l_1 = +1;
				 l_2 = -57; end
		4165: begin l_1 = -1;
				 l_2 = +57; end
		46694: begin l_1 = -1;
				 l_2 = -57; end
		8333: begin l_1 = +1;
				 l_2 = +58; end
		42530: begin l_1 = +1;
				 l_2 = -58; end
		8331: begin l_1 = -1;
				 l_2 = +58; end
		42528: begin l_1 = -1;
				 l_2 = -58; end
		16665: begin l_1 = +1;
				 l_2 = +59; end
		34198: begin l_1 = +1;
				 l_2 = -59; end
		16663: begin l_1 = -1;
				 l_2 = +59; end
		34196: begin l_1 = -1;
				 l_2 = -59; end
		33329: begin l_1 = +1;
				 l_2 = +60; end
		17534: begin l_1 = +1;
				 l_2 = -60; end
		33327: begin l_1 = -1;
				 l_2 = +60; end
		17532: begin l_1 = -1;
				 l_2 = -60; end
		15796: begin l_1 = +1;
				 l_2 = +61; end
		35067: begin l_1 = +1;
				 l_2 = -61; end
		15794: begin l_1 = -1;
				 l_2 = +61; end
		35065: begin l_1 = -1;
				 l_2 = -61; end
		31591: begin l_1 = +1;
				 l_2 = +62; end
		19272: begin l_1 = +1;
				 l_2 = -62; end
		31589: begin l_1 = -1;
				 l_2 = +62; end
		19270: begin l_1 = -1;
				 l_2 = -62; end
		12320: begin l_1 = +1;
				 l_2 = +63; end
		38543: begin l_1 = +1;
				 l_2 = -63; end
		12318: begin l_1 = -1;
				 l_2 = +63; end
		38541: begin l_1 = -1;
				 l_2 = -63; end
		24639: begin l_1 = +1;
				 l_2 = +64; end
		26224: begin l_1 = +1;
				 l_2 = -64; end
		24637: begin l_1 = -1;
				 l_2 = +64; end
		26222: begin l_1 = -1;
				 l_2 = -64; end
		49277: begin l_1 = +1;
				 l_2 = +65; end
		1586: begin l_1 = +1;
				 l_2 = -65; end
		49275: begin l_1 = -1;
				 l_2 = +65; end
		1584: begin l_1 = -1;
				 l_2 = -65; end
		47692: begin l_1 = +1;
				 l_2 = +66; end
		3171: begin l_1 = +1;
				 l_2 = -66; end
		47690: begin l_1 = -1;
				 l_2 = +66; end
		3169: begin l_1 = -1;
				 l_2 = -66; end
		44522: begin l_1 = +1;
				 l_2 = +67; end
		6341: begin l_1 = +1;
				 l_2 = -67; end
		44520: begin l_1 = -1;
				 l_2 = +67; end
		6339: begin l_1 = -1;
				 l_2 = -67; end
		38182: begin l_1 = +1;
				 l_2 = +68; end
		12681: begin l_1 = +1;
				 l_2 = -68; end
		38180: begin l_1 = -1;
				 l_2 = +68; end
		12679: begin l_1 = -1;
				 l_2 = -68; end
		6: begin l_1 = -2;
				 l_2 = +4; end
		50855: begin l_1 = -2;
				 l_2 = -3; end
		10: begin l_1 = +2;
				 l_2 = +4; end
		50851: begin l_1 = -2;
				 l_2 = -4; end
		18: begin l_1 = +2;
				 l_2 = +5; end
		50847: begin l_1 = +2;
				 l_2 = -5; end
		14: begin l_1 = -2;
				 l_2 = +5; end
		50843: begin l_1 = -2;
				 l_2 = -5; end
		34: begin l_1 = +2;
				 l_2 = +6; end
		50831: begin l_1 = +2;
				 l_2 = -6; end
		30: begin l_1 = -2;
				 l_2 = +6; end
		50827: begin l_1 = -2;
				 l_2 = -6; end
		66: begin l_1 = +2;
				 l_2 = +7; end
		50799: begin l_1 = +2;
				 l_2 = -7; end
		62: begin l_1 = -2;
				 l_2 = +7; end
		50795: begin l_1 = -2;
				 l_2 = -7; end
		130: begin l_1 = +2;
				 l_2 = +8; end
		50735: begin l_1 = +2;
				 l_2 = -8; end
		126: begin l_1 = -2;
				 l_2 = +8; end
		50731: begin l_1 = -2;
				 l_2 = -8; end
		258: begin l_1 = +2;
				 l_2 = +9; end
		50607: begin l_1 = +2;
				 l_2 = -9; end
		254: begin l_1 = -2;
				 l_2 = +9; end
		50603: begin l_1 = -2;
				 l_2 = -9; end
		514: begin l_1 = +2;
				 l_2 = +10; end
		50351: begin l_1 = +2;
				 l_2 = -10; end
		510: begin l_1 = -2;
				 l_2 = +10; end
		50347: begin l_1 = -2;
				 l_2 = -10; end
		1026: begin l_1 = +2;
				 l_2 = +11; end
		49839: begin l_1 = +2;
				 l_2 = -11; end
		1022: begin l_1 = -2;
				 l_2 = +11; end
		49835: begin l_1 = -2;
				 l_2 = -11; end
		2050: begin l_1 = +2;
				 l_2 = +12; end
		48815: begin l_1 = +2;
				 l_2 = -12; end
		2046: begin l_1 = -2;
				 l_2 = +12; end
		48811: begin l_1 = -2;
				 l_2 = -12; end
		4098: begin l_1 = +2;
				 l_2 = +13; end
		46767: begin l_1 = +2;
				 l_2 = -13; end
		4094: begin l_1 = -2;
				 l_2 = +13; end
		46763: begin l_1 = -2;
				 l_2 = -13; end
		8194: begin l_1 = +2;
				 l_2 = +14; end
		42671: begin l_1 = +2;
				 l_2 = -14; end
		8190: begin l_1 = -2;
				 l_2 = +14; end
		42667: begin l_1 = -2;
				 l_2 = -14; end
		16386: begin l_1 = +2;
				 l_2 = +15; end
		34479: begin l_1 = +2;
				 l_2 = -15; end
		16382: begin l_1 = -2;
				 l_2 = +15; end
		34475: begin l_1 = -2;
				 l_2 = -15; end
		32770: begin l_1 = +2;
				 l_2 = +16; end
		18095: begin l_1 = +2;
				 l_2 = -16; end
		32766: begin l_1 = -2;
				 l_2 = +16; end
		18091: begin l_1 = -2;
				 l_2 = -16; end
		14677: begin l_1 = +2;
				 l_2 = +17; end
		36188: begin l_1 = +2;
				 l_2 = -17; end
		14673: begin l_1 = -2;
				 l_2 = +17; end
		36184: begin l_1 = -2;
				 l_2 = -17; end
		29352: begin l_1 = +2;
				 l_2 = +18; end
		21513: begin l_1 = +2;
				 l_2 = -18; end
		29348: begin l_1 = -2;
				 l_2 = +18; end
		21509: begin l_1 = -2;
				 l_2 = -18; end
		7841: begin l_1 = +2;
				 l_2 = +19; end
		43024: begin l_1 = +2;
				 l_2 = -19; end
		7837: begin l_1 = -2;
				 l_2 = +19; end
		43020: begin l_1 = -2;
				 l_2 = -19; end
		15680: begin l_1 = +2;
				 l_2 = +20; end
		35185: begin l_1 = +2;
				 l_2 = -20; end
		15676: begin l_1 = -2;
				 l_2 = +20; end
		35181: begin l_1 = -2;
				 l_2 = -20; end
		31358: begin l_1 = +2;
				 l_2 = +21; end
		19507: begin l_1 = +2;
				 l_2 = -21; end
		31354: begin l_1 = -2;
				 l_2 = +21; end
		19503: begin l_1 = -2;
				 l_2 = -21; end
		11853: begin l_1 = +2;
				 l_2 = +22; end
		39012: begin l_1 = +2;
				 l_2 = -22; end
		11849: begin l_1 = -2;
				 l_2 = +22; end
		39008: begin l_1 = -2;
				 l_2 = -22; end
		23704: begin l_1 = +2;
				 l_2 = +23; end
		27161: begin l_1 = +2;
				 l_2 = -23; end
		23700: begin l_1 = -2;
				 l_2 = +23; end
		27157: begin l_1 = -2;
				 l_2 = -23; end
		47406: begin l_1 = +2;
				 l_2 = +24; end
		3459: begin l_1 = +2;
				 l_2 = -24; end
		47402: begin l_1 = -2;
				 l_2 = +24; end
		3455: begin l_1 = -2;
				 l_2 = -24; end
		43949: begin l_1 = +2;
				 l_2 = +25; end
		6916: begin l_1 = +2;
				 l_2 = -25; end
		43945: begin l_1 = -2;
				 l_2 = +25; end
		6912: begin l_1 = -2;
				 l_2 = -25; end
		37035: begin l_1 = +2;
				 l_2 = +26; end
		13830: begin l_1 = +2;
				 l_2 = -26; end
		37031: begin l_1 = -2;
				 l_2 = +26; end
		13826: begin l_1 = -2;
				 l_2 = -26; end
		23207: begin l_1 = +2;
				 l_2 = +27; end
		27658: begin l_1 = +2;
				 l_2 = -27; end
		23203: begin l_1 = -2;
				 l_2 = +27; end
		27654: begin l_1 = -2;
				 l_2 = -27; end
		46412: begin l_1 = +2;
				 l_2 = +28; end
		4453: begin l_1 = +2;
				 l_2 = -28; end
		46408: begin l_1 = -2;
				 l_2 = +28; end
		4449: begin l_1 = -2;
				 l_2 = -28; end
		41961: begin l_1 = +2;
				 l_2 = +29; end
		8904: begin l_1 = +2;
				 l_2 = -29; end
		41957: begin l_1 = -2;
				 l_2 = +29; end
		8900: begin l_1 = -2;
				 l_2 = -29; end
		33059: begin l_1 = +2;
				 l_2 = +30; end
		17806: begin l_1 = +2;
				 l_2 = -30; end
		33055: begin l_1 = -2;
				 l_2 = +30; end
		17802: begin l_1 = -2;
				 l_2 = -30; end
		15255: begin l_1 = +2;
				 l_2 = +31; end
		35610: begin l_1 = +2;
				 l_2 = -31; end
		15251: begin l_1 = -2;
				 l_2 = +31; end
		35606: begin l_1 = -2;
				 l_2 = -31; end
		30508: begin l_1 = +2;
				 l_2 = +32; end
		20357: begin l_1 = +2;
				 l_2 = -32; end
		30504: begin l_1 = -2;
				 l_2 = +32; end
		20353: begin l_1 = -2;
				 l_2 = -32; end
		10153: begin l_1 = +2;
				 l_2 = +33; end
		40712: begin l_1 = +2;
				 l_2 = -33; end
		10149: begin l_1 = -2;
				 l_2 = +33; end
		40708: begin l_1 = -2;
				 l_2 = -33; end
		20304: begin l_1 = +2;
				 l_2 = +34; end
		30561: begin l_1 = +2;
				 l_2 = -34; end
		20300: begin l_1 = -2;
				 l_2 = +34; end
		30557: begin l_1 = -2;
				 l_2 = -34; end
		40606: begin l_1 = +2;
				 l_2 = +35; end
		10259: begin l_1 = +2;
				 l_2 = -35; end
		40602: begin l_1 = -2;
				 l_2 = +35; end
		10255: begin l_1 = -2;
				 l_2 = -35; end
		30349: begin l_1 = +2;
				 l_2 = +36; end
		20516: begin l_1 = +2;
				 l_2 = -36; end
		30345: begin l_1 = -2;
				 l_2 = +36; end
		20512: begin l_1 = -2;
				 l_2 = -36; end
		9835: begin l_1 = +2;
				 l_2 = +37; end
		41030: begin l_1 = +2;
				 l_2 = -37; end
		9831: begin l_1 = -2;
				 l_2 = +37; end
		41026: begin l_1 = -2;
				 l_2 = -37; end
		19668: begin l_1 = +2;
				 l_2 = +38; end
		31197: begin l_1 = +2;
				 l_2 = -38; end
		19664: begin l_1 = -2;
				 l_2 = +38; end
		31193: begin l_1 = -2;
				 l_2 = -38; end
		39334: begin l_1 = +2;
				 l_2 = +39; end
		11531: begin l_1 = +2;
				 l_2 = -39; end
		39330: begin l_1 = -2;
				 l_2 = +39; end
		11527: begin l_1 = -2;
				 l_2 = -39; end
		27805: begin l_1 = +2;
				 l_2 = +40; end
		23060: begin l_1 = +2;
				 l_2 = -40; end
		27801: begin l_1 = -2;
				 l_2 = +40; end
		23056: begin l_1 = -2;
				 l_2 = -40; end
		4747: begin l_1 = +2;
				 l_2 = +41; end
		46118: begin l_1 = +2;
				 l_2 = -41; end
		4743: begin l_1 = -2;
				 l_2 = +41; end
		46114: begin l_1 = -2;
				 l_2 = -41; end
		9492: begin l_1 = +2;
				 l_2 = +42; end
		41373: begin l_1 = +2;
				 l_2 = -42; end
		9488: begin l_1 = -2;
				 l_2 = +42; end
		41369: begin l_1 = -2;
				 l_2 = -42; end
		18982: begin l_1 = +2;
				 l_2 = +43; end
		31883: begin l_1 = +2;
				 l_2 = -43; end
		18978: begin l_1 = -2;
				 l_2 = +43; end
		31879: begin l_1 = -2;
				 l_2 = -43; end
		37962: begin l_1 = +2;
				 l_2 = +44; end
		12903: begin l_1 = +2;
				 l_2 = -44; end
		37958: begin l_1 = -2;
				 l_2 = +44; end
		12899: begin l_1 = -2;
				 l_2 = -44; end
		25061: begin l_1 = +2;
				 l_2 = +45; end
		25804: begin l_1 = +2;
				 l_2 = -45; end
		25057: begin l_1 = -2;
				 l_2 = +45; end
		25800: begin l_1 = -2;
				 l_2 = -45; end
		50120: begin l_1 = +2;
				 l_2 = +46; end
		745: begin l_1 = +2;
				 l_2 = -46; end
		50116: begin l_1 = -2;
				 l_2 = +46; end
		741: begin l_1 = -2;
				 l_2 = -46; end
		49377: begin l_1 = +2;
				 l_2 = +47; end
		1488: begin l_1 = +2;
				 l_2 = -47; end
		49373: begin l_1 = -2;
				 l_2 = +47; end
		1484: begin l_1 = -2;
				 l_2 = -47; end
		47891: begin l_1 = +2;
				 l_2 = +48; end
		2974: begin l_1 = +2;
				 l_2 = -48; end
		47887: begin l_1 = -2;
				 l_2 = +48; end
		2970: begin l_1 = -2;
				 l_2 = -48; end
		44919: begin l_1 = +2;
				 l_2 = +49; end
		5946: begin l_1 = +2;
				 l_2 = -49; end
		44915: begin l_1 = -2;
				 l_2 = +49; end
		5942: begin l_1 = -2;
				 l_2 = -49; end
		38975: begin l_1 = +2;
				 l_2 = +50; end
		11890: begin l_1 = +2;
				 l_2 = -50; end
		38971: begin l_1 = -2;
				 l_2 = +50; end
		11886: begin l_1 = -2;
				 l_2 = -50; end
		27087: begin l_1 = +2;
				 l_2 = +51; end
		23778: begin l_1 = +2;
				 l_2 = -51; end
		27083: begin l_1 = -2;
				 l_2 = +51; end
		23774: begin l_1 = -2;
				 l_2 = -51; end
		3311: begin l_1 = +2;
				 l_2 = +52; end
		47554: begin l_1 = +2;
				 l_2 = -52; end
		3307: begin l_1 = -2;
				 l_2 = +52; end
		47550: begin l_1 = -2;
				 l_2 = -52; end
		6620: begin l_1 = +2;
				 l_2 = +53; end
		44245: begin l_1 = +2;
				 l_2 = -53; end
		6616: begin l_1 = -2;
				 l_2 = +53; end
		44241: begin l_1 = -2;
				 l_2 = -53; end
		13238: begin l_1 = +2;
				 l_2 = +54; end
		37627: begin l_1 = +2;
				 l_2 = -54; end
		13234: begin l_1 = -2;
				 l_2 = +54; end
		37623: begin l_1 = -2;
				 l_2 = -54; end
		26474: begin l_1 = +2;
				 l_2 = +55; end
		24391: begin l_1 = +2;
				 l_2 = -55; end
		26470: begin l_1 = -2;
				 l_2 = +55; end
		24387: begin l_1 = -2;
				 l_2 = -55; end
		2085: begin l_1 = +2;
				 l_2 = +56; end
		48780: begin l_1 = +2;
				 l_2 = -56; end
		2081: begin l_1 = -2;
				 l_2 = +56; end
		48776: begin l_1 = -2;
				 l_2 = -56; end
		4168: begin l_1 = +2;
				 l_2 = +57; end
		46697: begin l_1 = +2;
				 l_2 = -57; end
		4164: begin l_1 = -2;
				 l_2 = +57; end
		46693: begin l_1 = -2;
				 l_2 = -57; end
		8334: begin l_1 = +2;
				 l_2 = +58; end
		42531: begin l_1 = +2;
				 l_2 = -58; end
		8330: begin l_1 = -2;
				 l_2 = +58; end
		42527: begin l_1 = -2;
				 l_2 = -58; end
		16666: begin l_1 = +2;
				 l_2 = +59; end
		34199: begin l_1 = +2;
				 l_2 = -59; end
		16662: begin l_1 = -2;
				 l_2 = +59; end
		34195: begin l_1 = -2;
				 l_2 = -59; end
		33330: begin l_1 = +2;
				 l_2 = +60; end
		17535: begin l_1 = +2;
				 l_2 = -60; end
		33326: begin l_1 = -2;
				 l_2 = +60; end
		17531: begin l_1 = -2;
				 l_2 = -60; end
		15797: begin l_1 = +2;
				 l_2 = +61; end
		35068: begin l_1 = +2;
				 l_2 = -61; end
		15793: begin l_1 = -2;
				 l_2 = +61; end
		35064: begin l_1 = -2;
				 l_2 = -61; end
		31592: begin l_1 = +2;
				 l_2 = +62; end
		19273: begin l_1 = +2;
				 l_2 = -62; end
		31588: begin l_1 = -2;
				 l_2 = +62; end
		19269: begin l_1 = -2;
				 l_2 = -62; end
		12321: begin l_1 = +2;
				 l_2 = +63; end
		38544: begin l_1 = +2;
				 l_2 = -63; end
		12317: begin l_1 = -2;
				 l_2 = +63; end
		38540: begin l_1 = -2;
				 l_2 = -63; end
		24640: begin l_1 = +2;
				 l_2 = +64; end
		26225: begin l_1 = +2;
				 l_2 = -64; end
		24636: begin l_1 = -2;
				 l_2 = +64; end
		26221: begin l_1 = -2;
				 l_2 = -64; end
		49278: begin l_1 = +2;
				 l_2 = +65; end
		1587: begin l_1 = +2;
				 l_2 = -65; end
		49274: begin l_1 = -2;
				 l_2 = +65; end
		1583: begin l_1 = -2;
				 l_2 = -65; end
		47693: begin l_1 = +2;
				 l_2 = +66; end
		3172: begin l_1 = +2;
				 l_2 = -66; end
		47689: begin l_1 = -2;
				 l_2 = +66; end
		3168: begin l_1 = -2;
				 l_2 = -66; end
		44523: begin l_1 = +2;
				 l_2 = +67; end
		6342: begin l_1 = +2;
				 l_2 = -67; end
		44519: begin l_1 = -2;
				 l_2 = +67; end
		6338: begin l_1 = -2;
				 l_2 = -67; end
		38183: begin l_1 = +2;
				 l_2 = +68; end
		12682: begin l_1 = +2;
				 l_2 = -68; end
		38179: begin l_1 = -2;
				 l_2 = +68; end
		12678: begin l_1 = -2;
				 l_2 = -68; end
		12: begin l_1 = -3;
				 l_2 = +5; end
		50849: begin l_1 = -3;
				 l_2 = -4; end
		20: begin l_1 = +3;
				 l_2 = +5; end
		50841: begin l_1 = -3;
				 l_2 = -5; end
		36: begin l_1 = +3;
				 l_2 = +6; end
		50833: begin l_1 = +3;
				 l_2 = -6; end
		28: begin l_1 = -3;
				 l_2 = +6; end
		50825: begin l_1 = -3;
				 l_2 = -6; end
		68: begin l_1 = +3;
				 l_2 = +7; end
		50801: begin l_1 = +3;
				 l_2 = -7; end
		60: begin l_1 = -3;
				 l_2 = +7; end
		50793: begin l_1 = -3;
				 l_2 = -7; end
		132: begin l_1 = +3;
				 l_2 = +8; end
		50737: begin l_1 = +3;
				 l_2 = -8; end
		124: begin l_1 = -3;
				 l_2 = +8; end
		50729: begin l_1 = -3;
				 l_2 = -8; end
		260: begin l_1 = +3;
				 l_2 = +9; end
		50609: begin l_1 = +3;
				 l_2 = -9; end
		252: begin l_1 = -3;
				 l_2 = +9; end
		50601: begin l_1 = -3;
				 l_2 = -9; end
		516: begin l_1 = +3;
				 l_2 = +10; end
		50353: begin l_1 = +3;
				 l_2 = -10; end
		508: begin l_1 = -3;
				 l_2 = +10; end
		50345: begin l_1 = -3;
				 l_2 = -10; end
		1028: begin l_1 = +3;
				 l_2 = +11; end
		49841: begin l_1 = +3;
				 l_2 = -11; end
		1020: begin l_1 = -3;
				 l_2 = +11; end
		49833: begin l_1 = -3;
				 l_2 = -11; end
		2052: begin l_1 = +3;
				 l_2 = +12; end
		48817: begin l_1 = +3;
				 l_2 = -12; end
		2044: begin l_1 = -3;
				 l_2 = +12; end
		48809: begin l_1 = -3;
				 l_2 = -12; end
		4100: begin l_1 = +3;
				 l_2 = +13; end
		46769: begin l_1 = +3;
				 l_2 = -13; end
		4092: begin l_1 = -3;
				 l_2 = +13; end
		46761: begin l_1 = -3;
				 l_2 = -13; end
		8196: begin l_1 = +3;
				 l_2 = +14; end
		42673: begin l_1 = +3;
				 l_2 = -14; end
		8188: begin l_1 = -3;
				 l_2 = +14; end
		42665: begin l_1 = -3;
				 l_2 = -14; end
		16388: begin l_1 = +3;
				 l_2 = +15; end
		34481: begin l_1 = +3;
				 l_2 = -15; end
		16380: begin l_1 = -3;
				 l_2 = +15; end
		34473: begin l_1 = -3;
				 l_2 = -15; end
		32772: begin l_1 = +3;
				 l_2 = +16; end
		18097: begin l_1 = +3;
				 l_2 = -16; end
		32764: begin l_1 = -3;
				 l_2 = +16; end
		18089: begin l_1 = -3;
				 l_2 = -16; end
		14679: begin l_1 = +3;
				 l_2 = +17; end
		36190: begin l_1 = +3;
				 l_2 = -17; end
		14671: begin l_1 = -3;
				 l_2 = +17; end
		36182: begin l_1 = -3;
				 l_2 = -17; end
		29354: begin l_1 = +3;
				 l_2 = +18; end
		21515: begin l_1 = +3;
				 l_2 = -18; end
		29346: begin l_1 = -3;
				 l_2 = +18; end
		21507: begin l_1 = -3;
				 l_2 = -18; end
		7843: begin l_1 = +3;
				 l_2 = +19; end
		43026: begin l_1 = +3;
				 l_2 = -19; end
		7835: begin l_1 = -3;
				 l_2 = +19; end
		43018: begin l_1 = -3;
				 l_2 = -19; end
		15682: begin l_1 = +3;
				 l_2 = +20; end
		35187: begin l_1 = +3;
				 l_2 = -20; end
		15674: begin l_1 = -3;
				 l_2 = +20; end
		35179: begin l_1 = -3;
				 l_2 = -20; end
		31360: begin l_1 = +3;
				 l_2 = +21; end
		19509: begin l_1 = +3;
				 l_2 = -21; end
		31352: begin l_1 = -3;
				 l_2 = +21; end
		19501: begin l_1 = -3;
				 l_2 = -21; end
		11855: begin l_1 = +3;
				 l_2 = +22; end
		39014: begin l_1 = +3;
				 l_2 = -22; end
		11847: begin l_1 = -3;
				 l_2 = +22; end
		39006: begin l_1 = -3;
				 l_2 = -22; end
		23706: begin l_1 = +3;
				 l_2 = +23; end
		27163: begin l_1 = +3;
				 l_2 = -23; end
		23698: begin l_1 = -3;
				 l_2 = +23; end
		27155: begin l_1 = -3;
				 l_2 = -23; end
		47408: begin l_1 = +3;
				 l_2 = +24; end
		3461: begin l_1 = +3;
				 l_2 = -24; end
		47400: begin l_1 = -3;
				 l_2 = +24; end
		3453: begin l_1 = -3;
				 l_2 = -24; end
		43951: begin l_1 = +3;
				 l_2 = +25; end
		6918: begin l_1 = +3;
				 l_2 = -25; end
		43943: begin l_1 = -3;
				 l_2 = +25; end
		6910: begin l_1 = -3;
				 l_2 = -25; end
		37037: begin l_1 = +3;
				 l_2 = +26; end
		13832: begin l_1 = +3;
				 l_2 = -26; end
		37029: begin l_1 = -3;
				 l_2 = +26; end
		13824: begin l_1 = -3;
				 l_2 = -26; end
		23209: begin l_1 = +3;
				 l_2 = +27; end
		27660: begin l_1 = +3;
				 l_2 = -27; end
		23201: begin l_1 = -3;
				 l_2 = +27; end
		27652: begin l_1 = -3;
				 l_2 = -27; end
		46414: begin l_1 = +3;
				 l_2 = +28; end
		4455: begin l_1 = +3;
				 l_2 = -28; end
		46406: begin l_1 = -3;
				 l_2 = +28; end
		4447: begin l_1 = -3;
				 l_2 = -28; end
		41963: begin l_1 = +3;
				 l_2 = +29; end
		8906: begin l_1 = +3;
				 l_2 = -29; end
		41955: begin l_1 = -3;
				 l_2 = +29; end
		8898: begin l_1 = -3;
				 l_2 = -29; end
		33061: begin l_1 = +3;
				 l_2 = +30; end
		17808: begin l_1 = +3;
				 l_2 = -30; end
		33053: begin l_1 = -3;
				 l_2 = +30; end
		17800: begin l_1 = -3;
				 l_2 = -30; end
		15257: begin l_1 = +3;
				 l_2 = +31; end
		35612: begin l_1 = +3;
				 l_2 = -31; end
		15249: begin l_1 = -3;
				 l_2 = +31; end
		35604: begin l_1 = -3;
				 l_2 = -31; end
		30510: begin l_1 = +3;
				 l_2 = +32; end
		20359: begin l_1 = +3;
				 l_2 = -32; end
		30502: begin l_1 = -3;
				 l_2 = +32; end
		20351: begin l_1 = -3;
				 l_2 = -32; end
		10155: begin l_1 = +3;
				 l_2 = +33; end
		40714: begin l_1 = +3;
				 l_2 = -33; end
		10147: begin l_1 = -3;
				 l_2 = +33; end
		40706: begin l_1 = -3;
				 l_2 = -33; end
		20306: begin l_1 = +3;
				 l_2 = +34; end
		30563: begin l_1 = +3;
				 l_2 = -34; end
		20298: begin l_1 = -3;
				 l_2 = +34; end
		30555: begin l_1 = -3;
				 l_2 = -34; end
		40608: begin l_1 = +3;
				 l_2 = +35; end
		10261: begin l_1 = +3;
				 l_2 = -35; end
		40600: begin l_1 = -3;
				 l_2 = +35; end
		10253: begin l_1 = -3;
				 l_2 = -35; end
		30351: begin l_1 = +3;
				 l_2 = +36; end
		20518: begin l_1 = +3;
				 l_2 = -36; end
		30343: begin l_1 = -3;
				 l_2 = +36; end
		20510: begin l_1 = -3;
				 l_2 = -36; end
		9837: begin l_1 = +3;
				 l_2 = +37; end
		41032: begin l_1 = +3;
				 l_2 = -37; end
		9829: begin l_1 = -3;
				 l_2 = +37; end
		41024: begin l_1 = -3;
				 l_2 = -37; end
		19670: begin l_1 = +3;
				 l_2 = +38; end
		31199: begin l_1 = +3;
				 l_2 = -38; end
		19662: begin l_1 = -3;
				 l_2 = +38; end
		31191: begin l_1 = -3;
				 l_2 = -38; end
		39336: begin l_1 = +3;
				 l_2 = +39; end
		11533: begin l_1 = +3;
				 l_2 = -39; end
		39328: begin l_1 = -3;
				 l_2 = +39; end
		11525: begin l_1 = -3;
				 l_2 = -39; end
		27807: begin l_1 = +3;
				 l_2 = +40; end
		23062: begin l_1 = +3;
				 l_2 = -40; end
		27799: begin l_1 = -3;
				 l_2 = +40; end
		23054: begin l_1 = -3;
				 l_2 = -40; end
		4749: begin l_1 = +3;
				 l_2 = +41; end
		46120: begin l_1 = +3;
				 l_2 = -41; end
		4741: begin l_1 = -3;
				 l_2 = +41; end
		46112: begin l_1 = -3;
				 l_2 = -41; end
		9494: begin l_1 = +3;
				 l_2 = +42; end
		41375: begin l_1 = +3;
				 l_2 = -42; end
		9486: begin l_1 = -3;
				 l_2 = +42; end
		41367: begin l_1 = -3;
				 l_2 = -42; end
		18984: begin l_1 = +3;
				 l_2 = +43; end
		31885: begin l_1 = +3;
				 l_2 = -43; end
		18976: begin l_1 = -3;
				 l_2 = +43; end
		31877: begin l_1 = -3;
				 l_2 = -43; end
		37964: begin l_1 = +3;
				 l_2 = +44; end
		12905: begin l_1 = +3;
				 l_2 = -44; end
		37956: begin l_1 = -3;
				 l_2 = +44; end
		12897: begin l_1 = -3;
				 l_2 = -44; end
		25063: begin l_1 = +3;
				 l_2 = +45; end
		25806: begin l_1 = +3;
				 l_2 = -45; end
		25055: begin l_1 = -3;
				 l_2 = +45; end
		25798: begin l_1 = -3;
				 l_2 = -45; end
		50122: begin l_1 = +3;
				 l_2 = +46; end
		747: begin l_1 = +3;
				 l_2 = -46; end
		50114: begin l_1 = -3;
				 l_2 = +46; end
		739: begin l_1 = -3;
				 l_2 = -46; end
		49379: begin l_1 = +3;
				 l_2 = +47; end
		1490: begin l_1 = +3;
				 l_2 = -47; end
		49371: begin l_1 = -3;
				 l_2 = +47; end
		1482: begin l_1 = -3;
				 l_2 = -47; end
		47893: begin l_1 = +3;
				 l_2 = +48; end
		2976: begin l_1 = +3;
				 l_2 = -48; end
		47885: begin l_1 = -3;
				 l_2 = +48; end
		2968: begin l_1 = -3;
				 l_2 = -48; end
		44921: begin l_1 = +3;
				 l_2 = +49; end
		5948: begin l_1 = +3;
				 l_2 = -49; end
		44913: begin l_1 = -3;
				 l_2 = +49; end
		5940: begin l_1 = -3;
				 l_2 = -49; end
		38977: begin l_1 = +3;
				 l_2 = +50; end
		11892: begin l_1 = +3;
				 l_2 = -50; end
		38969: begin l_1 = -3;
				 l_2 = +50; end
		11884: begin l_1 = -3;
				 l_2 = -50; end
		27089: begin l_1 = +3;
				 l_2 = +51; end
		23780: begin l_1 = +3;
				 l_2 = -51; end
		27081: begin l_1 = -3;
				 l_2 = +51; end
		23772: begin l_1 = -3;
				 l_2 = -51; end
		3313: begin l_1 = +3;
				 l_2 = +52; end
		47556: begin l_1 = +3;
				 l_2 = -52; end
		3305: begin l_1 = -3;
				 l_2 = +52; end
		47548: begin l_1 = -3;
				 l_2 = -52; end
		6622: begin l_1 = +3;
				 l_2 = +53; end
		44247: begin l_1 = +3;
				 l_2 = -53; end
		6614: begin l_1 = -3;
				 l_2 = +53; end
		44239: begin l_1 = -3;
				 l_2 = -53; end
		13240: begin l_1 = +3;
				 l_2 = +54; end
		37629: begin l_1 = +3;
				 l_2 = -54; end
		13232: begin l_1 = -3;
				 l_2 = +54; end
		37621: begin l_1 = -3;
				 l_2 = -54; end
		26476: begin l_1 = +3;
				 l_2 = +55; end
		24393: begin l_1 = +3;
				 l_2 = -55; end
		26468: begin l_1 = -3;
				 l_2 = +55; end
		24385: begin l_1 = -3;
				 l_2 = -55; end
		2087: begin l_1 = +3;
				 l_2 = +56; end
		48782: begin l_1 = +3;
				 l_2 = -56; end
		2079: begin l_1 = -3;
				 l_2 = +56; end
		48774: begin l_1 = -3;
				 l_2 = -56; end
		4170: begin l_1 = +3;
				 l_2 = +57; end
		46699: begin l_1 = +3;
				 l_2 = -57; end
		4162: begin l_1 = -3;
				 l_2 = +57; end
		46691: begin l_1 = -3;
				 l_2 = -57; end
		8336: begin l_1 = +3;
				 l_2 = +58; end
		42533: begin l_1 = +3;
				 l_2 = -58; end
		8328: begin l_1 = -3;
				 l_2 = +58; end
		42525: begin l_1 = -3;
				 l_2 = -58; end
		16668: begin l_1 = +3;
				 l_2 = +59; end
		34201: begin l_1 = +3;
				 l_2 = -59; end
		16660: begin l_1 = -3;
				 l_2 = +59; end
		34193: begin l_1 = -3;
				 l_2 = -59; end
		33332: begin l_1 = +3;
				 l_2 = +60; end
		17537: begin l_1 = +3;
				 l_2 = -60; end
		33324: begin l_1 = -3;
				 l_2 = +60; end
		17529: begin l_1 = -3;
				 l_2 = -60; end
		15799: begin l_1 = +3;
				 l_2 = +61; end
		35070: begin l_1 = +3;
				 l_2 = -61; end
		15791: begin l_1 = -3;
				 l_2 = +61; end
		35062: begin l_1 = -3;
				 l_2 = -61; end
		31594: begin l_1 = +3;
				 l_2 = +62; end
		19275: begin l_1 = +3;
				 l_2 = -62; end
		31586: begin l_1 = -3;
				 l_2 = +62; end
		19267: begin l_1 = -3;
				 l_2 = -62; end
		12323: begin l_1 = +3;
				 l_2 = +63; end
		38546: begin l_1 = +3;
				 l_2 = -63; end
		12315: begin l_1 = -3;
				 l_2 = +63; end
		38538: begin l_1 = -3;
				 l_2 = -63; end
		24642: begin l_1 = +3;
				 l_2 = +64; end
		26227: begin l_1 = +3;
				 l_2 = -64; end
		24634: begin l_1 = -3;
				 l_2 = +64; end
		26219: begin l_1 = -3;
				 l_2 = -64; end
		49280: begin l_1 = +3;
				 l_2 = +65; end
		1589: begin l_1 = +3;
				 l_2 = -65; end
		49272: begin l_1 = -3;
				 l_2 = +65; end
		1581: begin l_1 = -3;
				 l_2 = -65; end
		47695: begin l_1 = +3;
				 l_2 = +66; end
		3174: begin l_1 = +3;
				 l_2 = -66; end
		47687: begin l_1 = -3;
				 l_2 = +66; end
		3166: begin l_1 = -3;
				 l_2 = -66; end
		44525: begin l_1 = +3;
				 l_2 = +67; end
		6344: begin l_1 = +3;
				 l_2 = -67; end
		44517: begin l_1 = -3;
				 l_2 = +67; end
		6336: begin l_1 = -3;
				 l_2 = -67; end
		38185: begin l_1 = +3;
				 l_2 = +68; end
		12684: begin l_1 = +3;
				 l_2 = -68; end
		38177: begin l_1 = -3;
				 l_2 = +68; end
		12676: begin l_1 = -3;
				 l_2 = -68; end
		24: begin l_1 = -4;
				 l_2 = +6; end
		50837: begin l_1 = -4;
				 l_2 = -5; end
		40: begin l_1 = +4;
				 l_2 = +6; end
		50821: begin l_1 = -4;
				 l_2 = -6; end
		72: begin l_1 = +4;
				 l_2 = +7; end
		50805: begin l_1 = +4;
				 l_2 = -7; end
		56: begin l_1 = -4;
				 l_2 = +7; end
		50789: begin l_1 = -4;
				 l_2 = -7; end
		136: begin l_1 = +4;
				 l_2 = +8; end
		50741: begin l_1 = +4;
				 l_2 = -8; end
		120: begin l_1 = -4;
				 l_2 = +8; end
		50725: begin l_1 = -4;
				 l_2 = -8; end
		264: begin l_1 = +4;
				 l_2 = +9; end
		50613: begin l_1 = +4;
				 l_2 = -9; end
		248: begin l_1 = -4;
				 l_2 = +9; end
		50597: begin l_1 = -4;
				 l_2 = -9; end
		520: begin l_1 = +4;
				 l_2 = +10; end
		50357: begin l_1 = +4;
				 l_2 = -10; end
		504: begin l_1 = -4;
				 l_2 = +10; end
		50341: begin l_1 = -4;
				 l_2 = -10; end
		1032: begin l_1 = +4;
				 l_2 = +11; end
		49845: begin l_1 = +4;
				 l_2 = -11; end
		1016: begin l_1 = -4;
				 l_2 = +11; end
		49829: begin l_1 = -4;
				 l_2 = -11; end
		2056: begin l_1 = +4;
				 l_2 = +12; end
		48821: begin l_1 = +4;
				 l_2 = -12; end
		2040: begin l_1 = -4;
				 l_2 = +12; end
		48805: begin l_1 = -4;
				 l_2 = -12; end
		4104: begin l_1 = +4;
				 l_2 = +13; end
		46773: begin l_1 = +4;
				 l_2 = -13; end
		4088: begin l_1 = -4;
				 l_2 = +13; end
		46757: begin l_1 = -4;
				 l_2 = -13; end
		8200: begin l_1 = +4;
				 l_2 = +14; end
		42677: begin l_1 = +4;
				 l_2 = -14; end
		8184: begin l_1 = -4;
				 l_2 = +14; end
		42661: begin l_1 = -4;
				 l_2 = -14; end
		16392: begin l_1 = +4;
				 l_2 = +15; end
		34485: begin l_1 = +4;
				 l_2 = -15; end
		16376: begin l_1 = -4;
				 l_2 = +15; end
		34469: begin l_1 = -4;
				 l_2 = -15; end
		32776: begin l_1 = +4;
				 l_2 = +16; end
		18101: begin l_1 = +4;
				 l_2 = -16; end
		32760: begin l_1 = -4;
				 l_2 = +16; end
		18085: begin l_1 = -4;
				 l_2 = -16; end
		14683: begin l_1 = +4;
				 l_2 = +17; end
		36194: begin l_1 = +4;
				 l_2 = -17; end
		14667: begin l_1 = -4;
				 l_2 = +17; end
		36178: begin l_1 = -4;
				 l_2 = -17; end
		29358: begin l_1 = +4;
				 l_2 = +18; end
		21519: begin l_1 = +4;
				 l_2 = -18; end
		29342: begin l_1 = -4;
				 l_2 = +18; end
		21503: begin l_1 = -4;
				 l_2 = -18; end
		7847: begin l_1 = +4;
				 l_2 = +19; end
		43030: begin l_1 = +4;
				 l_2 = -19; end
		7831: begin l_1 = -4;
				 l_2 = +19; end
		43014: begin l_1 = -4;
				 l_2 = -19; end
		15686: begin l_1 = +4;
				 l_2 = +20; end
		35191: begin l_1 = +4;
				 l_2 = -20; end
		15670: begin l_1 = -4;
				 l_2 = +20; end
		35175: begin l_1 = -4;
				 l_2 = -20; end
		31364: begin l_1 = +4;
				 l_2 = +21; end
		19513: begin l_1 = +4;
				 l_2 = -21; end
		31348: begin l_1 = -4;
				 l_2 = +21; end
		19497: begin l_1 = -4;
				 l_2 = -21; end
		11859: begin l_1 = +4;
				 l_2 = +22; end
		39018: begin l_1 = +4;
				 l_2 = -22; end
		11843: begin l_1 = -4;
				 l_2 = +22; end
		39002: begin l_1 = -4;
				 l_2 = -22; end
		23710: begin l_1 = +4;
				 l_2 = +23; end
		27167: begin l_1 = +4;
				 l_2 = -23; end
		23694: begin l_1 = -4;
				 l_2 = +23; end
		27151: begin l_1 = -4;
				 l_2 = -23; end
		47412: begin l_1 = +4;
				 l_2 = +24; end
		3465: begin l_1 = +4;
				 l_2 = -24; end
		47396: begin l_1 = -4;
				 l_2 = +24; end
		3449: begin l_1 = -4;
				 l_2 = -24; end
		43955: begin l_1 = +4;
				 l_2 = +25; end
		6922: begin l_1 = +4;
				 l_2 = -25; end
		43939: begin l_1 = -4;
				 l_2 = +25; end
		6906: begin l_1 = -4;
				 l_2 = -25; end
		37041: begin l_1 = +4;
				 l_2 = +26; end
		13836: begin l_1 = +4;
				 l_2 = -26; end
		37025: begin l_1 = -4;
				 l_2 = +26; end
		13820: begin l_1 = -4;
				 l_2 = -26; end
		23213: begin l_1 = +4;
				 l_2 = +27; end
		27664: begin l_1 = +4;
				 l_2 = -27; end
		23197: begin l_1 = -4;
				 l_2 = +27; end
		27648: begin l_1 = -4;
				 l_2 = -27; end
		46418: begin l_1 = +4;
				 l_2 = +28; end
		4459: begin l_1 = +4;
				 l_2 = -28; end
		46402: begin l_1 = -4;
				 l_2 = +28; end
		4443: begin l_1 = -4;
				 l_2 = -28; end
		41967: begin l_1 = +4;
				 l_2 = +29; end
		8910: begin l_1 = +4;
				 l_2 = -29; end
		41951: begin l_1 = -4;
				 l_2 = +29; end
		8894: begin l_1 = -4;
				 l_2 = -29; end
		33065: begin l_1 = +4;
				 l_2 = +30; end
		17812: begin l_1 = +4;
				 l_2 = -30; end
		33049: begin l_1 = -4;
				 l_2 = +30; end
		17796: begin l_1 = -4;
				 l_2 = -30; end
		15261: begin l_1 = +4;
				 l_2 = +31; end
		35616: begin l_1 = +4;
				 l_2 = -31; end
		15245: begin l_1 = -4;
				 l_2 = +31; end
		35600: begin l_1 = -4;
				 l_2 = -31; end
		30514: begin l_1 = +4;
				 l_2 = +32; end
		20363: begin l_1 = +4;
				 l_2 = -32; end
		30498: begin l_1 = -4;
				 l_2 = +32; end
		20347: begin l_1 = -4;
				 l_2 = -32; end
		10159: begin l_1 = +4;
				 l_2 = +33; end
		40718: begin l_1 = +4;
				 l_2 = -33; end
		10143: begin l_1 = -4;
				 l_2 = +33; end
		40702: begin l_1 = -4;
				 l_2 = -33; end
		20310: begin l_1 = +4;
				 l_2 = +34; end
		30567: begin l_1 = +4;
				 l_2 = -34; end
		20294: begin l_1 = -4;
				 l_2 = +34; end
		30551: begin l_1 = -4;
				 l_2 = -34; end
		40612: begin l_1 = +4;
				 l_2 = +35; end
		10265: begin l_1 = +4;
				 l_2 = -35; end
		40596: begin l_1 = -4;
				 l_2 = +35; end
		10249: begin l_1 = -4;
				 l_2 = -35; end
		30355: begin l_1 = +4;
				 l_2 = +36; end
		20522: begin l_1 = +4;
				 l_2 = -36; end
		30339: begin l_1 = -4;
				 l_2 = +36; end
		20506: begin l_1 = -4;
				 l_2 = -36; end
		9841: begin l_1 = +4;
				 l_2 = +37; end
		41036: begin l_1 = +4;
				 l_2 = -37; end
		9825: begin l_1 = -4;
				 l_2 = +37; end
		41020: begin l_1 = -4;
				 l_2 = -37; end
		19674: begin l_1 = +4;
				 l_2 = +38; end
		31203: begin l_1 = +4;
				 l_2 = -38; end
		19658: begin l_1 = -4;
				 l_2 = +38; end
		31187: begin l_1 = -4;
				 l_2 = -38; end
		39340: begin l_1 = +4;
				 l_2 = +39; end
		11537: begin l_1 = +4;
				 l_2 = -39; end
		39324: begin l_1 = -4;
				 l_2 = +39; end
		11521: begin l_1 = -4;
				 l_2 = -39; end
		27811: begin l_1 = +4;
				 l_2 = +40; end
		23066: begin l_1 = +4;
				 l_2 = -40; end
		27795: begin l_1 = -4;
				 l_2 = +40; end
		23050: begin l_1 = -4;
				 l_2 = -40; end
		4753: begin l_1 = +4;
				 l_2 = +41; end
		46124: begin l_1 = +4;
				 l_2 = -41; end
		4737: begin l_1 = -4;
				 l_2 = +41; end
		46108: begin l_1 = -4;
				 l_2 = -41; end
		9498: begin l_1 = +4;
				 l_2 = +42; end
		41379: begin l_1 = +4;
				 l_2 = -42; end
		9482: begin l_1 = -4;
				 l_2 = +42; end
		41363: begin l_1 = -4;
				 l_2 = -42; end
		18988: begin l_1 = +4;
				 l_2 = +43; end
		31889: begin l_1 = +4;
				 l_2 = -43; end
		18972: begin l_1 = -4;
				 l_2 = +43; end
		31873: begin l_1 = -4;
				 l_2 = -43; end
		37968: begin l_1 = +4;
				 l_2 = +44; end
		12909: begin l_1 = +4;
				 l_2 = -44; end
		37952: begin l_1 = -4;
				 l_2 = +44; end
		12893: begin l_1 = -4;
				 l_2 = -44; end
		25067: begin l_1 = +4;
				 l_2 = +45; end
		25810: begin l_1 = +4;
				 l_2 = -45; end
		25051: begin l_1 = -4;
				 l_2 = +45; end
		25794: begin l_1 = -4;
				 l_2 = -45; end
		50126: begin l_1 = +4;
				 l_2 = +46; end
		751: begin l_1 = +4;
				 l_2 = -46; end
		50110: begin l_1 = -4;
				 l_2 = +46; end
		735: begin l_1 = -4;
				 l_2 = -46; end
		49383: begin l_1 = +4;
				 l_2 = +47; end
		1494: begin l_1 = +4;
				 l_2 = -47; end
		49367: begin l_1 = -4;
				 l_2 = +47; end
		1478: begin l_1 = -4;
				 l_2 = -47; end
		47897: begin l_1 = +4;
				 l_2 = +48; end
		2980: begin l_1 = +4;
				 l_2 = -48; end
		47881: begin l_1 = -4;
				 l_2 = +48; end
		2964: begin l_1 = -4;
				 l_2 = -48; end
		44925: begin l_1 = +4;
				 l_2 = +49; end
		5952: begin l_1 = +4;
				 l_2 = -49; end
		44909: begin l_1 = -4;
				 l_2 = +49; end
		5936: begin l_1 = -4;
				 l_2 = -49; end
		38981: begin l_1 = +4;
				 l_2 = +50; end
		11896: begin l_1 = +4;
				 l_2 = -50; end
		38965: begin l_1 = -4;
				 l_2 = +50; end
		11880: begin l_1 = -4;
				 l_2 = -50; end
		27093: begin l_1 = +4;
				 l_2 = +51; end
		23784: begin l_1 = +4;
				 l_2 = -51; end
		27077: begin l_1 = -4;
				 l_2 = +51; end
		23768: begin l_1 = -4;
				 l_2 = -51; end
		3317: begin l_1 = +4;
				 l_2 = +52; end
		47560: begin l_1 = +4;
				 l_2 = -52; end
		3301: begin l_1 = -4;
				 l_2 = +52; end
		47544: begin l_1 = -4;
				 l_2 = -52; end
		6626: begin l_1 = +4;
				 l_2 = +53; end
		44251: begin l_1 = +4;
				 l_2 = -53; end
		6610: begin l_1 = -4;
				 l_2 = +53; end
		44235: begin l_1 = -4;
				 l_2 = -53; end
		13244: begin l_1 = +4;
				 l_2 = +54; end
		37633: begin l_1 = +4;
				 l_2 = -54; end
		13228: begin l_1 = -4;
				 l_2 = +54; end
		37617: begin l_1 = -4;
				 l_2 = -54; end
		26480: begin l_1 = +4;
				 l_2 = +55; end
		24397: begin l_1 = +4;
				 l_2 = -55; end
		26464: begin l_1 = -4;
				 l_2 = +55; end
		24381: begin l_1 = -4;
				 l_2 = -55; end
		2091: begin l_1 = +4;
				 l_2 = +56; end
		48786: begin l_1 = +4;
				 l_2 = -56; end
		2075: begin l_1 = -4;
				 l_2 = +56; end
		48770: begin l_1 = -4;
				 l_2 = -56; end
		4174: begin l_1 = +4;
				 l_2 = +57; end
		46703: begin l_1 = +4;
				 l_2 = -57; end
		4158: begin l_1 = -4;
				 l_2 = +57; end
		46687: begin l_1 = -4;
				 l_2 = -57; end
		8340: begin l_1 = +4;
				 l_2 = +58; end
		42537: begin l_1 = +4;
				 l_2 = -58; end
		8324: begin l_1 = -4;
				 l_2 = +58; end
		42521: begin l_1 = -4;
				 l_2 = -58; end
		16672: begin l_1 = +4;
				 l_2 = +59; end
		34205: begin l_1 = +4;
				 l_2 = -59; end
		16656: begin l_1 = -4;
				 l_2 = +59; end
		34189: begin l_1 = -4;
				 l_2 = -59; end
		33336: begin l_1 = +4;
				 l_2 = +60; end
		17541: begin l_1 = +4;
				 l_2 = -60; end
		33320: begin l_1 = -4;
				 l_2 = +60; end
		17525: begin l_1 = -4;
				 l_2 = -60; end
		15803: begin l_1 = +4;
				 l_2 = +61; end
		35074: begin l_1 = +4;
				 l_2 = -61; end
		15787: begin l_1 = -4;
				 l_2 = +61; end
		35058: begin l_1 = -4;
				 l_2 = -61; end
		31598: begin l_1 = +4;
				 l_2 = +62; end
		19279: begin l_1 = +4;
				 l_2 = -62; end
		31582: begin l_1 = -4;
				 l_2 = +62; end
		19263: begin l_1 = -4;
				 l_2 = -62; end
		12327: begin l_1 = +4;
				 l_2 = +63; end
		38550: begin l_1 = +4;
				 l_2 = -63; end
		12311: begin l_1 = -4;
				 l_2 = +63; end
		38534: begin l_1 = -4;
				 l_2 = -63; end
		24646: begin l_1 = +4;
				 l_2 = +64; end
		26231: begin l_1 = +4;
				 l_2 = -64; end
		24630: begin l_1 = -4;
				 l_2 = +64; end
		26215: begin l_1 = -4;
				 l_2 = -64; end
		49284: begin l_1 = +4;
				 l_2 = +65; end
		1593: begin l_1 = +4;
				 l_2 = -65; end
		49268: begin l_1 = -4;
				 l_2 = +65; end
		1577: begin l_1 = -4;
				 l_2 = -65; end
		47699: begin l_1 = +4;
				 l_2 = +66; end
		3178: begin l_1 = +4;
				 l_2 = -66; end
		47683: begin l_1 = -4;
				 l_2 = +66; end
		3162: begin l_1 = -4;
				 l_2 = -66; end
		44529: begin l_1 = +4;
				 l_2 = +67; end
		6348: begin l_1 = +4;
				 l_2 = -67; end
		44513: begin l_1 = -4;
				 l_2 = +67; end
		6332: begin l_1 = -4;
				 l_2 = -67; end
		38189: begin l_1 = +4;
				 l_2 = +68; end
		12688: begin l_1 = +4;
				 l_2 = -68; end
		38173: begin l_1 = -4;
				 l_2 = +68; end
		12672: begin l_1 = -4;
				 l_2 = -68; end
		48: begin l_1 = -5;
				 l_2 = +7; end
		50813: begin l_1 = -5;
				 l_2 = -6; end
		80: begin l_1 = +5;
				 l_2 = +7; end
		50781: begin l_1 = -5;
				 l_2 = -7; end
		144: begin l_1 = +5;
				 l_2 = +8; end
		50749: begin l_1 = +5;
				 l_2 = -8; end
		112: begin l_1 = -5;
				 l_2 = +8; end
		50717: begin l_1 = -5;
				 l_2 = -8; end
		272: begin l_1 = +5;
				 l_2 = +9; end
		50621: begin l_1 = +5;
				 l_2 = -9; end
		240: begin l_1 = -5;
				 l_2 = +9; end
		50589: begin l_1 = -5;
				 l_2 = -9; end
		528: begin l_1 = +5;
				 l_2 = +10; end
		50365: begin l_1 = +5;
				 l_2 = -10; end
		496: begin l_1 = -5;
				 l_2 = +10; end
		50333: begin l_1 = -5;
				 l_2 = -10; end
		1040: begin l_1 = +5;
				 l_2 = +11; end
		49853: begin l_1 = +5;
				 l_2 = -11; end
		1008: begin l_1 = -5;
				 l_2 = +11; end
		49821: begin l_1 = -5;
				 l_2 = -11; end
		2064: begin l_1 = +5;
				 l_2 = +12; end
		48829: begin l_1 = +5;
				 l_2 = -12; end
		2032: begin l_1 = -5;
				 l_2 = +12; end
		48797: begin l_1 = -5;
				 l_2 = -12; end
		4112: begin l_1 = +5;
				 l_2 = +13; end
		46781: begin l_1 = +5;
				 l_2 = -13; end
		4080: begin l_1 = -5;
				 l_2 = +13; end
		46749: begin l_1 = -5;
				 l_2 = -13; end
		8208: begin l_1 = +5;
				 l_2 = +14; end
		42685: begin l_1 = +5;
				 l_2 = -14; end
		8176: begin l_1 = -5;
				 l_2 = +14; end
		42653: begin l_1 = -5;
				 l_2 = -14; end
		16400: begin l_1 = +5;
				 l_2 = +15; end
		34493: begin l_1 = +5;
				 l_2 = -15; end
		16368: begin l_1 = -5;
				 l_2 = +15; end
		34461: begin l_1 = -5;
				 l_2 = -15; end
		32784: begin l_1 = +5;
				 l_2 = +16; end
		18109: begin l_1 = +5;
				 l_2 = -16; end
		32752: begin l_1 = -5;
				 l_2 = +16; end
		18077: begin l_1 = -5;
				 l_2 = -16; end
		14691: begin l_1 = +5;
				 l_2 = +17; end
		36202: begin l_1 = +5;
				 l_2 = -17; end
		14659: begin l_1 = -5;
				 l_2 = +17; end
		36170: begin l_1 = -5;
				 l_2 = -17; end
		29366: begin l_1 = +5;
				 l_2 = +18; end
		21527: begin l_1 = +5;
				 l_2 = -18; end
		29334: begin l_1 = -5;
				 l_2 = +18; end
		21495: begin l_1 = -5;
				 l_2 = -18; end
		7855: begin l_1 = +5;
				 l_2 = +19; end
		43038: begin l_1 = +5;
				 l_2 = -19; end
		7823: begin l_1 = -5;
				 l_2 = +19; end
		43006: begin l_1 = -5;
				 l_2 = -19; end
		15694: begin l_1 = +5;
				 l_2 = +20; end
		35199: begin l_1 = +5;
				 l_2 = -20; end
		15662: begin l_1 = -5;
				 l_2 = +20; end
		35167: begin l_1 = -5;
				 l_2 = -20; end
		31372: begin l_1 = +5;
				 l_2 = +21; end
		19521: begin l_1 = +5;
				 l_2 = -21; end
		31340: begin l_1 = -5;
				 l_2 = +21; end
		19489: begin l_1 = -5;
				 l_2 = -21; end
		11867: begin l_1 = +5;
				 l_2 = +22; end
		39026: begin l_1 = +5;
				 l_2 = -22; end
		11835: begin l_1 = -5;
				 l_2 = +22; end
		38994: begin l_1 = -5;
				 l_2 = -22; end
		23718: begin l_1 = +5;
				 l_2 = +23; end
		27175: begin l_1 = +5;
				 l_2 = -23; end
		23686: begin l_1 = -5;
				 l_2 = +23; end
		27143: begin l_1 = -5;
				 l_2 = -23; end
		47420: begin l_1 = +5;
				 l_2 = +24; end
		3473: begin l_1 = +5;
				 l_2 = -24; end
		47388: begin l_1 = -5;
				 l_2 = +24; end
		3441: begin l_1 = -5;
				 l_2 = -24; end
		43963: begin l_1 = +5;
				 l_2 = +25; end
		6930: begin l_1 = +5;
				 l_2 = -25; end
		43931: begin l_1 = -5;
				 l_2 = +25; end
		6898: begin l_1 = -5;
				 l_2 = -25; end
		37049: begin l_1 = +5;
				 l_2 = +26; end
		13844: begin l_1 = +5;
				 l_2 = -26; end
		37017: begin l_1 = -5;
				 l_2 = +26; end
		13812: begin l_1 = -5;
				 l_2 = -26; end
		23221: begin l_1 = +5;
				 l_2 = +27; end
		27672: begin l_1 = +5;
				 l_2 = -27; end
		23189: begin l_1 = -5;
				 l_2 = +27; end
		27640: begin l_1 = -5;
				 l_2 = -27; end
		46426: begin l_1 = +5;
				 l_2 = +28; end
		4467: begin l_1 = +5;
				 l_2 = -28; end
		46394: begin l_1 = -5;
				 l_2 = +28; end
		4435: begin l_1 = -5;
				 l_2 = -28; end
		41975: begin l_1 = +5;
				 l_2 = +29; end
		8918: begin l_1 = +5;
				 l_2 = -29; end
		41943: begin l_1 = -5;
				 l_2 = +29; end
		8886: begin l_1 = -5;
				 l_2 = -29; end
		33073: begin l_1 = +5;
				 l_2 = +30; end
		17820: begin l_1 = +5;
				 l_2 = -30; end
		33041: begin l_1 = -5;
				 l_2 = +30; end
		17788: begin l_1 = -5;
				 l_2 = -30; end
		15269: begin l_1 = +5;
				 l_2 = +31; end
		35624: begin l_1 = +5;
				 l_2 = -31; end
		15237: begin l_1 = -5;
				 l_2 = +31; end
		35592: begin l_1 = -5;
				 l_2 = -31; end
		30522: begin l_1 = +5;
				 l_2 = +32; end
		20371: begin l_1 = +5;
				 l_2 = -32; end
		30490: begin l_1 = -5;
				 l_2 = +32; end
		20339: begin l_1 = -5;
				 l_2 = -32; end
		10167: begin l_1 = +5;
				 l_2 = +33; end
		40726: begin l_1 = +5;
				 l_2 = -33; end
		10135: begin l_1 = -5;
				 l_2 = +33; end
		40694: begin l_1 = -5;
				 l_2 = -33; end
		20318: begin l_1 = +5;
				 l_2 = +34; end
		30575: begin l_1 = +5;
				 l_2 = -34; end
		20286: begin l_1 = -5;
				 l_2 = +34; end
		30543: begin l_1 = -5;
				 l_2 = -34; end
		40620: begin l_1 = +5;
				 l_2 = +35; end
		10273: begin l_1 = +5;
				 l_2 = -35; end
		40588: begin l_1 = -5;
				 l_2 = +35; end
		10241: begin l_1 = -5;
				 l_2 = -35; end
		30363: begin l_1 = +5;
				 l_2 = +36; end
		20530: begin l_1 = +5;
				 l_2 = -36; end
		30331: begin l_1 = -5;
				 l_2 = +36; end
		20498: begin l_1 = -5;
				 l_2 = -36; end
		9849: begin l_1 = +5;
				 l_2 = +37; end
		41044: begin l_1 = +5;
				 l_2 = -37; end
		9817: begin l_1 = -5;
				 l_2 = +37; end
		41012: begin l_1 = -5;
				 l_2 = -37; end
		19682: begin l_1 = +5;
				 l_2 = +38; end
		31211: begin l_1 = +5;
				 l_2 = -38; end
		19650: begin l_1 = -5;
				 l_2 = +38; end
		31179: begin l_1 = -5;
				 l_2 = -38; end
		39348: begin l_1 = +5;
				 l_2 = +39; end
		11545: begin l_1 = +5;
				 l_2 = -39; end
		39316: begin l_1 = -5;
				 l_2 = +39; end
		11513: begin l_1 = -5;
				 l_2 = -39; end
		27819: begin l_1 = +5;
				 l_2 = +40; end
		23074: begin l_1 = +5;
				 l_2 = -40; end
		27787: begin l_1 = -5;
				 l_2 = +40; end
		23042: begin l_1 = -5;
				 l_2 = -40; end
		4761: begin l_1 = +5;
				 l_2 = +41; end
		46132: begin l_1 = +5;
				 l_2 = -41; end
		4729: begin l_1 = -5;
				 l_2 = +41; end
		46100: begin l_1 = -5;
				 l_2 = -41; end
		9506: begin l_1 = +5;
				 l_2 = +42; end
		41387: begin l_1 = +5;
				 l_2 = -42; end
		9474: begin l_1 = -5;
				 l_2 = +42; end
		41355: begin l_1 = -5;
				 l_2 = -42; end
		18996: begin l_1 = +5;
				 l_2 = +43; end
		31897: begin l_1 = +5;
				 l_2 = -43; end
		18964: begin l_1 = -5;
				 l_2 = +43; end
		31865: begin l_1 = -5;
				 l_2 = -43; end
		37976: begin l_1 = +5;
				 l_2 = +44; end
		12917: begin l_1 = +5;
				 l_2 = -44; end
		37944: begin l_1 = -5;
				 l_2 = +44; end
		12885: begin l_1 = -5;
				 l_2 = -44; end
		25075: begin l_1 = +5;
				 l_2 = +45; end
		25818: begin l_1 = +5;
				 l_2 = -45; end
		25043: begin l_1 = -5;
				 l_2 = +45; end
		25786: begin l_1 = -5;
				 l_2 = -45; end
		50134: begin l_1 = +5;
				 l_2 = +46; end
		759: begin l_1 = +5;
				 l_2 = -46; end
		50102: begin l_1 = -5;
				 l_2 = +46; end
		727: begin l_1 = -5;
				 l_2 = -46; end
		49391: begin l_1 = +5;
				 l_2 = +47; end
		1502: begin l_1 = +5;
				 l_2 = -47; end
		49359: begin l_1 = -5;
				 l_2 = +47; end
		1470: begin l_1 = -5;
				 l_2 = -47; end
		47905: begin l_1 = +5;
				 l_2 = +48; end
		2988: begin l_1 = +5;
				 l_2 = -48; end
		47873: begin l_1 = -5;
				 l_2 = +48; end
		2956: begin l_1 = -5;
				 l_2 = -48; end
		44933: begin l_1 = +5;
				 l_2 = +49; end
		5960: begin l_1 = +5;
				 l_2 = -49; end
		44901: begin l_1 = -5;
				 l_2 = +49; end
		5928: begin l_1 = -5;
				 l_2 = -49; end
		38989: begin l_1 = +5;
				 l_2 = +50; end
		11904: begin l_1 = +5;
				 l_2 = -50; end
		38957: begin l_1 = -5;
				 l_2 = +50; end
		11872: begin l_1 = -5;
				 l_2 = -50; end
		27101: begin l_1 = +5;
				 l_2 = +51; end
		23792: begin l_1 = +5;
				 l_2 = -51; end
		27069: begin l_1 = -5;
				 l_2 = +51; end
		23760: begin l_1 = -5;
				 l_2 = -51; end
		3325: begin l_1 = +5;
				 l_2 = +52; end
		47568: begin l_1 = +5;
				 l_2 = -52; end
		3293: begin l_1 = -5;
				 l_2 = +52; end
		47536: begin l_1 = -5;
				 l_2 = -52; end
		6634: begin l_1 = +5;
				 l_2 = +53; end
		44259: begin l_1 = +5;
				 l_2 = -53; end
		6602: begin l_1 = -5;
				 l_2 = +53; end
		44227: begin l_1 = -5;
				 l_2 = -53; end
		13252: begin l_1 = +5;
				 l_2 = +54; end
		37641: begin l_1 = +5;
				 l_2 = -54; end
		13220: begin l_1 = -5;
				 l_2 = +54; end
		37609: begin l_1 = -5;
				 l_2 = -54; end
		26488: begin l_1 = +5;
				 l_2 = +55; end
		24405: begin l_1 = +5;
				 l_2 = -55; end
		26456: begin l_1 = -5;
				 l_2 = +55; end
		24373: begin l_1 = -5;
				 l_2 = -55; end
		2099: begin l_1 = +5;
				 l_2 = +56; end
		48794: begin l_1 = +5;
				 l_2 = -56; end
		2067: begin l_1 = -5;
				 l_2 = +56; end
		48762: begin l_1 = -5;
				 l_2 = -56; end
		4182: begin l_1 = +5;
				 l_2 = +57; end
		46711: begin l_1 = +5;
				 l_2 = -57; end
		4150: begin l_1 = -5;
				 l_2 = +57; end
		46679: begin l_1 = -5;
				 l_2 = -57; end
		8348: begin l_1 = +5;
				 l_2 = +58; end
		42545: begin l_1 = +5;
				 l_2 = -58; end
		8316: begin l_1 = -5;
				 l_2 = +58; end
		42513: begin l_1 = -5;
				 l_2 = -58; end
		16680: begin l_1 = +5;
				 l_2 = +59; end
		34213: begin l_1 = +5;
				 l_2 = -59; end
		16648: begin l_1 = -5;
				 l_2 = +59; end
		34181: begin l_1 = -5;
				 l_2 = -59; end
		33344: begin l_1 = +5;
				 l_2 = +60; end
		17549: begin l_1 = +5;
				 l_2 = -60; end
		33312: begin l_1 = -5;
				 l_2 = +60; end
		17517: begin l_1 = -5;
				 l_2 = -60; end
		15811: begin l_1 = +5;
				 l_2 = +61; end
		35082: begin l_1 = +5;
				 l_2 = -61; end
		15779: begin l_1 = -5;
				 l_2 = +61; end
		35050: begin l_1 = -5;
				 l_2 = -61; end
		31606: begin l_1 = +5;
				 l_2 = +62; end
		19287: begin l_1 = +5;
				 l_2 = -62; end
		31574: begin l_1 = -5;
				 l_2 = +62; end
		19255: begin l_1 = -5;
				 l_2 = -62; end
		12335: begin l_1 = +5;
				 l_2 = +63; end
		38558: begin l_1 = +5;
				 l_2 = -63; end
		12303: begin l_1 = -5;
				 l_2 = +63; end
		38526: begin l_1 = -5;
				 l_2 = -63; end
		24654: begin l_1 = +5;
				 l_2 = +64; end
		26239: begin l_1 = +5;
				 l_2 = -64; end
		24622: begin l_1 = -5;
				 l_2 = +64; end
		26207: begin l_1 = -5;
				 l_2 = -64; end
		49292: begin l_1 = +5;
				 l_2 = +65; end
		1601: begin l_1 = +5;
				 l_2 = -65; end
		49260: begin l_1 = -5;
				 l_2 = +65; end
		1569: begin l_1 = -5;
				 l_2 = -65; end
		47707: begin l_1 = +5;
				 l_2 = +66; end
		3186: begin l_1 = +5;
				 l_2 = -66; end
		47675: begin l_1 = -5;
				 l_2 = +66; end
		3154: begin l_1 = -5;
				 l_2 = -66; end
		44537: begin l_1 = +5;
				 l_2 = +67; end
		6356: begin l_1 = +5;
				 l_2 = -67; end
		44505: begin l_1 = -5;
				 l_2 = +67; end
		6324: begin l_1 = -5;
				 l_2 = -67; end
		38197: begin l_1 = +5;
				 l_2 = +68; end
		12696: begin l_1 = +5;
				 l_2 = -68; end
		38165: begin l_1 = -5;
				 l_2 = +68; end
		12664: begin l_1 = -5;
				 l_2 = -68; end
		96: begin l_1 = -6;
				 l_2 = +8; end
		50765: begin l_1 = -6;
				 l_2 = -7; end
		160: begin l_1 = +6;
				 l_2 = +8; end
		50701: begin l_1 = -6;
				 l_2 = -8; end
		288: begin l_1 = +6;
				 l_2 = +9; end
		50637: begin l_1 = +6;
				 l_2 = -9; end
		224: begin l_1 = -6;
				 l_2 = +9; end
		50573: begin l_1 = -6;
				 l_2 = -9; end
		544: begin l_1 = +6;
				 l_2 = +10; end
		50381: begin l_1 = +6;
				 l_2 = -10; end
		480: begin l_1 = -6;
				 l_2 = +10; end
		50317: begin l_1 = -6;
				 l_2 = -10; end
		1056: begin l_1 = +6;
				 l_2 = +11; end
		49869: begin l_1 = +6;
				 l_2 = -11; end
		992: begin l_1 = -6;
				 l_2 = +11; end
		49805: begin l_1 = -6;
				 l_2 = -11; end
		2080: begin l_1 = +6;
				 l_2 = +12; end
		48845: begin l_1 = +6;
				 l_2 = -12; end
		2016: begin l_1 = -6;
				 l_2 = +12; end
		48781: begin l_1 = -6;
				 l_2 = -12; end
		4128: begin l_1 = +6;
				 l_2 = +13; end
		46797: begin l_1 = +6;
				 l_2 = -13; end
		4064: begin l_1 = -6;
				 l_2 = +13; end
		46733: begin l_1 = -6;
				 l_2 = -13; end
		8224: begin l_1 = +6;
				 l_2 = +14; end
		42701: begin l_1 = +6;
				 l_2 = -14; end
		8160: begin l_1 = -6;
				 l_2 = +14; end
		42637: begin l_1 = -6;
				 l_2 = -14; end
		16416: begin l_1 = +6;
				 l_2 = +15; end
		34509: begin l_1 = +6;
				 l_2 = -15; end
		16352: begin l_1 = -6;
				 l_2 = +15; end
		34445: begin l_1 = -6;
				 l_2 = -15; end
		32800: begin l_1 = +6;
				 l_2 = +16; end
		18125: begin l_1 = +6;
				 l_2 = -16; end
		32736: begin l_1 = -6;
				 l_2 = +16; end
		18061: begin l_1 = -6;
				 l_2 = -16; end
		14707: begin l_1 = +6;
				 l_2 = +17; end
		36218: begin l_1 = +6;
				 l_2 = -17; end
		14643: begin l_1 = -6;
				 l_2 = +17; end
		36154: begin l_1 = -6;
				 l_2 = -17; end
		29382: begin l_1 = +6;
				 l_2 = +18; end
		21543: begin l_1 = +6;
				 l_2 = -18; end
		29318: begin l_1 = -6;
				 l_2 = +18; end
		21479: begin l_1 = -6;
				 l_2 = -18; end
		7871: begin l_1 = +6;
				 l_2 = +19; end
		43054: begin l_1 = +6;
				 l_2 = -19; end
		7807: begin l_1 = -6;
				 l_2 = +19; end
		42990: begin l_1 = -6;
				 l_2 = -19; end
		15710: begin l_1 = +6;
				 l_2 = +20; end
		35215: begin l_1 = +6;
				 l_2 = -20; end
		15646: begin l_1 = -6;
				 l_2 = +20; end
		35151: begin l_1 = -6;
				 l_2 = -20; end
		31388: begin l_1 = +6;
				 l_2 = +21; end
		19537: begin l_1 = +6;
				 l_2 = -21; end
		31324: begin l_1 = -6;
				 l_2 = +21; end
		19473: begin l_1 = -6;
				 l_2 = -21; end
		11883: begin l_1 = +6;
				 l_2 = +22; end
		39042: begin l_1 = +6;
				 l_2 = -22; end
		11819: begin l_1 = -6;
				 l_2 = +22; end
		38978: begin l_1 = -6;
				 l_2 = -22; end
		23734: begin l_1 = +6;
				 l_2 = +23; end
		27191: begin l_1 = +6;
				 l_2 = -23; end
		23670: begin l_1 = -6;
				 l_2 = +23; end
		27127: begin l_1 = -6;
				 l_2 = -23; end
		47436: begin l_1 = +6;
				 l_2 = +24; end
		3489: begin l_1 = +6;
				 l_2 = -24; end
		47372: begin l_1 = -6;
				 l_2 = +24; end
		3425: begin l_1 = -6;
				 l_2 = -24; end
		43979: begin l_1 = +6;
				 l_2 = +25; end
		6946: begin l_1 = +6;
				 l_2 = -25; end
		43915: begin l_1 = -6;
				 l_2 = +25; end
		6882: begin l_1 = -6;
				 l_2 = -25; end
		37065: begin l_1 = +6;
				 l_2 = +26; end
		13860: begin l_1 = +6;
				 l_2 = -26; end
		37001: begin l_1 = -6;
				 l_2 = +26; end
		13796: begin l_1 = -6;
				 l_2 = -26; end
		23237: begin l_1 = +6;
				 l_2 = +27; end
		27688: begin l_1 = +6;
				 l_2 = -27; end
		23173: begin l_1 = -6;
				 l_2 = +27; end
		27624: begin l_1 = -6;
				 l_2 = -27; end
		46442: begin l_1 = +6;
				 l_2 = +28; end
		4483: begin l_1 = +6;
				 l_2 = -28; end
		46378: begin l_1 = -6;
				 l_2 = +28; end
		4419: begin l_1 = -6;
				 l_2 = -28; end
		41991: begin l_1 = +6;
				 l_2 = +29; end
		8934: begin l_1 = +6;
				 l_2 = -29; end
		41927: begin l_1 = -6;
				 l_2 = +29; end
		8870: begin l_1 = -6;
				 l_2 = -29; end
		33089: begin l_1 = +6;
				 l_2 = +30; end
		17836: begin l_1 = +6;
				 l_2 = -30; end
		33025: begin l_1 = -6;
				 l_2 = +30; end
		17772: begin l_1 = -6;
				 l_2 = -30; end
		15285: begin l_1 = +6;
				 l_2 = +31; end
		35640: begin l_1 = +6;
				 l_2 = -31; end
		15221: begin l_1 = -6;
				 l_2 = +31; end
		35576: begin l_1 = -6;
				 l_2 = -31; end
		30538: begin l_1 = +6;
				 l_2 = +32; end
		20387: begin l_1 = +6;
				 l_2 = -32; end
		30474: begin l_1 = -6;
				 l_2 = +32; end
		20323: begin l_1 = -6;
				 l_2 = -32; end
		10183: begin l_1 = +6;
				 l_2 = +33; end
		40742: begin l_1 = +6;
				 l_2 = -33; end
		10119: begin l_1 = -6;
				 l_2 = +33; end
		40678: begin l_1 = -6;
				 l_2 = -33; end
		20334: begin l_1 = +6;
				 l_2 = +34; end
		30591: begin l_1 = +6;
				 l_2 = -34; end
		20270: begin l_1 = -6;
				 l_2 = +34; end
		30527: begin l_1 = -6;
				 l_2 = -34; end
		40636: begin l_1 = +6;
				 l_2 = +35; end
		10289: begin l_1 = +6;
				 l_2 = -35; end
		40572: begin l_1 = -6;
				 l_2 = +35; end
		10225: begin l_1 = -6;
				 l_2 = -35; end
		30379: begin l_1 = +6;
				 l_2 = +36; end
		20546: begin l_1 = +6;
				 l_2 = -36; end
		30315: begin l_1 = -6;
				 l_2 = +36; end
		20482: begin l_1 = -6;
				 l_2 = -36; end
		9865: begin l_1 = +6;
				 l_2 = +37; end
		41060: begin l_1 = +6;
				 l_2 = -37; end
		9801: begin l_1 = -6;
				 l_2 = +37; end
		40996: begin l_1 = -6;
				 l_2 = -37; end
		19698: begin l_1 = +6;
				 l_2 = +38; end
		31227: begin l_1 = +6;
				 l_2 = -38; end
		19634: begin l_1 = -6;
				 l_2 = +38; end
		31163: begin l_1 = -6;
				 l_2 = -38; end
		39364: begin l_1 = +6;
				 l_2 = +39; end
		11561: begin l_1 = +6;
				 l_2 = -39; end
		39300: begin l_1 = -6;
				 l_2 = +39; end
		11497: begin l_1 = -6;
				 l_2 = -39; end
		27835: begin l_1 = +6;
				 l_2 = +40; end
		23090: begin l_1 = +6;
				 l_2 = -40; end
		27771: begin l_1 = -6;
				 l_2 = +40; end
		23026: begin l_1 = -6;
				 l_2 = -40; end
		4777: begin l_1 = +6;
				 l_2 = +41; end
		46148: begin l_1 = +6;
				 l_2 = -41; end
		4713: begin l_1 = -6;
				 l_2 = +41; end
		46084: begin l_1 = -6;
				 l_2 = -41; end
		9522: begin l_1 = +6;
				 l_2 = +42; end
		41403: begin l_1 = +6;
				 l_2 = -42; end
		9458: begin l_1 = -6;
				 l_2 = +42; end
		41339: begin l_1 = -6;
				 l_2 = -42; end
		19012: begin l_1 = +6;
				 l_2 = +43; end
		31913: begin l_1 = +6;
				 l_2 = -43; end
		18948: begin l_1 = -6;
				 l_2 = +43; end
		31849: begin l_1 = -6;
				 l_2 = -43; end
		37992: begin l_1 = +6;
				 l_2 = +44; end
		12933: begin l_1 = +6;
				 l_2 = -44; end
		37928: begin l_1 = -6;
				 l_2 = +44; end
		12869: begin l_1 = -6;
				 l_2 = -44; end
		25091: begin l_1 = +6;
				 l_2 = +45; end
		25834: begin l_1 = +6;
				 l_2 = -45; end
		25027: begin l_1 = -6;
				 l_2 = +45; end
		25770: begin l_1 = -6;
				 l_2 = -45; end
		50150: begin l_1 = +6;
				 l_2 = +46; end
		775: begin l_1 = +6;
				 l_2 = -46; end
		50086: begin l_1 = -6;
				 l_2 = +46; end
		711: begin l_1 = -6;
				 l_2 = -46; end
		49407: begin l_1 = +6;
				 l_2 = +47; end
		1518: begin l_1 = +6;
				 l_2 = -47; end
		49343: begin l_1 = -6;
				 l_2 = +47; end
		1454: begin l_1 = -6;
				 l_2 = -47; end
		47921: begin l_1 = +6;
				 l_2 = +48; end
		3004: begin l_1 = +6;
				 l_2 = -48; end
		47857: begin l_1 = -6;
				 l_2 = +48; end
		2940: begin l_1 = -6;
				 l_2 = -48; end
		44949: begin l_1 = +6;
				 l_2 = +49; end
		5976: begin l_1 = +6;
				 l_2 = -49; end
		44885: begin l_1 = -6;
				 l_2 = +49; end
		5912: begin l_1 = -6;
				 l_2 = -49; end
		39005: begin l_1 = +6;
				 l_2 = +50; end
		11920: begin l_1 = +6;
				 l_2 = -50; end
		38941: begin l_1 = -6;
				 l_2 = +50; end
		11856: begin l_1 = -6;
				 l_2 = -50; end
		27117: begin l_1 = +6;
				 l_2 = +51; end
		23808: begin l_1 = +6;
				 l_2 = -51; end
		27053: begin l_1 = -6;
				 l_2 = +51; end
		23744: begin l_1 = -6;
				 l_2 = -51; end
		3341: begin l_1 = +6;
				 l_2 = +52; end
		47584: begin l_1 = +6;
				 l_2 = -52; end
		3277: begin l_1 = -6;
				 l_2 = +52; end
		47520: begin l_1 = -6;
				 l_2 = -52; end
		6650: begin l_1 = +6;
				 l_2 = +53; end
		44275: begin l_1 = +6;
				 l_2 = -53; end
		6586: begin l_1 = -6;
				 l_2 = +53; end
		44211: begin l_1 = -6;
				 l_2 = -53; end
		13268: begin l_1 = +6;
				 l_2 = +54; end
		37657: begin l_1 = +6;
				 l_2 = -54; end
		13204: begin l_1 = -6;
				 l_2 = +54; end
		37593: begin l_1 = -6;
				 l_2 = -54; end
		26504: begin l_1 = +6;
				 l_2 = +55; end
		24421: begin l_1 = +6;
				 l_2 = -55; end
		26440: begin l_1 = -6;
				 l_2 = +55; end
		24357: begin l_1 = -6;
				 l_2 = -55; end
		2115: begin l_1 = +6;
				 l_2 = +56; end
		48810: begin l_1 = +6;
				 l_2 = -56; end
		2051: begin l_1 = -6;
				 l_2 = +56; end
		48746: begin l_1 = -6;
				 l_2 = -56; end
		4198: begin l_1 = +6;
				 l_2 = +57; end
		46727: begin l_1 = +6;
				 l_2 = -57; end
		4134: begin l_1 = -6;
				 l_2 = +57; end
		46663: begin l_1 = -6;
				 l_2 = -57; end
		8364: begin l_1 = +6;
				 l_2 = +58; end
		42561: begin l_1 = +6;
				 l_2 = -58; end
		8300: begin l_1 = -6;
				 l_2 = +58; end
		42497: begin l_1 = -6;
				 l_2 = -58; end
		16696: begin l_1 = +6;
				 l_2 = +59; end
		34229: begin l_1 = +6;
				 l_2 = -59; end
		16632: begin l_1 = -6;
				 l_2 = +59; end
		34165: begin l_1 = -6;
				 l_2 = -59; end
		33360: begin l_1 = +6;
				 l_2 = +60; end
		17565: begin l_1 = +6;
				 l_2 = -60; end
		33296: begin l_1 = -6;
				 l_2 = +60; end
		17501: begin l_1 = -6;
				 l_2 = -60; end
		15827: begin l_1 = +6;
				 l_2 = +61; end
		35098: begin l_1 = +6;
				 l_2 = -61; end
		15763: begin l_1 = -6;
				 l_2 = +61; end
		35034: begin l_1 = -6;
				 l_2 = -61; end
		31622: begin l_1 = +6;
				 l_2 = +62; end
		19303: begin l_1 = +6;
				 l_2 = -62; end
		31558: begin l_1 = -6;
				 l_2 = +62; end
		19239: begin l_1 = -6;
				 l_2 = -62; end
		12351: begin l_1 = +6;
				 l_2 = +63; end
		38574: begin l_1 = +6;
				 l_2 = -63; end
		12287: begin l_1 = -6;
				 l_2 = +63; end
		38510: begin l_1 = -6;
				 l_2 = -63; end
		24670: begin l_1 = +6;
				 l_2 = +64; end
		26255: begin l_1 = +6;
				 l_2 = -64; end
		24606: begin l_1 = -6;
				 l_2 = +64; end
		26191: begin l_1 = -6;
				 l_2 = -64; end
		49308: begin l_1 = +6;
				 l_2 = +65; end
		1617: begin l_1 = +6;
				 l_2 = -65; end
		49244: begin l_1 = -6;
				 l_2 = +65; end
		1553: begin l_1 = -6;
				 l_2 = -65; end
		47723: begin l_1 = +6;
				 l_2 = +66; end
		3202: begin l_1 = +6;
				 l_2 = -66; end
		47659: begin l_1 = -6;
				 l_2 = +66; end
		3138: begin l_1 = -6;
				 l_2 = -66; end
		44553: begin l_1 = +6;
				 l_2 = +67; end
		6372: begin l_1 = +6;
				 l_2 = -67; end
		44489: begin l_1 = -6;
				 l_2 = +67; end
		6308: begin l_1 = -6;
				 l_2 = -67; end
		38213: begin l_1 = +6;
				 l_2 = +68; end
		12712: begin l_1 = +6;
				 l_2 = -68; end
		38149: begin l_1 = -6;
				 l_2 = +68; end
		12648: begin l_1 = -6;
				 l_2 = -68; end
		192: begin l_1 = -7;
				 l_2 = +9; end
		50669: begin l_1 = -7;
				 l_2 = -8; end
		320: begin l_1 = +7;
				 l_2 = +9; end
		50541: begin l_1 = -7;
				 l_2 = -9; end
		576: begin l_1 = +7;
				 l_2 = +10; end
		50413: begin l_1 = +7;
				 l_2 = -10; end
		448: begin l_1 = -7;
				 l_2 = +10; end
		50285: begin l_1 = -7;
				 l_2 = -10; end
		1088: begin l_1 = +7;
				 l_2 = +11; end
		49901: begin l_1 = +7;
				 l_2 = -11; end
		960: begin l_1 = -7;
				 l_2 = +11; end
		49773: begin l_1 = -7;
				 l_2 = -11; end
		2112: begin l_1 = +7;
				 l_2 = +12; end
		48877: begin l_1 = +7;
				 l_2 = -12; end
		1984: begin l_1 = -7;
				 l_2 = +12; end
		48749: begin l_1 = -7;
				 l_2 = -12; end
		4160: begin l_1 = +7;
				 l_2 = +13; end
		46829: begin l_1 = +7;
				 l_2 = -13; end
		4032: begin l_1 = -7;
				 l_2 = +13; end
		46701: begin l_1 = -7;
				 l_2 = -13; end
		8256: begin l_1 = +7;
				 l_2 = +14; end
		42733: begin l_1 = +7;
				 l_2 = -14; end
		8128: begin l_1 = -7;
				 l_2 = +14; end
		42605: begin l_1 = -7;
				 l_2 = -14; end
		16448: begin l_1 = +7;
				 l_2 = +15; end
		34541: begin l_1 = +7;
				 l_2 = -15; end
		16320: begin l_1 = -7;
				 l_2 = +15; end
		34413: begin l_1 = -7;
				 l_2 = -15; end
		32832: begin l_1 = +7;
				 l_2 = +16; end
		18157: begin l_1 = +7;
				 l_2 = -16; end
		32704: begin l_1 = -7;
				 l_2 = +16; end
		18029: begin l_1 = -7;
				 l_2 = -16; end
		14739: begin l_1 = +7;
				 l_2 = +17; end
		36250: begin l_1 = +7;
				 l_2 = -17; end
		14611: begin l_1 = -7;
				 l_2 = +17; end
		36122: begin l_1 = -7;
				 l_2 = -17; end
		29414: begin l_1 = +7;
				 l_2 = +18; end
		21575: begin l_1 = +7;
				 l_2 = -18; end
		29286: begin l_1 = -7;
				 l_2 = +18; end
		21447: begin l_1 = -7;
				 l_2 = -18; end
		7903: begin l_1 = +7;
				 l_2 = +19; end
		43086: begin l_1 = +7;
				 l_2 = -19; end
		7775: begin l_1 = -7;
				 l_2 = +19; end
		42958: begin l_1 = -7;
				 l_2 = -19; end
		15742: begin l_1 = +7;
				 l_2 = +20; end
		35247: begin l_1 = +7;
				 l_2 = -20; end
		15614: begin l_1 = -7;
				 l_2 = +20; end
		35119: begin l_1 = -7;
				 l_2 = -20; end
		31420: begin l_1 = +7;
				 l_2 = +21; end
		19569: begin l_1 = +7;
				 l_2 = -21; end
		31292: begin l_1 = -7;
				 l_2 = +21; end
		19441: begin l_1 = -7;
				 l_2 = -21; end
		11915: begin l_1 = +7;
				 l_2 = +22; end
		39074: begin l_1 = +7;
				 l_2 = -22; end
		11787: begin l_1 = -7;
				 l_2 = +22; end
		38946: begin l_1 = -7;
				 l_2 = -22; end
		23766: begin l_1 = +7;
				 l_2 = +23; end
		27223: begin l_1 = +7;
				 l_2 = -23; end
		23638: begin l_1 = -7;
				 l_2 = +23; end
		27095: begin l_1 = -7;
				 l_2 = -23; end
		47468: begin l_1 = +7;
				 l_2 = +24; end
		3521: begin l_1 = +7;
				 l_2 = -24; end
		47340: begin l_1 = -7;
				 l_2 = +24; end
		3393: begin l_1 = -7;
				 l_2 = -24; end
		44011: begin l_1 = +7;
				 l_2 = +25; end
		6978: begin l_1 = +7;
				 l_2 = -25; end
		43883: begin l_1 = -7;
				 l_2 = +25; end
		6850: begin l_1 = -7;
				 l_2 = -25; end
		37097: begin l_1 = +7;
				 l_2 = +26; end
		13892: begin l_1 = +7;
				 l_2 = -26; end
		36969: begin l_1 = -7;
				 l_2 = +26; end
		13764: begin l_1 = -7;
				 l_2 = -26; end
		23269: begin l_1 = +7;
				 l_2 = +27; end
		27720: begin l_1 = +7;
				 l_2 = -27; end
		23141: begin l_1 = -7;
				 l_2 = +27; end
		27592: begin l_1 = -7;
				 l_2 = -27; end
		46474: begin l_1 = +7;
				 l_2 = +28; end
		4515: begin l_1 = +7;
				 l_2 = -28; end
		46346: begin l_1 = -7;
				 l_2 = +28; end
		4387: begin l_1 = -7;
				 l_2 = -28; end
		42023: begin l_1 = +7;
				 l_2 = +29; end
		8966: begin l_1 = +7;
				 l_2 = -29; end
		41895: begin l_1 = -7;
				 l_2 = +29; end
		8838: begin l_1 = -7;
				 l_2 = -29; end
		33121: begin l_1 = +7;
				 l_2 = +30; end
		17868: begin l_1 = +7;
				 l_2 = -30; end
		32993: begin l_1 = -7;
				 l_2 = +30; end
		17740: begin l_1 = -7;
				 l_2 = -30; end
		15317: begin l_1 = +7;
				 l_2 = +31; end
		35672: begin l_1 = +7;
				 l_2 = -31; end
		15189: begin l_1 = -7;
				 l_2 = +31; end
		35544: begin l_1 = -7;
				 l_2 = -31; end
		30570: begin l_1 = +7;
				 l_2 = +32; end
		20419: begin l_1 = +7;
				 l_2 = -32; end
		30442: begin l_1 = -7;
				 l_2 = +32; end
		20291: begin l_1 = -7;
				 l_2 = -32; end
		10215: begin l_1 = +7;
				 l_2 = +33; end
		40774: begin l_1 = +7;
				 l_2 = -33; end
		10087: begin l_1 = -7;
				 l_2 = +33; end
		40646: begin l_1 = -7;
				 l_2 = -33; end
		20366: begin l_1 = +7;
				 l_2 = +34; end
		30623: begin l_1 = +7;
				 l_2 = -34; end
		20238: begin l_1 = -7;
				 l_2 = +34; end
		30495: begin l_1 = -7;
				 l_2 = -34; end
		40668: begin l_1 = +7;
				 l_2 = +35; end
		10321: begin l_1 = +7;
				 l_2 = -35; end
		40540: begin l_1 = -7;
				 l_2 = +35; end
		10193: begin l_1 = -7;
				 l_2 = -35; end
		30411: begin l_1 = +7;
				 l_2 = +36; end
		20578: begin l_1 = +7;
				 l_2 = -36; end
		30283: begin l_1 = -7;
				 l_2 = +36; end
		20450: begin l_1 = -7;
				 l_2 = -36; end
		9897: begin l_1 = +7;
				 l_2 = +37; end
		41092: begin l_1 = +7;
				 l_2 = -37; end
		9769: begin l_1 = -7;
				 l_2 = +37; end
		40964: begin l_1 = -7;
				 l_2 = -37; end
		19730: begin l_1 = +7;
				 l_2 = +38; end
		31259: begin l_1 = +7;
				 l_2 = -38; end
		19602: begin l_1 = -7;
				 l_2 = +38; end
		31131: begin l_1 = -7;
				 l_2 = -38; end
		39396: begin l_1 = +7;
				 l_2 = +39; end
		11593: begin l_1 = +7;
				 l_2 = -39; end
		39268: begin l_1 = -7;
				 l_2 = +39; end
		11465: begin l_1 = -7;
				 l_2 = -39; end
		27867: begin l_1 = +7;
				 l_2 = +40; end
		23122: begin l_1 = +7;
				 l_2 = -40; end
		27739: begin l_1 = -7;
				 l_2 = +40; end
		22994: begin l_1 = -7;
				 l_2 = -40; end
		4809: begin l_1 = +7;
				 l_2 = +41; end
		46180: begin l_1 = +7;
				 l_2 = -41; end
		4681: begin l_1 = -7;
				 l_2 = +41; end
		46052: begin l_1 = -7;
				 l_2 = -41; end
		9554: begin l_1 = +7;
				 l_2 = +42; end
		41435: begin l_1 = +7;
				 l_2 = -42; end
		9426: begin l_1 = -7;
				 l_2 = +42; end
		41307: begin l_1 = -7;
				 l_2 = -42; end
		19044: begin l_1 = +7;
				 l_2 = +43; end
		31945: begin l_1 = +7;
				 l_2 = -43; end
		18916: begin l_1 = -7;
				 l_2 = +43; end
		31817: begin l_1 = -7;
				 l_2 = -43; end
		38024: begin l_1 = +7;
				 l_2 = +44; end
		12965: begin l_1 = +7;
				 l_2 = -44; end
		37896: begin l_1 = -7;
				 l_2 = +44; end
		12837: begin l_1 = -7;
				 l_2 = -44; end
		25123: begin l_1 = +7;
				 l_2 = +45; end
		25866: begin l_1 = +7;
				 l_2 = -45; end
		24995: begin l_1 = -7;
				 l_2 = +45; end
		25738: begin l_1 = -7;
				 l_2 = -45; end
		50182: begin l_1 = +7;
				 l_2 = +46; end
		807: begin l_1 = +7;
				 l_2 = -46; end
		50054: begin l_1 = -7;
				 l_2 = +46; end
		679: begin l_1 = -7;
				 l_2 = -46; end
		49439: begin l_1 = +7;
				 l_2 = +47; end
		1550: begin l_1 = +7;
				 l_2 = -47; end
		49311: begin l_1 = -7;
				 l_2 = +47; end
		1422: begin l_1 = -7;
				 l_2 = -47; end
		47953: begin l_1 = +7;
				 l_2 = +48; end
		3036: begin l_1 = +7;
				 l_2 = -48; end
		47825: begin l_1 = -7;
				 l_2 = +48; end
		2908: begin l_1 = -7;
				 l_2 = -48; end
		44981: begin l_1 = +7;
				 l_2 = +49; end
		6008: begin l_1 = +7;
				 l_2 = -49; end
		44853: begin l_1 = -7;
				 l_2 = +49; end
		5880: begin l_1 = -7;
				 l_2 = -49; end
		39037: begin l_1 = +7;
				 l_2 = +50; end
		11952: begin l_1 = +7;
				 l_2 = -50; end
		38909: begin l_1 = -7;
				 l_2 = +50; end
		11824: begin l_1 = -7;
				 l_2 = -50; end
		27149: begin l_1 = +7;
				 l_2 = +51; end
		23840: begin l_1 = +7;
				 l_2 = -51; end
		27021: begin l_1 = -7;
				 l_2 = +51; end
		23712: begin l_1 = -7;
				 l_2 = -51; end
		3373: begin l_1 = +7;
				 l_2 = +52; end
		47616: begin l_1 = +7;
				 l_2 = -52; end
		3245: begin l_1 = -7;
				 l_2 = +52; end
		47488: begin l_1 = -7;
				 l_2 = -52; end
		6682: begin l_1 = +7;
				 l_2 = +53; end
		44307: begin l_1 = +7;
				 l_2 = -53; end
		6554: begin l_1 = -7;
				 l_2 = +53; end
		44179: begin l_1 = -7;
				 l_2 = -53; end
		13300: begin l_1 = +7;
				 l_2 = +54; end
		37689: begin l_1 = +7;
				 l_2 = -54; end
		13172: begin l_1 = -7;
				 l_2 = +54; end
		37561: begin l_1 = -7;
				 l_2 = -54; end
		26536: begin l_1 = +7;
				 l_2 = +55; end
		24453: begin l_1 = +7;
				 l_2 = -55; end
		26408: begin l_1 = -7;
				 l_2 = +55; end
		24325: begin l_1 = -7;
				 l_2 = -55; end
		2147: begin l_1 = +7;
				 l_2 = +56; end
		48842: begin l_1 = +7;
				 l_2 = -56; end
		2019: begin l_1 = -7;
				 l_2 = +56; end
		48714: begin l_1 = -7;
				 l_2 = -56; end
		4230: begin l_1 = +7;
				 l_2 = +57; end
		46759: begin l_1 = +7;
				 l_2 = -57; end
		4102: begin l_1 = -7;
				 l_2 = +57; end
		46631: begin l_1 = -7;
				 l_2 = -57; end
		8396: begin l_1 = +7;
				 l_2 = +58; end
		42593: begin l_1 = +7;
				 l_2 = -58; end
		8268: begin l_1 = -7;
				 l_2 = +58; end
		42465: begin l_1 = -7;
				 l_2 = -58; end
		16728: begin l_1 = +7;
				 l_2 = +59; end
		34261: begin l_1 = +7;
				 l_2 = -59; end
		16600: begin l_1 = -7;
				 l_2 = +59; end
		34133: begin l_1 = -7;
				 l_2 = -59; end
		33392: begin l_1 = +7;
				 l_2 = +60; end
		17597: begin l_1 = +7;
				 l_2 = -60; end
		33264: begin l_1 = -7;
				 l_2 = +60; end
		17469: begin l_1 = -7;
				 l_2 = -60; end
		15859: begin l_1 = +7;
				 l_2 = +61; end
		35130: begin l_1 = +7;
				 l_2 = -61; end
		15731: begin l_1 = -7;
				 l_2 = +61; end
		35002: begin l_1 = -7;
				 l_2 = -61; end
		31654: begin l_1 = +7;
				 l_2 = +62; end
		19335: begin l_1 = +7;
				 l_2 = -62; end
		31526: begin l_1 = -7;
				 l_2 = +62; end
		19207: begin l_1 = -7;
				 l_2 = -62; end
		12383: begin l_1 = +7;
				 l_2 = +63; end
		38606: begin l_1 = +7;
				 l_2 = -63; end
		12255: begin l_1 = -7;
				 l_2 = +63; end
		38478: begin l_1 = -7;
				 l_2 = -63; end
		24702: begin l_1 = +7;
				 l_2 = +64; end
		26287: begin l_1 = +7;
				 l_2 = -64; end
		24574: begin l_1 = -7;
				 l_2 = +64; end
		26159: begin l_1 = -7;
				 l_2 = -64; end
		49340: begin l_1 = +7;
				 l_2 = +65; end
		1649: begin l_1 = +7;
				 l_2 = -65; end
		49212: begin l_1 = -7;
				 l_2 = +65; end
		1521: begin l_1 = -7;
				 l_2 = -65; end
		47755: begin l_1 = +7;
				 l_2 = +66; end
		3234: begin l_1 = +7;
				 l_2 = -66; end
		47627: begin l_1 = -7;
				 l_2 = +66; end
		3106: begin l_1 = -7;
				 l_2 = -66; end
		44585: begin l_1 = +7;
				 l_2 = +67; end
		6404: begin l_1 = +7;
				 l_2 = -67; end
		44457: begin l_1 = -7;
				 l_2 = +67; end
		6276: begin l_1 = -7;
				 l_2 = -67; end
		38245: begin l_1 = +7;
				 l_2 = +68; end
		12744: begin l_1 = +7;
				 l_2 = -68; end
		38117: begin l_1 = -7;
				 l_2 = +68; end
		12616: begin l_1 = -7;
				 l_2 = -68; end
		384: begin l_1 = -8;
				 l_2 = +10; end
		50477: begin l_1 = -8;
				 l_2 = -9; end
		640: begin l_1 = +8;
				 l_2 = +10; end
		50221: begin l_1 = -8;
				 l_2 = -10; end
		1152: begin l_1 = +8;
				 l_2 = +11; end
		49965: begin l_1 = +8;
				 l_2 = -11; end
		896: begin l_1 = -8;
				 l_2 = +11; end
		49709: begin l_1 = -8;
				 l_2 = -11; end
		2176: begin l_1 = +8;
				 l_2 = +12; end
		48941: begin l_1 = +8;
				 l_2 = -12; end
		1920: begin l_1 = -8;
				 l_2 = +12; end
		48685: begin l_1 = -8;
				 l_2 = -12; end
		4224: begin l_1 = +8;
				 l_2 = +13; end
		46893: begin l_1 = +8;
				 l_2 = -13; end
		3968: begin l_1 = -8;
				 l_2 = +13; end
		46637: begin l_1 = -8;
				 l_2 = -13; end
		8320: begin l_1 = +8;
				 l_2 = +14; end
		42797: begin l_1 = +8;
				 l_2 = -14; end
		8064: begin l_1 = -8;
				 l_2 = +14; end
		42541: begin l_1 = -8;
				 l_2 = -14; end
		16512: begin l_1 = +8;
				 l_2 = +15; end
		34605: begin l_1 = +8;
				 l_2 = -15; end
		16256: begin l_1 = -8;
				 l_2 = +15; end
		34349: begin l_1 = -8;
				 l_2 = -15; end
		32896: begin l_1 = +8;
				 l_2 = +16; end
		18221: begin l_1 = +8;
				 l_2 = -16; end
		32640: begin l_1 = -8;
				 l_2 = +16; end
		17965: begin l_1 = -8;
				 l_2 = -16; end
		14803: begin l_1 = +8;
				 l_2 = +17; end
		36314: begin l_1 = +8;
				 l_2 = -17; end
		14547: begin l_1 = -8;
				 l_2 = +17; end
		36058: begin l_1 = -8;
				 l_2 = -17; end
		29478: begin l_1 = +8;
				 l_2 = +18; end
		21639: begin l_1 = +8;
				 l_2 = -18; end
		29222: begin l_1 = -8;
				 l_2 = +18; end
		21383: begin l_1 = -8;
				 l_2 = -18; end
		7967: begin l_1 = +8;
				 l_2 = +19; end
		43150: begin l_1 = +8;
				 l_2 = -19; end
		7711: begin l_1 = -8;
				 l_2 = +19; end
		42894: begin l_1 = -8;
				 l_2 = -19; end
		15806: begin l_1 = +8;
				 l_2 = +20; end
		35311: begin l_1 = +8;
				 l_2 = -20; end
		15550: begin l_1 = -8;
				 l_2 = +20; end
		35055: begin l_1 = -8;
				 l_2 = -20; end
		31484: begin l_1 = +8;
				 l_2 = +21; end
		19633: begin l_1 = +8;
				 l_2 = -21; end
		31228: begin l_1 = -8;
				 l_2 = +21; end
		19377: begin l_1 = -8;
				 l_2 = -21; end
		11979: begin l_1 = +8;
				 l_2 = +22; end
		39138: begin l_1 = +8;
				 l_2 = -22; end
		11723: begin l_1 = -8;
				 l_2 = +22; end
		38882: begin l_1 = -8;
				 l_2 = -22; end
		23830: begin l_1 = +8;
				 l_2 = +23; end
		27287: begin l_1 = +8;
				 l_2 = -23; end
		23574: begin l_1 = -8;
				 l_2 = +23; end
		27031: begin l_1 = -8;
				 l_2 = -23; end
		47532: begin l_1 = +8;
				 l_2 = +24; end
		3585: begin l_1 = +8;
				 l_2 = -24; end
		47276: begin l_1 = -8;
				 l_2 = +24; end
		3329: begin l_1 = -8;
				 l_2 = -24; end
		44075: begin l_1 = +8;
				 l_2 = +25; end
		7042: begin l_1 = +8;
				 l_2 = -25; end
		43819: begin l_1 = -8;
				 l_2 = +25; end
		6786: begin l_1 = -8;
				 l_2 = -25; end
		37161: begin l_1 = +8;
				 l_2 = +26; end
		13956: begin l_1 = +8;
				 l_2 = -26; end
		36905: begin l_1 = -8;
				 l_2 = +26; end
		13700: begin l_1 = -8;
				 l_2 = -26; end
		23333: begin l_1 = +8;
				 l_2 = +27; end
		27784: begin l_1 = +8;
				 l_2 = -27; end
		23077: begin l_1 = -8;
				 l_2 = +27; end
		27528: begin l_1 = -8;
				 l_2 = -27; end
		46538: begin l_1 = +8;
				 l_2 = +28; end
		4579: begin l_1 = +8;
				 l_2 = -28; end
		46282: begin l_1 = -8;
				 l_2 = +28; end
		4323: begin l_1 = -8;
				 l_2 = -28; end
		42087: begin l_1 = +8;
				 l_2 = +29; end
		9030: begin l_1 = +8;
				 l_2 = -29; end
		41831: begin l_1 = -8;
				 l_2 = +29; end
		8774: begin l_1 = -8;
				 l_2 = -29; end
		33185: begin l_1 = +8;
				 l_2 = +30; end
		17932: begin l_1 = +8;
				 l_2 = -30; end
		32929: begin l_1 = -8;
				 l_2 = +30; end
		17676: begin l_1 = -8;
				 l_2 = -30; end
		15381: begin l_1 = +8;
				 l_2 = +31; end
		35736: begin l_1 = +8;
				 l_2 = -31; end
		15125: begin l_1 = -8;
				 l_2 = +31; end
		35480: begin l_1 = -8;
				 l_2 = -31; end
		30634: begin l_1 = +8;
				 l_2 = +32; end
		20483: begin l_1 = +8;
				 l_2 = -32; end
		30378: begin l_1 = -8;
				 l_2 = +32; end
		20227: begin l_1 = -8;
				 l_2 = -32; end
		10279: begin l_1 = +8;
				 l_2 = +33; end
		40838: begin l_1 = +8;
				 l_2 = -33; end
		10023: begin l_1 = -8;
				 l_2 = +33; end
		40582: begin l_1 = -8;
				 l_2 = -33; end
		20430: begin l_1 = +8;
				 l_2 = +34; end
		30687: begin l_1 = +8;
				 l_2 = -34; end
		20174: begin l_1 = -8;
				 l_2 = +34; end
		30431: begin l_1 = -8;
				 l_2 = -34; end
		40732: begin l_1 = +8;
				 l_2 = +35; end
		10385: begin l_1 = +8;
				 l_2 = -35; end
		40476: begin l_1 = -8;
				 l_2 = +35; end
		10129: begin l_1 = -8;
				 l_2 = -35; end
		30475: begin l_1 = +8;
				 l_2 = +36; end
		20642: begin l_1 = +8;
				 l_2 = -36; end
		30219: begin l_1 = -8;
				 l_2 = +36; end
		20386: begin l_1 = -8;
				 l_2 = -36; end
		9961: begin l_1 = +8;
				 l_2 = +37; end
		41156: begin l_1 = +8;
				 l_2 = -37; end
		9705: begin l_1 = -8;
				 l_2 = +37; end
		40900: begin l_1 = -8;
				 l_2 = -37; end
		19794: begin l_1 = +8;
				 l_2 = +38; end
		31323: begin l_1 = +8;
				 l_2 = -38; end
		19538: begin l_1 = -8;
				 l_2 = +38; end
		31067: begin l_1 = -8;
				 l_2 = -38; end
		39460: begin l_1 = +8;
				 l_2 = +39; end
		11657: begin l_1 = +8;
				 l_2 = -39; end
		39204: begin l_1 = -8;
				 l_2 = +39; end
		11401: begin l_1 = -8;
				 l_2 = -39; end
		27931: begin l_1 = +8;
				 l_2 = +40; end
		23186: begin l_1 = +8;
				 l_2 = -40; end
		27675: begin l_1 = -8;
				 l_2 = +40; end
		22930: begin l_1 = -8;
				 l_2 = -40; end
		4873: begin l_1 = +8;
				 l_2 = +41; end
		46244: begin l_1 = +8;
				 l_2 = -41; end
		4617: begin l_1 = -8;
				 l_2 = +41; end
		45988: begin l_1 = -8;
				 l_2 = -41; end
		9618: begin l_1 = +8;
				 l_2 = +42; end
		41499: begin l_1 = +8;
				 l_2 = -42; end
		9362: begin l_1 = -8;
				 l_2 = +42; end
		41243: begin l_1 = -8;
				 l_2 = -42; end
		19108: begin l_1 = +8;
				 l_2 = +43; end
		32009: begin l_1 = +8;
				 l_2 = -43; end
		18852: begin l_1 = -8;
				 l_2 = +43; end
		31753: begin l_1 = -8;
				 l_2 = -43; end
		38088: begin l_1 = +8;
				 l_2 = +44; end
		13029: begin l_1 = +8;
				 l_2 = -44; end
		37832: begin l_1 = -8;
				 l_2 = +44; end
		12773: begin l_1 = -8;
				 l_2 = -44; end
		25187: begin l_1 = +8;
				 l_2 = +45; end
		25930: begin l_1 = +8;
				 l_2 = -45; end
		24931: begin l_1 = -8;
				 l_2 = +45; end
		25674: begin l_1 = -8;
				 l_2 = -45; end
		50246: begin l_1 = +8;
				 l_2 = +46; end
		871: begin l_1 = +8;
				 l_2 = -46; end
		49990: begin l_1 = -8;
				 l_2 = +46; end
		615: begin l_1 = -8;
				 l_2 = -46; end
		49503: begin l_1 = +8;
				 l_2 = +47; end
		1614: begin l_1 = +8;
				 l_2 = -47; end
		49247: begin l_1 = -8;
				 l_2 = +47; end
		1358: begin l_1 = -8;
				 l_2 = -47; end
		48017: begin l_1 = +8;
				 l_2 = +48; end
		3100: begin l_1 = +8;
				 l_2 = -48; end
		47761: begin l_1 = -8;
				 l_2 = +48; end
		2844: begin l_1 = -8;
				 l_2 = -48; end
		45045: begin l_1 = +8;
				 l_2 = +49; end
		6072: begin l_1 = +8;
				 l_2 = -49; end
		44789: begin l_1 = -8;
				 l_2 = +49; end
		5816: begin l_1 = -8;
				 l_2 = -49; end
		39101: begin l_1 = +8;
				 l_2 = +50; end
		12016: begin l_1 = +8;
				 l_2 = -50; end
		38845: begin l_1 = -8;
				 l_2 = +50; end
		11760: begin l_1 = -8;
				 l_2 = -50; end
		27213: begin l_1 = +8;
				 l_2 = +51; end
		23904: begin l_1 = +8;
				 l_2 = -51; end
		26957: begin l_1 = -8;
				 l_2 = +51; end
		23648: begin l_1 = -8;
				 l_2 = -51; end
		3437: begin l_1 = +8;
				 l_2 = +52; end
		47680: begin l_1 = +8;
				 l_2 = -52; end
		3181: begin l_1 = -8;
				 l_2 = +52; end
		47424: begin l_1 = -8;
				 l_2 = -52; end
		6746: begin l_1 = +8;
				 l_2 = +53; end
		44371: begin l_1 = +8;
				 l_2 = -53; end
		6490: begin l_1 = -8;
				 l_2 = +53; end
		44115: begin l_1 = -8;
				 l_2 = -53; end
		13364: begin l_1 = +8;
				 l_2 = +54; end
		37753: begin l_1 = +8;
				 l_2 = -54; end
		13108: begin l_1 = -8;
				 l_2 = +54; end
		37497: begin l_1 = -8;
				 l_2 = -54; end
		26600: begin l_1 = +8;
				 l_2 = +55; end
		24517: begin l_1 = +8;
				 l_2 = -55; end
		26344: begin l_1 = -8;
				 l_2 = +55; end
		24261: begin l_1 = -8;
				 l_2 = -55; end
		2211: begin l_1 = +8;
				 l_2 = +56; end
		48906: begin l_1 = +8;
				 l_2 = -56; end
		1955: begin l_1 = -8;
				 l_2 = +56; end
		48650: begin l_1 = -8;
				 l_2 = -56; end
		4294: begin l_1 = +8;
				 l_2 = +57; end
		46823: begin l_1 = +8;
				 l_2 = -57; end
		4038: begin l_1 = -8;
				 l_2 = +57; end
		46567: begin l_1 = -8;
				 l_2 = -57; end
		8460: begin l_1 = +8;
				 l_2 = +58; end
		42657: begin l_1 = +8;
				 l_2 = -58; end
		8204: begin l_1 = -8;
				 l_2 = +58; end
		42401: begin l_1 = -8;
				 l_2 = -58; end
		16792: begin l_1 = +8;
				 l_2 = +59; end
		34325: begin l_1 = +8;
				 l_2 = -59; end
		16536: begin l_1 = -8;
				 l_2 = +59; end
		34069: begin l_1 = -8;
				 l_2 = -59; end
		33456: begin l_1 = +8;
				 l_2 = +60; end
		17661: begin l_1 = +8;
				 l_2 = -60; end
		33200: begin l_1 = -8;
				 l_2 = +60; end
		17405: begin l_1 = -8;
				 l_2 = -60; end
		15923: begin l_1 = +8;
				 l_2 = +61; end
		35194: begin l_1 = +8;
				 l_2 = -61; end
		15667: begin l_1 = -8;
				 l_2 = +61; end
		34938: begin l_1 = -8;
				 l_2 = -61; end
		31718: begin l_1 = +8;
				 l_2 = +62; end
		19399: begin l_1 = +8;
				 l_2 = -62; end
		31462: begin l_1 = -8;
				 l_2 = +62; end
		19143: begin l_1 = -8;
				 l_2 = -62; end
		12447: begin l_1 = +8;
				 l_2 = +63; end
		38670: begin l_1 = +8;
				 l_2 = -63; end
		12191: begin l_1 = -8;
				 l_2 = +63; end
		38414: begin l_1 = -8;
				 l_2 = -63; end
		24766: begin l_1 = +8;
				 l_2 = +64; end
		26351: begin l_1 = +8;
				 l_2 = -64; end
		24510: begin l_1 = -8;
				 l_2 = +64; end
		26095: begin l_1 = -8;
				 l_2 = -64; end
		49404: begin l_1 = +8;
				 l_2 = +65; end
		1713: begin l_1 = +8;
				 l_2 = -65; end
		49148: begin l_1 = -8;
				 l_2 = +65; end
		1457: begin l_1 = -8;
				 l_2 = -65; end
		47819: begin l_1 = +8;
				 l_2 = +66; end
		3298: begin l_1 = +8;
				 l_2 = -66; end
		47563: begin l_1 = -8;
				 l_2 = +66; end
		3042: begin l_1 = -8;
				 l_2 = -66; end
		44649: begin l_1 = +8;
				 l_2 = +67; end
		6468: begin l_1 = +8;
				 l_2 = -67; end
		44393: begin l_1 = -8;
				 l_2 = +67; end
		6212: begin l_1 = -8;
				 l_2 = -67; end
		38309: begin l_1 = +8;
				 l_2 = +68; end
		12808: begin l_1 = +8;
				 l_2 = -68; end
		38053: begin l_1 = -8;
				 l_2 = +68; end
		12552: begin l_1 = -8;
				 l_2 = -68; end
		768: begin l_1 = -9;
				 l_2 = +11; end
		50093: begin l_1 = -9;
				 l_2 = -10; end
		1280: begin l_1 = +9;
				 l_2 = +11; end
		49581: begin l_1 = -9;
				 l_2 = -11; end
		2304: begin l_1 = +9;
				 l_2 = +12; end
		49069: begin l_1 = +9;
				 l_2 = -12; end
		1792: begin l_1 = -9;
				 l_2 = +12; end
		48557: begin l_1 = -9;
				 l_2 = -12; end
		4352: begin l_1 = +9;
				 l_2 = +13; end
		47021: begin l_1 = +9;
				 l_2 = -13; end
		3840: begin l_1 = -9;
				 l_2 = +13; end
		46509: begin l_1 = -9;
				 l_2 = -13; end
		8448: begin l_1 = +9;
				 l_2 = +14; end
		42925: begin l_1 = +9;
				 l_2 = -14; end
		7936: begin l_1 = -9;
				 l_2 = +14; end
		42413: begin l_1 = -9;
				 l_2 = -14; end
		16640: begin l_1 = +9;
				 l_2 = +15; end
		34733: begin l_1 = +9;
				 l_2 = -15; end
		16128: begin l_1 = -9;
				 l_2 = +15; end
		34221: begin l_1 = -9;
				 l_2 = -15; end
		33024: begin l_1 = +9;
				 l_2 = +16; end
		18349: begin l_1 = +9;
				 l_2 = -16; end
		32512: begin l_1 = -9;
				 l_2 = +16; end
		17837: begin l_1 = -9;
				 l_2 = -16; end
		14931: begin l_1 = +9;
				 l_2 = +17; end
		36442: begin l_1 = +9;
				 l_2 = -17; end
		14419: begin l_1 = -9;
				 l_2 = +17; end
		35930: begin l_1 = -9;
				 l_2 = -17; end
		29606: begin l_1 = +9;
				 l_2 = +18; end
		21767: begin l_1 = +9;
				 l_2 = -18; end
		29094: begin l_1 = -9;
				 l_2 = +18; end
		21255: begin l_1 = -9;
				 l_2 = -18; end
		8095: begin l_1 = +9;
				 l_2 = +19; end
		43278: begin l_1 = +9;
				 l_2 = -19; end
		7583: begin l_1 = -9;
				 l_2 = +19; end
		42766: begin l_1 = -9;
				 l_2 = -19; end
		15934: begin l_1 = +9;
				 l_2 = +20; end
		35439: begin l_1 = +9;
				 l_2 = -20; end
		15422: begin l_1 = -9;
				 l_2 = +20; end
		34927: begin l_1 = -9;
				 l_2 = -20; end
		31612: begin l_1 = +9;
				 l_2 = +21; end
		19761: begin l_1 = +9;
				 l_2 = -21; end
		31100: begin l_1 = -9;
				 l_2 = +21; end
		19249: begin l_1 = -9;
				 l_2 = -21; end
		12107: begin l_1 = +9;
				 l_2 = +22; end
		39266: begin l_1 = +9;
				 l_2 = -22; end
		11595: begin l_1 = -9;
				 l_2 = +22; end
		38754: begin l_1 = -9;
				 l_2 = -22; end
		23958: begin l_1 = +9;
				 l_2 = +23; end
		27415: begin l_1 = +9;
				 l_2 = -23; end
		23446: begin l_1 = -9;
				 l_2 = +23; end
		26903: begin l_1 = -9;
				 l_2 = -23; end
		47660: begin l_1 = +9;
				 l_2 = +24; end
		3713: begin l_1 = +9;
				 l_2 = -24; end
		47148: begin l_1 = -9;
				 l_2 = +24; end
		3201: begin l_1 = -9;
				 l_2 = -24; end
		44203: begin l_1 = +9;
				 l_2 = +25; end
		7170: begin l_1 = +9;
				 l_2 = -25; end
		43691: begin l_1 = -9;
				 l_2 = +25; end
		6658: begin l_1 = -9;
				 l_2 = -25; end
		37289: begin l_1 = +9;
				 l_2 = +26; end
		14084: begin l_1 = +9;
				 l_2 = -26; end
		36777: begin l_1 = -9;
				 l_2 = +26; end
		13572: begin l_1 = -9;
				 l_2 = -26; end
		23461: begin l_1 = +9;
				 l_2 = +27; end
		27912: begin l_1 = +9;
				 l_2 = -27; end
		22949: begin l_1 = -9;
				 l_2 = +27; end
		27400: begin l_1 = -9;
				 l_2 = -27; end
		46666: begin l_1 = +9;
				 l_2 = +28; end
		4707: begin l_1 = +9;
				 l_2 = -28; end
		46154: begin l_1 = -9;
				 l_2 = +28; end
		4195: begin l_1 = -9;
				 l_2 = -28; end
		42215: begin l_1 = +9;
				 l_2 = +29; end
		9158: begin l_1 = +9;
				 l_2 = -29; end
		41703: begin l_1 = -9;
				 l_2 = +29; end
		8646: begin l_1 = -9;
				 l_2 = -29; end
		33313: begin l_1 = +9;
				 l_2 = +30; end
		18060: begin l_1 = +9;
				 l_2 = -30; end
		32801: begin l_1 = -9;
				 l_2 = +30; end
		17548: begin l_1 = -9;
				 l_2 = -30; end
		15509: begin l_1 = +9;
				 l_2 = +31; end
		35864: begin l_1 = +9;
				 l_2 = -31; end
		14997: begin l_1 = -9;
				 l_2 = +31; end
		35352: begin l_1 = -9;
				 l_2 = -31; end
		30762: begin l_1 = +9;
				 l_2 = +32; end
		20611: begin l_1 = +9;
				 l_2 = -32; end
		30250: begin l_1 = -9;
				 l_2 = +32; end
		20099: begin l_1 = -9;
				 l_2 = -32; end
		10407: begin l_1 = +9;
				 l_2 = +33; end
		40966: begin l_1 = +9;
				 l_2 = -33; end
		9895: begin l_1 = -9;
				 l_2 = +33; end
		40454: begin l_1 = -9;
				 l_2 = -33; end
		20558: begin l_1 = +9;
				 l_2 = +34; end
		30815: begin l_1 = +9;
				 l_2 = -34; end
		20046: begin l_1 = -9;
				 l_2 = +34; end
		30303: begin l_1 = -9;
				 l_2 = -34; end
		40860: begin l_1 = +9;
				 l_2 = +35; end
		10513: begin l_1 = +9;
				 l_2 = -35; end
		40348: begin l_1 = -9;
				 l_2 = +35; end
		10001: begin l_1 = -9;
				 l_2 = -35; end
		30603: begin l_1 = +9;
				 l_2 = +36; end
		20770: begin l_1 = +9;
				 l_2 = -36; end
		30091: begin l_1 = -9;
				 l_2 = +36; end
		20258: begin l_1 = -9;
				 l_2 = -36; end
		10089: begin l_1 = +9;
				 l_2 = +37; end
		41284: begin l_1 = +9;
				 l_2 = -37; end
		9577: begin l_1 = -9;
				 l_2 = +37; end
		40772: begin l_1 = -9;
				 l_2 = -37; end
		19922: begin l_1 = +9;
				 l_2 = +38; end
		31451: begin l_1 = +9;
				 l_2 = -38; end
		19410: begin l_1 = -9;
				 l_2 = +38; end
		30939: begin l_1 = -9;
				 l_2 = -38; end
		39588: begin l_1 = +9;
				 l_2 = +39; end
		11785: begin l_1 = +9;
				 l_2 = -39; end
		39076: begin l_1 = -9;
				 l_2 = +39; end
		11273: begin l_1 = -9;
				 l_2 = -39; end
		28059: begin l_1 = +9;
				 l_2 = +40; end
		23314: begin l_1 = +9;
				 l_2 = -40; end
		27547: begin l_1 = -9;
				 l_2 = +40; end
		22802: begin l_1 = -9;
				 l_2 = -40; end
		5001: begin l_1 = +9;
				 l_2 = +41; end
		46372: begin l_1 = +9;
				 l_2 = -41; end
		4489: begin l_1 = -9;
				 l_2 = +41; end
		45860: begin l_1 = -9;
				 l_2 = -41; end
		9746: begin l_1 = +9;
				 l_2 = +42; end
		41627: begin l_1 = +9;
				 l_2 = -42; end
		9234: begin l_1 = -9;
				 l_2 = +42; end
		41115: begin l_1 = -9;
				 l_2 = -42; end
		19236: begin l_1 = +9;
				 l_2 = +43; end
		32137: begin l_1 = +9;
				 l_2 = -43; end
		18724: begin l_1 = -9;
				 l_2 = +43; end
		31625: begin l_1 = -9;
				 l_2 = -43; end
		38216: begin l_1 = +9;
				 l_2 = +44; end
		13157: begin l_1 = +9;
				 l_2 = -44; end
		37704: begin l_1 = -9;
				 l_2 = +44; end
		12645: begin l_1 = -9;
				 l_2 = -44; end
		25315: begin l_1 = +9;
				 l_2 = +45; end
		26058: begin l_1 = +9;
				 l_2 = -45; end
		24803: begin l_1 = -9;
				 l_2 = +45; end
		25546: begin l_1 = -9;
				 l_2 = -45; end
		50374: begin l_1 = +9;
				 l_2 = +46; end
		999: begin l_1 = +9;
				 l_2 = -46; end
		49862: begin l_1 = -9;
				 l_2 = +46; end
		487: begin l_1 = -9;
				 l_2 = -46; end
		49631: begin l_1 = +9;
				 l_2 = +47; end
		1742: begin l_1 = +9;
				 l_2 = -47; end
		49119: begin l_1 = -9;
				 l_2 = +47; end
		1230: begin l_1 = -9;
				 l_2 = -47; end
		48145: begin l_1 = +9;
				 l_2 = +48; end
		3228: begin l_1 = +9;
				 l_2 = -48; end
		47633: begin l_1 = -9;
				 l_2 = +48; end
		2716: begin l_1 = -9;
				 l_2 = -48; end
		45173: begin l_1 = +9;
				 l_2 = +49; end
		6200: begin l_1 = +9;
				 l_2 = -49; end
		44661: begin l_1 = -9;
				 l_2 = +49; end
		5688: begin l_1 = -9;
				 l_2 = -49; end
		39229: begin l_1 = +9;
				 l_2 = +50; end
		12144: begin l_1 = +9;
				 l_2 = -50; end
		38717: begin l_1 = -9;
				 l_2 = +50; end
		11632: begin l_1 = -9;
				 l_2 = -50; end
		27341: begin l_1 = +9;
				 l_2 = +51; end
		24032: begin l_1 = +9;
				 l_2 = -51; end
		26829: begin l_1 = -9;
				 l_2 = +51; end
		23520: begin l_1 = -9;
				 l_2 = -51; end
		3565: begin l_1 = +9;
				 l_2 = +52; end
		47808: begin l_1 = +9;
				 l_2 = -52; end
		3053: begin l_1 = -9;
				 l_2 = +52; end
		47296: begin l_1 = -9;
				 l_2 = -52; end
		6874: begin l_1 = +9;
				 l_2 = +53; end
		44499: begin l_1 = +9;
				 l_2 = -53; end
		6362: begin l_1 = -9;
				 l_2 = +53; end
		43987: begin l_1 = -9;
				 l_2 = -53; end
		13492: begin l_1 = +9;
				 l_2 = +54; end
		37881: begin l_1 = +9;
				 l_2 = -54; end
		12980: begin l_1 = -9;
				 l_2 = +54; end
		37369: begin l_1 = -9;
				 l_2 = -54; end
		26728: begin l_1 = +9;
				 l_2 = +55; end
		24645: begin l_1 = +9;
				 l_2 = -55; end
		26216: begin l_1 = -9;
				 l_2 = +55; end
		24133: begin l_1 = -9;
				 l_2 = -55; end
		2339: begin l_1 = +9;
				 l_2 = +56; end
		49034: begin l_1 = +9;
				 l_2 = -56; end
		1827: begin l_1 = -9;
				 l_2 = +56; end
		48522: begin l_1 = -9;
				 l_2 = -56; end
		4422: begin l_1 = +9;
				 l_2 = +57; end
		46951: begin l_1 = +9;
				 l_2 = -57; end
		3910: begin l_1 = -9;
				 l_2 = +57; end
		46439: begin l_1 = -9;
				 l_2 = -57; end
		8588: begin l_1 = +9;
				 l_2 = +58; end
		42785: begin l_1 = +9;
				 l_2 = -58; end
		8076: begin l_1 = -9;
				 l_2 = +58; end
		42273: begin l_1 = -9;
				 l_2 = -58; end
		16920: begin l_1 = +9;
				 l_2 = +59; end
		34453: begin l_1 = +9;
				 l_2 = -59; end
		16408: begin l_1 = -9;
				 l_2 = +59; end
		33941: begin l_1 = -9;
				 l_2 = -59; end
		33584: begin l_1 = +9;
				 l_2 = +60; end
		17789: begin l_1 = +9;
				 l_2 = -60; end
		33072: begin l_1 = -9;
				 l_2 = +60; end
		17277: begin l_1 = -9;
				 l_2 = -60; end
		16051: begin l_1 = +9;
				 l_2 = +61; end
		35322: begin l_1 = +9;
				 l_2 = -61; end
		15539: begin l_1 = -9;
				 l_2 = +61; end
		34810: begin l_1 = -9;
				 l_2 = -61; end
		31846: begin l_1 = +9;
				 l_2 = +62; end
		19527: begin l_1 = +9;
				 l_2 = -62; end
		31334: begin l_1 = -9;
				 l_2 = +62; end
		19015: begin l_1 = -9;
				 l_2 = -62; end
		12575: begin l_1 = +9;
				 l_2 = +63; end
		38798: begin l_1 = +9;
				 l_2 = -63; end
		12063: begin l_1 = -9;
				 l_2 = +63; end
		38286: begin l_1 = -9;
				 l_2 = -63; end
		24894: begin l_1 = +9;
				 l_2 = +64; end
		26479: begin l_1 = +9;
				 l_2 = -64; end
		24382: begin l_1 = -9;
				 l_2 = +64; end
		25967: begin l_1 = -9;
				 l_2 = -64; end
		49532: begin l_1 = +9;
				 l_2 = +65; end
		1841: begin l_1 = +9;
				 l_2 = -65; end
		49020: begin l_1 = -9;
				 l_2 = +65; end
		1329: begin l_1 = -9;
				 l_2 = -65; end
		47947: begin l_1 = +9;
				 l_2 = +66; end
		3426: begin l_1 = +9;
				 l_2 = -66; end
		47435: begin l_1 = -9;
				 l_2 = +66; end
		2914: begin l_1 = -9;
				 l_2 = -66; end
		44777: begin l_1 = +9;
				 l_2 = +67; end
		6596: begin l_1 = +9;
				 l_2 = -67; end
		44265: begin l_1 = -9;
				 l_2 = +67; end
		6084: begin l_1 = -9;
				 l_2 = -67; end
		38437: begin l_1 = +9;
				 l_2 = +68; end
		12936: begin l_1 = +9;
				 l_2 = -68; end
		37925: begin l_1 = -9;
				 l_2 = +68; end
		12424: begin l_1 = -9;
				 l_2 = -68; end
		1536: begin l_1 = -10;
				 l_2 = +12; end
		49325: begin l_1 = -10;
				 l_2 = -11; end
		2560: begin l_1 = +10;
				 l_2 = +12; end
		48301: begin l_1 = -10;
				 l_2 = -12; end
		4608: begin l_1 = +10;
				 l_2 = +13; end
		47277: begin l_1 = +10;
				 l_2 = -13; end
		3584: begin l_1 = -10;
				 l_2 = +13; end
		46253: begin l_1 = -10;
				 l_2 = -13; end
		8704: begin l_1 = +10;
				 l_2 = +14; end
		43181: begin l_1 = +10;
				 l_2 = -14; end
		7680: begin l_1 = -10;
				 l_2 = +14; end
		42157: begin l_1 = -10;
				 l_2 = -14; end
		16896: begin l_1 = +10;
				 l_2 = +15; end
		34989: begin l_1 = +10;
				 l_2 = -15; end
		15872: begin l_1 = -10;
				 l_2 = +15; end
		33965: begin l_1 = -10;
				 l_2 = -15; end
		33280: begin l_1 = +10;
				 l_2 = +16; end
		18605: begin l_1 = +10;
				 l_2 = -16; end
		32256: begin l_1 = -10;
				 l_2 = +16; end
		17581: begin l_1 = -10;
				 l_2 = -16; end
		15187: begin l_1 = +10;
				 l_2 = +17; end
		36698: begin l_1 = +10;
				 l_2 = -17; end
		14163: begin l_1 = -10;
				 l_2 = +17; end
		35674: begin l_1 = -10;
				 l_2 = -17; end
		29862: begin l_1 = +10;
				 l_2 = +18; end
		22023: begin l_1 = +10;
				 l_2 = -18; end
		28838: begin l_1 = -10;
				 l_2 = +18; end
		20999: begin l_1 = -10;
				 l_2 = -18; end
		8351: begin l_1 = +10;
				 l_2 = +19; end
		43534: begin l_1 = +10;
				 l_2 = -19; end
		7327: begin l_1 = -10;
				 l_2 = +19; end
		42510: begin l_1 = -10;
				 l_2 = -19; end
		16190: begin l_1 = +10;
				 l_2 = +20; end
		35695: begin l_1 = +10;
				 l_2 = -20; end
		15166: begin l_1 = -10;
				 l_2 = +20; end
		34671: begin l_1 = -10;
				 l_2 = -20; end
		31868: begin l_1 = +10;
				 l_2 = +21; end
		20017: begin l_1 = +10;
				 l_2 = -21; end
		30844: begin l_1 = -10;
				 l_2 = +21; end
		18993: begin l_1 = -10;
				 l_2 = -21; end
		12363: begin l_1 = +10;
				 l_2 = +22; end
		39522: begin l_1 = +10;
				 l_2 = -22; end
		11339: begin l_1 = -10;
				 l_2 = +22; end
		38498: begin l_1 = -10;
				 l_2 = -22; end
		24214: begin l_1 = +10;
				 l_2 = +23; end
		27671: begin l_1 = +10;
				 l_2 = -23; end
		23190: begin l_1 = -10;
				 l_2 = +23; end
		26647: begin l_1 = -10;
				 l_2 = -23; end
		47916: begin l_1 = +10;
				 l_2 = +24; end
		3969: begin l_1 = +10;
				 l_2 = -24; end
		46892: begin l_1 = -10;
				 l_2 = +24; end
		2945: begin l_1 = -10;
				 l_2 = -24; end
		44459: begin l_1 = +10;
				 l_2 = +25; end
		7426: begin l_1 = +10;
				 l_2 = -25; end
		43435: begin l_1 = -10;
				 l_2 = +25; end
		6402: begin l_1 = -10;
				 l_2 = -25; end
		37545: begin l_1 = +10;
				 l_2 = +26; end
		14340: begin l_1 = +10;
				 l_2 = -26; end
		36521: begin l_1 = -10;
				 l_2 = +26; end
		13316: begin l_1 = -10;
				 l_2 = -26; end
		23717: begin l_1 = +10;
				 l_2 = +27; end
		28168: begin l_1 = +10;
				 l_2 = -27; end
		22693: begin l_1 = -10;
				 l_2 = +27; end
		27144: begin l_1 = -10;
				 l_2 = -27; end
		46922: begin l_1 = +10;
				 l_2 = +28; end
		4963: begin l_1 = +10;
				 l_2 = -28; end
		45898: begin l_1 = -10;
				 l_2 = +28; end
		3939: begin l_1 = -10;
				 l_2 = -28; end
		42471: begin l_1 = +10;
				 l_2 = +29; end
		9414: begin l_1 = +10;
				 l_2 = -29; end
		41447: begin l_1 = -10;
				 l_2 = +29; end
		8390: begin l_1 = -10;
				 l_2 = -29; end
		33569: begin l_1 = +10;
				 l_2 = +30; end
		18316: begin l_1 = +10;
				 l_2 = -30; end
		32545: begin l_1 = -10;
				 l_2 = +30; end
		17292: begin l_1 = -10;
				 l_2 = -30; end
		15765: begin l_1 = +10;
				 l_2 = +31; end
		36120: begin l_1 = +10;
				 l_2 = -31; end
		14741: begin l_1 = -10;
				 l_2 = +31; end
		35096: begin l_1 = -10;
				 l_2 = -31; end
		31018: begin l_1 = +10;
				 l_2 = +32; end
		20867: begin l_1 = +10;
				 l_2 = -32; end
		29994: begin l_1 = -10;
				 l_2 = +32; end
		19843: begin l_1 = -10;
				 l_2 = -32; end
		10663: begin l_1 = +10;
				 l_2 = +33; end
		41222: begin l_1 = +10;
				 l_2 = -33; end
		9639: begin l_1 = -10;
				 l_2 = +33; end
		40198: begin l_1 = -10;
				 l_2 = -33; end
		20814: begin l_1 = +10;
				 l_2 = +34; end
		31071: begin l_1 = +10;
				 l_2 = -34; end
		19790: begin l_1 = -10;
				 l_2 = +34; end
		30047: begin l_1 = -10;
				 l_2 = -34; end
		41116: begin l_1 = +10;
				 l_2 = +35; end
		10769: begin l_1 = +10;
				 l_2 = -35; end
		40092: begin l_1 = -10;
				 l_2 = +35; end
		9745: begin l_1 = -10;
				 l_2 = -35; end
		30859: begin l_1 = +10;
				 l_2 = +36; end
		21026: begin l_1 = +10;
				 l_2 = -36; end
		29835: begin l_1 = -10;
				 l_2 = +36; end
		20002: begin l_1 = -10;
				 l_2 = -36; end
		10345: begin l_1 = +10;
				 l_2 = +37; end
		41540: begin l_1 = +10;
				 l_2 = -37; end
		9321: begin l_1 = -10;
				 l_2 = +37; end
		40516: begin l_1 = -10;
				 l_2 = -37; end
		20178: begin l_1 = +10;
				 l_2 = +38; end
		31707: begin l_1 = +10;
				 l_2 = -38; end
		19154: begin l_1 = -10;
				 l_2 = +38; end
		30683: begin l_1 = -10;
				 l_2 = -38; end
		39844: begin l_1 = +10;
				 l_2 = +39; end
		12041: begin l_1 = +10;
				 l_2 = -39; end
		38820: begin l_1 = -10;
				 l_2 = +39; end
		11017: begin l_1 = -10;
				 l_2 = -39; end
		28315: begin l_1 = +10;
				 l_2 = +40; end
		23570: begin l_1 = +10;
				 l_2 = -40; end
		27291: begin l_1 = -10;
				 l_2 = +40; end
		22546: begin l_1 = -10;
				 l_2 = -40; end
		5257: begin l_1 = +10;
				 l_2 = +41; end
		46628: begin l_1 = +10;
				 l_2 = -41; end
		4233: begin l_1 = -10;
				 l_2 = +41; end
		45604: begin l_1 = -10;
				 l_2 = -41; end
		10002: begin l_1 = +10;
				 l_2 = +42; end
		41883: begin l_1 = +10;
				 l_2 = -42; end
		8978: begin l_1 = -10;
				 l_2 = +42; end
		40859: begin l_1 = -10;
				 l_2 = -42; end
		19492: begin l_1 = +10;
				 l_2 = +43; end
		32393: begin l_1 = +10;
				 l_2 = -43; end
		18468: begin l_1 = -10;
				 l_2 = +43; end
		31369: begin l_1 = -10;
				 l_2 = -43; end
		38472: begin l_1 = +10;
				 l_2 = +44; end
		13413: begin l_1 = +10;
				 l_2 = -44; end
		37448: begin l_1 = -10;
				 l_2 = +44; end
		12389: begin l_1 = -10;
				 l_2 = -44; end
		25571: begin l_1 = +10;
				 l_2 = +45; end
		26314: begin l_1 = +10;
				 l_2 = -45; end
		24547: begin l_1 = -10;
				 l_2 = +45; end
		25290: begin l_1 = -10;
				 l_2 = -45; end
		50630: begin l_1 = +10;
				 l_2 = +46; end
		1255: begin l_1 = +10;
				 l_2 = -46; end
		49606: begin l_1 = -10;
				 l_2 = +46; end
		231: begin l_1 = -10;
				 l_2 = -46; end
		49887: begin l_1 = +10;
				 l_2 = +47; end
		1998: begin l_1 = +10;
				 l_2 = -47; end
		48863: begin l_1 = -10;
				 l_2 = +47; end
		974: begin l_1 = -10;
				 l_2 = -47; end
		48401: begin l_1 = +10;
				 l_2 = +48; end
		3484: begin l_1 = +10;
				 l_2 = -48; end
		47377: begin l_1 = -10;
				 l_2 = +48; end
		2460: begin l_1 = -10;
				 l_2 = -48; end
		45429: begin l_1 = +10;
				 l_2 = +49; end
		6456: begin l_1 = +10;
				 l_2 = -49; end
		44405: begin l_1 = -10;
				 l_2 = +49; end
		5432: begin l_1 = -10;
				 l_2 = -49; end
		39485: begin l_1 = +10;
				 l_2 = +50; end
		12400: begin l_1 = +10;
				 l_2 = -50; end
		38461: begin l_1 = -10;
				 l_2 = +50; end
		11376: begin l_1 = -10;
				 l_2 = -50; end
		27597: begin l_1 = +10;
				 l_2 = +51; end
		24288: begin l_1 = +10;
				 l_2 = -51; end
		26573: begin l_1 = -10;
				 l_2 = +51; end
		23264: begin l_1 = -10;
				 l_2 = -51; end
		3821: begin l_1 = +10;
				 l_2 = +52; end
		48064: begin l_1 = +10;
				 l_2 = -52; end
		2797: begin l_1 = -10;
				 l_2 = +52; end
		47040: begin l_1 = -10;
				 l_2 = -52; end
		7130: begin l_1 = +10;
				 l_2 = +53; end
		44755: begin l_1 = +10;
				 l_2 = -53; end
		6106: begin l_1 = -10;
				 l_2 = +53; end
		43731: begin l_1 = -10;
				 l_2 = -53; end
		13748: begin l_1 = +10;
				 l_2 = +54; end
		38137: begin l_1 = +10;
				 l_2 = -54; end
		12724: begin l_1 = -10;
				 l_2 = +54; end
		37113: begin l_1 = -10;
				 l_2 = -54; end
		26984: begin l_1 = +10;
				 l_2 = +55; end
		24901: begin l_1 = +10;
				 l_2 = -55; end
		25960: begin l_1 = -10;
				 l_2 = +55; end
		23877: begin l_1 = -10;
				 l_2 = -55; end
		2595: begin l_1 = +10;
				 l_2 = +56; end
		49290: begin l_1 = +10;
				 l_2 = -56; end
		1571: begin l_1 = -10;
				 l_2 = +56; end
		48266: begin l_1 = -10;
				 l_2 = -56; end
		4678: begin l_1 = +10;
				 l_2 = +57; end
		47207: begin l_1 = +10;
				 l_2 = -57; end
		3654: begin l_1 = -10;
				 l_2 = +57; end
		46183: begin l_1 = -10;
				 l_2 = -57; end
		8844: begin l_1 = +10;
				 l_2 = +58; end
		43041: begin l_1 = +10;
				 l_2 = -58; end
		7820: begin l_1 = -10;
				 l_2 = +58; end
		42017: begin l_1 = -10;
				 l_2 = -58; end
		17176: begin l_1 = +10;
				 l_2 = +59; end
		34709: begin l_1 = +10;
				 l_2 = -59; end
		16152: begin l_1 = -10;
				 l_2 = +59; end
		33685: begin l_1 = -10;
				 l_2 = -59; end
		33840: begin l_1 = +10;
				 l_2 = +60; end
		18045: begin l_1 = +10;
				 l_2 = -60; end
		32816: begin l_1 = -10;
				 l_2 = +60; end
		17021: begin l_1 = -10;
				 l_2 = -60; end
		16307: begin l_1 = +10;
				 l_2 = +61; end
		35578: begin l_1 = +10;
				 l_2 = -61; end
		15283: begin l_1 = -10;
				 l_2 = +61; end
		34554: begin l_1 = -10;
				 l_2 = -61; end
		32102: begin l_1 = +10;
				 l_2 = +62; end
		19783: begin l_1 = +10;
				 l_2 = -62; end
		31078: begin l_1 = -10;
				 l_2 = +62; end
		18759: begin l_1 = -10;
				 l_2 = -62; end
		12831: begin l_1 = +10;
				 l_2 = +63; end
		39054: begin l_1 = +10;
				 l_2 = -63; end
		11807: begin l_1 = -10;
				 l_2 = +63; end
		38030: begin l_1 = -10;
				 l_2 = -63; end
		25150: begin l_1 = +10;
				 l_2 = +64; end
		26735: begin l_1 = +10;
				 l_2 = -64; end
		24126: begin l_1 = -10;
				 l_2 = +64; end
		25711: begin l_1 = -10;
				 l_2 = -64; end
		49788: begin l_1 = +10;
				 l_2 = +65; end
		2097: begin l_1 = +10;
				 l_2 = -65; end
		48764: begin l_1 = -10;
				 l_2 = +65; end
		1073: begin l_1 = -10;
				 l_2 = -65; end
		48203: begin l_1 = +10;
				 l_2 = +66; end
		3682: begin l_1 = +10;
				 l_2 = -66; end
		47179: begin l_1 = -10;
				 l_2 = +66; end
		2658: begin l_1 = -10;
				 l_2 = -66; end
		45033: begin l_1 = +10;
				 l_2 = +67; end
		6852: begin l_1 = +10;
				 l_2 = -67; end
		44009: begin l_1 = -10;
				 l_2 = +67; end
		5828: begin l_1 = -10;
				 l_2 = -67; end
		38693: begin l_1 = +10;
				 l_2 = +68; end
		13192: begin l_1 = +10;
				 l_2 = -68; end
		37669: begin l_1 = -10;
				 l_2 = +68; end
		12168: begin l_1 = -10;
				 l_2 = -68; end
		3072: begin l_1 = -11;
				 l_2 = +13; end
		47789: begin l_1 = -11;
				 l_2 = -12; end
		5120: begin l_1 = +11;
				 l_2 = +13; end
		45741: begin l_1 = -11;
				 l_2 = -13; end
		9216: begin l_1 = +11;
				 l_2 = +14; end
		43693: begin l_1 = +11;
				 l_2 = -14; end
		7168: begin l_1 = -11;
				 l_2 = +14; end
		41645: begin l_1 = -11;
				 l_2 = -14; end
		17408: begin l_1 = +11;
				 l_2 = +15; end
		35501: begin l_1 = +11;
				 l_2 = -15; end
		15360: begin l_1 = -11;
				 l_2 = +15; end
		33453: begin l_1 = -11;
				 l_2 = -15; end
		33792: begin l_1 = +11;
				 l_2 = +16; end
		19117: begin l_1 = +11;
				 l_2 = -16; end
		31744: begin l_1 = -11;
				 l_2 = +16; end
		17069: begin l_1 = -11;
				 l_2 = -16; end
		15699: begin l_1 = +11;
				 l_2 = +17; end
		37210: begin l_1 = +11;
				 l_2 = -17; end
		13651: begin l_1 = -11;
				 l_2 = +17; end
		35162: begin l_1 = -11;
				 l_2 = -17; end
		30374: begin l_1 = +11;
				 l_2 = +18; end
		22535: begin l_1 = +11;
				 l_2 = -18; end
		28326: begin l_1 = -11;
				 l_2 = +18; end
		20487: begin l_1 = -11;
				 l_2 = -18; end
		8863: begin l_1 = +11;
				 l_2 = +19; end
		44046: begin l_1 = +11;
				 l_2 = -19; end
		6815: begin l_1 = -11;
				 l_2 = +19; end
		41998: begin l_1 = -11;
				 l_2 = -19; end
		16702: begin l_1 = +11;
				 l_2 = +20; end
		36207: begin l_1 = +11;
				 l_2 = -20; end
		14654: begin l_1 = -11;
				 l_2 = +20; end
		34159: begin l_1 = -11;
				 l_2 = -20; end
		32380: begin l_1 = +11;
				 l_2 = +21; end
		20529: begin l_1 = +11;
				 l_2 = -21; end
		30332: begin l_1 = -11;
				 l_2 = +21; end
		18481: begin l_1 = -11;
				 l_2 = -21; end
		12875: begin l_1 = +11;
				 l_2 = +22; end
		40034: begin l_1 = +11;
				 l_2 = -22; end
		10827: begin l_1 = -11;
				 l_2 = +22; end
		37986: begin l_1 = -11;
				 l_2 = -22; end
		24726: begin l_1 = +11;
				 l_2 = +23; end
		28183: begin l_1 = +11;
				 l_2 = -23; end
		22678: begin l_1 = -11;
				 l_2 = +23; end
		26135: begin l_1 = -11;
				 l_2 = -23; end
		48428: begin l_1 = +11;
				 l_2 = +24; end
		4481: begin l_1 = +11;
				 l_2 = -24; end
		46380: begin l_1 = -11;
				 l_2 = +24; end
		2433: begin l_1 = -11;
				 l_2 = -24; end
		44971: begin l_1 = +11;
				 l_2 = +25; end
		7938: begin l_1 = +11;
				 l_2 = -25; end
		42923: begin l_1 = -11;
				 l_2 = +25; end
		5890: begin l_1 = -11;
				 l_2 = -25; end
		38057: begin l_1 = +11;
				 l_2 = +26; end
		14852: begin l_1 = +11;
				 l_2 = -26; end
		36009: begin l_1 = -11;
				 l_2 = +26; end
		12804: begin l_1 = -11;
				 l_2 = -26; end
		24229: begin l_1 = +11;
				 l_2 = +27; end
		28680: begin l_1 = +11;
				 l_2 = -27; end
		22181: begin l_1 = -11;
				 l_2 = +27; end
		26632: begin l_1 = -11;
				 l_2 = -27; end
		47434: begin l_1 = +11;
				 l_2 = +28; end
		5475: begin l_1 = +11;
				 l_2 = -28; end
		45386: begin l_1 = -11;
				 l_2 = +28; end
		3427: begin l_1 = -11;
				 l_2 = -28; end
		42983: begin l_1 = +11;
				 l_2 = +29; end
		9926: begin l_1 = +11;
				 l_2 = -29; end
		40935: begin l_1 = -11;
				 l_2 = +29; end
		7878: begin l_1 = -11;
				 l_2 = -29; end
		34081: begin l_1 = +11;
				 l_2 = +30; end
		18828: begin l_1 = +11;
				 l_2 = -30; end
		32033: begin l_1 = -11;
				 l_2 = +30; end
		16780: begin l_1 = -11;
				 l_2 = -30; end
		16277: begin l_1 = +11;
				 l_2 = +31; end
		36632: begin l_1 = +11;
				 l_2 = -31; end
		14229: begin l_1 = -11;
				 l_2 = +31; end
		34584: begin l_1 = -11;
				 l_2 = -31; end
		31530: begin l_1 = +11;
				 l_2 = +32; end
		21379: begin l_1 = +11;
				 l_2 = -32; end
		29482: begin l_1 = -11;
				 l_2 = +32; end
		19331: begin l_1 = -11;
				 l_2 = -32; end
		11175: begin l_1 = +11;
				 l_2 = +33; end
		41734: begin l_1 = +11;
				 l_2 = -33; end
		9127: begin l_1 = -11;
				 l_2 = +33; end
		39686: begin l_1 = -11;
				 l_2 = -33; end
		21326: begin l_1 = +11;
				 l_2 = +34; end
		31583: begin l_1 = +11;
				 l_2 = -34; end
		19278: begin l_1 = -11;
				 l_2 = +34; end
		29535: begin l_1 = -11;
				 l_2 = -34; end
		41628: begin l_1 = +11;
				 l_2 = +35; end
		11281: begin l_1 = +11;
				 l_2 = -35; end
		39580: begin l_1 = -11;
				 l_2 = +35; end
		9233: begin l_1 = -11;
				 l_2 = -35; end
		31371: begin l_1 = +11;
				 l_2 = +36; end
		21538: begin l_1 = +11;
				 l_2 = -36; end
		29323: begin l_1 = -11;
				 l_2 = +36; end
		19490: begin l_1 = -11;
				 l_2 = -36; end
		10857: begin l_1 = +11;
				 l_2 = +37; end
		42052: begin l_1 = +11;
				 l_2 = -37; end
		8809: begin l_1 = -11;
				 l_2 = +37; end
		40004: begin l_1 = -11;
				 l_2 = -37; end
		20690: begin l_1 = +11;
				 l_2 = +38; end
		32219: begin l_1 = +11;
				 l_2 = -38; end
		18642: begin l_1 = -11;
				 l_2 = +38; end
		30171: begin l_1 = -11;
				 l_2 = -38; end
		40356: begin l_1 = +11;
				 l_2 = +39; end
		12553: begin l_1 = +11;
				 l_2 = -39; end
		38308: begin l_1 = -11;
				 l_2 = +39; end
		10505: begin l_1 = -11;
				 l_2 = -39; end
		28827: begin l_1 = +11;
				 l_2 = +40; end
		24082: begin l_1 = +11;
				 l_2 = -40; end
		26779: begin l_1 = -11;
				 l_2 = +40; end
		22034: begin l_1 = -11;
				 l_2 = -40; end
		5769: begin l_1 = +11;
				 l_2 = +41; end
		47140: begin l_1 = +11;
				 l_2 = -41; end
		3721: begin l_1 = -11;
				 l_2 = +41; end
		45092: begin l_1 = -11;
				 l_2 = -41; end
		10514: begin l_1 = +11;
				 l_2 = +42; end
		42395: begin l_1 = +11;
				 l_2 = -42; end
		8466: begin l_1 = -11;
				 l_2 = +42; end
		40347: begin l_1 = -11;
				 l_2 = -42; end
		20004: begin l_1 = +11;
				 l_2 = +43; end
		32905: begin l_1 = +11;
				 l_2 = -43; end
		17956: begin l_1 = -11;
				 l_2 = +43; end
		30857: begin l_1 = -11;
				 l_2 = -43; end
		38984: begin l_1 = +11;
				 l_2 = +44; end
		13925: begin l_1 = +11;
				 l_2 = -44; end
		36936: begin l_1 = -11;
				 l_2 = +44; end
		11877: begin l_1 = -11;
				 l_2 = -44; end
		26083: begin l_1 = +11;
				 l_2 = +45; end
		26826: begin l_1 = +11;
				 l_2 = -45; end
		24035: begin l_1 = -11;
				 l_2 = +45; end
		24778: begin l_1 = -11;
				 l_2 = -45; end
		281: begin l_1 = +11;
				 l_2 = +46; end
		1767: begin l_1 = +11;
				 l_2 = -46; end
		49094: begin l_1 = -11;
				 l_2 = +46; end
		50580: begin l_1 = -11;
				 l_2 = -46; end
		50399: begin l_1 = +11;
				 l_2 = +47; end
		2510: begin l_1 = +11;
				 l_2 = -47; end
		48351: begin l_1 = -11;
				 l_2 = +47; end
		462: begin l_1 = -11;
				 l_2 = -47; end
		48913: begin l_1 = +11;
				 l_2 = +48; end
		3996: begin l_1 = +11;
				 l_2 = -48; end
		46865: begin l_1 = -11;
				 l_2 = +48; end
		1948: begin l_1 = -11;
				 l_2 = -48; end
		45941: begin l_1 = +11;
				 l_2 = +49; end
		6968: begin l_1 = +11;
				 l_2 = -49; end
		43893: begin l_1 = -11;
				 l_2 = +49; end
		4920: begin l_1 = -11;
				 l_2 = -49; end
		39997: begin l_1 = +11;
				 l_2 = +50; end
		12912: begin l_1 = +11;
				 l_2 = -50; end
		37949: begin l_1 = -11;
				 l_2 = +50; end
		10864: begin l_1 = -11;
				 l_2 = -50; end
		28109: begin l_1 = +11;
				 l_2 = +51; end
		24800: begin l_1 = +11;
				 l_2 = -51; end
		26061: begin l_1 = -11;
				 l_2 = +51; end
		22752: begin l_1 = -11;
				 l_2 = -51; end
		4333: begin l_1 = +11;
				 l_2 = +52; end
		48576: begin l_1 = +11;
				 l_2 = -52; end
		2285: begin l_1 = -11;
				 l_2 = +52; end
		46528: begin l_1 = -11;
				 l_2 = -52; end
		7642: begin l_1 = +11;
				 l_2 = +53; end
		45267: begin l_1 = +11;
				 l_2 = -53; end
		5594: begin l_1 = -11;
				 l_2 = +53; end
		43219: begin l_1 = -11;
				 l_2 = -53; end
		14260: begin l_1 = +11;
				 l_2 = +54; end
		38649: begin l_1 = +11;
				 l_2 = -54; end
		12212: begin l_1 = -11;
				 l_2 = +54; end
		36601: begin l_1 = -11;
				 l_2 = -54; end
		27496: begin l_1 = +11;
				 l_2 = +55; end
		25413: begin l_1 = +11;
				 l_2 = -55; end
		25448: begin l_1 = -11;
				 l_2 = +55; end
		23365: begin l_1 = -11;
				 l_2 = -55; end
		3107: begin l_1 = +11;
				 l_2 = +56; end
		49802: begin l_1 = +11;
				 l_2 = -56; end
		1059: begin l_1 = -11;
				 l_2 = +56; end
		47754: begin l_1 = -11;
				 l_2 = -56; end
		5190: begin l_1 = +11;
				 l_2 = +57; end
		47719: begin l_1 = +11;
				 l_2 = -57; end
		3142: begin l_1 = -11;
				 l_2 = +57; end
		45671: begin l_1 = -11;
				 l_2 = -57; end
		9356: begin l_1 = +11;
				 l_2 = +58; end
		43553: begin l_1 = +11;
				 l_2 = -58; end
		7308: begin l_1 = -11;
				 l_2 = +58; end
		41505: begin l_1 = -11;
				 l_2 = -58; end
		17688: begin l_1 = +11;
				 l_2 = +59; end
		35221: begin l_1 = +11;
				 l_2 = -59; end
		15640: begin l_1 = -11;
				 l_2 = +59; end
		33173: begin l_1 = -11;
				 l_2 = -59; end
		34352: begin l_1 = +11;
				 l_2 = +60; end
		18557: begin l_1 = +11;
				 l_2 = -60; end
		32304: begin l_1 = -11;
				 l_2 = +60; end
		16509: begin l_1 = -11;
				 l_2 = -60; end
		16819: begin l_1 = +11;
				 l_2 = +61; end
		36090: begin l_1 = +11;
				 l_2 = -61; end
		14771: begin l_1 = -11;
				 l_2 = +61; end
		34042: begin l_1 = -11;
				 l_2 = -61; end
		32614: begin l_1 = +11;
				 l_2 = +62; end
		20295: begin l_1 = +11;
				 l_2 = -62; end
		30566: begin l_1 = -11;
				 l_2 = +62; end
		18247: begin l_1 = -11;
				 l_2 = -62; end
		13343: begin l_1 = +11;
				 l_2 = +63; end
		39566: begin l_1 = +11;
				 l_2 = -63; end
		11295: begin l_1 = -11;
				 l_2 = +63; end
		37518: begin l_1 = -11;
				 l_2 = -63; end
		25662: begin l_1 = +11;
				 l_2 = +64; end
		27247: begin l_1 = +11;
				 l_2 = -64; end
		23614: begin l_1 = -11;
				 l_2 = +64; end
		25199: begin l_1 = -11;
				 l_2 = -64; end
		50300: begin l_1 = +11;
				 l_2 = +65; end
		2609: begin l_1 = +11;
				 l_2 = -65; end
		48252: begin l_1 = -11;
				 l_2 = +65; end
		561: begin l_1 = -11;
				 l_2 = -65; end
		48715: begin l_1 = +11;
				 l_2 = +66; end
		4194: begin l_1 = +11;
				 l_2 = -66; end
		46667: begin l_1 = -11;
				 l_2 = +66; end
		2146: begin l_1 = -11;
				 l_2 = -66; end
		45545: begin l_1 = +11;
				 l_2 = +67; end
		7364: begin l_1 = +11;
				 l_2 = -67; end
		43497: begin l_1 = -11;
				 l_2 = +67; end
		5316: begin l_1 = -11;
				 l_2 = -67; end
		39205: begin l_1 = +11;
				 l_2 = +68; end
		13704: begin l_1 = +11;
				 l_2 = -68; end
		37157: begin l_1 = -11;
				 l_2 = +68; end
		11656: begin l_1 = -11;
				 l_2 = -68; end
		6144: begin l_1 = -12;
				 l_2 = +14; end
		44717: begin l_1 = -12;
				 l_2 = -13; end
		10240: begin l_1 = +12;
				 l_2 = +14; end
		40621: begin l_1 = -12;
				 l_2 = -14; end
		18432: begin l_1 = +12;
				 l_2 = +15; end
		36525: begin l_1 = +12;
				 l_2 = -15; end
		14336: begin l_1 = -12;
				 l_2 = +15; end
		32429: begin l_1 = -12;
				 l_2 = -15; end
		34816: begin l_1 = +12;
				 l_2 = +16; end
		20141: begin l_1 = +12;
				 l_2 = -16; end
		30720: begin l_1 = -12;
				 l_2 = +16; end
		16045: begin l_1 = -12;
				 l_2 = -16; end
		16723: begin l_1 = +12;
				 l_2 = +17; end
		38234: begin l_1 = +12;
				 l_2 = -17; end
		12627: begin l_1 = -12;
				 l_2 = +17; end
		34138: begin l_1 = -12;
				 l_2 = -17; end
		31398: begin l_1 = +12;
				 l_2 = +18; end
		23559: begin l_1 = +12;
				 l_2 = -18; end
		27302: begin l_1 = -12;
				 l_2 = +18; end
		19463: begin l_1 = -12;
				 l_2 = -18; end
		9887: begin l_1 = +12;
				 l_2 = +19; end
		45070: begin l_1 = +12;
				 l_2 = -19; end
		5791: begin l_1 = -12;
				 l_2 = +19; end
		40974: begin l_1 = -12;
				 l_2 = -19; end
		17726: begin l_1 = +12;
				 l_2 = +20; end
		37231: begin l_1 = +12;
				 l_2 = -20; end
		13630: begin l_1 = -12;
				 l_2 = +20; end
		33135: begin l_1 = -12;
				 l_2 = -20; end
		33404: begin l_1 = +12;
				 l_2 = +21; end
		21553: begin l_1 = +12;
				 l_2 = -21; end
		29308: begin l_1 = -12;
				 l_2 = +21; end
		17457: begin l_1 = -12;
				 l_2 = -21; end
		13899: begin l_1 = +12;
				 l_2 = +22; end
		41058: begin l_1 = +12;
				 l_2 = -22; end
		9803: begin l_1 = -12;
				 l_2 = +22; end
		36962: begin l_1 = -12;
				 l_2 = -22; end
		25750: begin l_1 = +12;
				 l_2 = +23; end
		29207: begin l_1 = +12;
				 l_2 = -23; end
		21654: begin l_1 = -12;
				 l_2 = +23; end
		25111: begin l_1 = -12;
				 l_2 = -23; end
		49452: begin l_1 = +12;
				 l_2 = +24; end
		5505: begin l_1 = +12;
				 l_2 = -24; end
		45356: begin l_1 = -12;
				 l_2 = +24; end
		1409: begin l_1 = -12;
				 l_2 = -24; end
		45995: begin l_1 = +12;
				 l_2 = +25; end
		8962: begin l_1 = +12;
				 l_2 = -25; end
		41899: begin l_1 = -12;
				 l_2 = +25; end
		4866: begin l_1 = -12;
				 l_2 = -25; end
		39081: begin l_1 = +12;
				 l_2 = +26; end
		15876: begin l_1 = +12;
				 l_2 = -26; end
		34985: begin l_1 = -12;
				 l_2 = +26; end
		11780: begin l_1 = -12;
				 l_2 = -26; end
		25253: begin l_1 = +12;
				 l_2 = +27; end
		29704: begin l_1 = +12;
				 l_2 = -27; end
		21157: begin l_1 = -12;
				 l_2 = +27; end
		25608: begin l_1 = -12;
				 l_2 = -27; end
		48458: begin l_1 = +12;
				 l_2 = +28; end
		6499: begin l_1 = +12;
				 l_2 = -28; end
		44362: begin l_1 = -12;
				 l_2 = +28; end
		2403: begin l_1 = -12;
				 l_2 = -28; end
		44007: begin l_1 = +12;
				 l_2 = +29; end
		10950: begin l_1 = +12;
				 l_2 = -29; end
		39911: begin l_1 = -12;
				 l_2 = +29; end
		6854: begin l_1 = -12;
				 l_2 = -29; end
		35105: begin l_1 = +12;
				 l_2 = +30; end
		19852: begin l_1 = +12;
				 l_2 = -30; end
		31009: begin l_1 = -12;
				 l_2 = +30; end
		15756: begin l_1 = -12;
				 l_2 = -30; end
		17301: begin l_1 = +12;
				 l_2 = +31; end
		37656: begin l_1 = +12;
				 l_2 = -31; end
		13205: begin l_1 = -12;
				 l_2 = +31; end
		33560: begin l_1 = -12;
				 l_2 = -31; end
		32554: begin l_1 = +12;
				 l_2 = +32; end
		22403: begin l_1 = +12;
				 l_2 = -32; end
		28458: begin l_1 = -12;
				 l_2 = +32; end
		18307: begin l_1 = -12;
				 l_2 = -32; end
		12199: begin l_1 = +12;
				 l_2 = +33; end
		42758: begin l_1 = +12;
				 l_2 = -33; end
		8103: begin l_1 = -12;
				 l_2 = +33; end
		38662: begin l_1 = -12;
				 l_2 = -33; end
		22350: begin l_1 = +12;
				 l_2 = +34; end
		32607: begin l_1 = +12;
				 l_2 = -34; end
		18254: begin l_1 = -12;
				 l_2 = +34; end
		28511: begin l_1 = -12;
				 l_2 = -34; end
		42652: begin l_1 = +12;
				 l_2 = +35; end
		12305: begin l_1 = +12;
				 l_2 = -35; end
		38556: begin l_1 = -12;
				 l_2 = +35; end
		8209: begin l_1 = -12;
				 l_2 = -35; end
		32395: begin l_1 = +12;
				 l_2 = +36; end
		22562: begin l_1 = +12;
				 l_2 = -36; end
		28299: begin l_1 = -12;
				 l_2 = +36; end
		18466: begin l_1 = -12;
				 l_2 = -36; end
		11881: begin l_1 = +12;
				 l_2 = +37; end
		43076: begin l_1 = +12;
				 l_2 = -37; end
		7785: begin l_1 = -12;
				 l_2 = +37; end
		38980: begin l_1 = -12;
				 l_2 = -37; end
		21714: begin l_1 = +12;
				 l_2 = +38; end
		33243: begin l_1 = +12;
				 l_2 = -38; end
		17618: begin l_1 = -12;
				 l_2 = +38; end
		29147: begin l_1 = -12;
				 l_2 = -38; end
		41380: begin l_1 = +12;
				 l_2 = +39; end
		13577: begin l_1 = +12;
				 l_2 = -39; end
		37284: begin l_1 = -12;
				 l_2 = +39; end
		9481: begin l_1 = -12;
				 l_2 = -39; end
		29851: begin l_1 = +12;
				 l_2 = +40; end
		25106: begin l_1 = +12;
				 l_2 = -40; end
		25755: begin l_1 = -12;
				 l_2 = +40; end
		21010: begin l_1 = -12;
				 l_2 = -40; end
		6793: begin l_1 = +12;
				 l_2 = +41; end
		48164: begin l_1 = +12;
				 l_2 = -41; end
		2697: begin l_1 = -12;
				 l_2 = +41; end
		44068: begin l_1 = -12;
				 l_2 = -41; end
		11538: begin l_1 = +12;
				 l_2 = +42; end
		43419: begin l_1 = +12;
				 l_2 = -42; end
		7442: begin l_1 = -12;
				 l_2 = +42; end
		39323: begin l_1 = -12;
				 l_2 = -42; end
		21028: begin l_1 = +12;
				 l_2 = +43; end
		33929: begin l_1 = +12;
				 l_2 = -43; end
		16932: begin l_1 = -12;
				 l_2 = +43; end
		29833: begin l_1 = -12;
				 l_2 = -43; end
		40008: begin l_1 = +12;
				 l_2 = +44; end
		14949: begin l_1 = +12;
				 l_2 = -44; end
		35912: begin l_1 = -12;
				 l_2 = +44; end
		10853: begin l_1 = -12;
				 l_2 = -44; end
		27107: begin l_1 = +12;
				 l_2 = +45; end
		27850: begin l_1 = +12;
				 l_2 = -45; end
		23011: begin l_1 = -12;
				 l_2 = +45; end
		23754: begin l_1 = -12;
				 l_2 = -45; end
		1305: begin l_1 = +12;
				 l_2 = +46; end
		2791: begin l_1 = +12;
				 l_2 = -46; end
		48070: begin l_1 = -12;
				 l_2 = +46; end
		49556: begin l_1 = -12;
				 l_2 = -46; end
		562: begin l_1 = +12;
				 l_2 = +47; end
		3534: begin l_1 = +12;
				 l_2 = -47; end
		47327: begin l_1 = -12;
				 l_2 = +47; end
		50299: begin l_1 = -12;
				 l_2 = -47; end
		49937: begin l_1 = +12;
				 l_2 = +48; end
		5020: begin l_1 = +12;
				 l_2 = -48; end
		45841: begin l_1 = -12;
				 l_2 = +48; end
		924: begin l_1 = -12;
				 l_2 = -48; end
		46965: begin l_1 = +12;
				 l_2 = +49; end
		7992: begin l_1 = +12;
				 l_2 = -49; end
		42869: begin l_1 = -12;
				 l_2 = +49; end
		3896: begin l_1 = -12;
				 l_2 = -49; end
		41021: begin l_1 = +12;
				 l_2 = +50; end
		13936: begin l_1 = +12;
				 l_2 = -50; end
		36925: begin l_1 = -12;
				 l_2 = +50; end
		9840: begin l_1 = -12;
				 l_2 = -50; end
		29133: begin l_1 = +12;
				 l_2 = +51; end
		25824: begin l_1 = +12;
				 l_2 = -51; end
		25037: begin l_1 = -12;
				 l_2 = +51; end
		21728: begin l_1 = -12;
				 l_2 = -51; end
		5357: begin l_1 = +12;
				 l_2 = +52; end
		49600: begin l_1 = +12;
				 l_2 = -52; end
		1261: begin l_1 = -12;
				 l_2 = +52; end
		45504: begin l_1 = -12;
				 l_2 = -52; end
		8666: begin l_1 = +12;
				 l_2 = +53; end
		46291: begin l_1 = +12;
				 l_2 = -53; end
		4570: begin l_1 = -12;
				 l_2 = +53; end
		42195: begin l_1 = -12;
				 l_2 = -53; end
		15284: begin l_1 = +12;
				 l_2 = +54; end
		39673: begin l_1 = +12;
				 l_2 = -54; end
		11188: begin l_1 = -12;
				 l_2 = +54; end
		35577: begin l_1 = -12;
				 l_2 = -54; end
		28520: begin l_1 = +12;
				 l_2 = +55; end
		26437: begin l_1 = +12;
				 l_2 = -55; end
		24424: begin l_1 = -12;
				 l_2 = +55; end
		22341: begin l_1 = -12;
				 l_2 = -55; end
		4131: begin l_1 = +12;
				 l_2 = +56; end
		50826: begin l_1 = +12;
				 l_2 = -56; end
		35: begin l_1 = -12;
				 l_2 = +56; end
		46730: begin l_1 = -12;
				 l_2 = -56; end
		6214: begin l_1 = +12;
				 l_2 = +57; end
		48743: begin l_1 = +12;
				 l_2 = -57; end
		2118: begin l_1 = -12;
				 l_2 = +57; end
		44647: begin l_1 = -12;
				 l_2 = -57; end
		10380: begin l_1 = +12;
				 l_2 = +58; end
		44577: begin l_1 = +12;
				 l_2 = -58; end
		6284: begin l_1 = -12;
				 l_2 = +58; end
		40481: begin l_1 = -12;
				 l_2 = -58; end
		18712: begin l_1 = +12;
				 l_2 = +59; end
		36245: begin l_1 = +12;
				 l_2 = -59; end
		14616: begin l_1 = -12;
				 l_2 = +59; end
		32149: begin l_1 = -12;
				 l_2 = -59; end
		35376: begin l_1 = +12;
				 l_2 = +60; end
		19581: begin l_1 = +12;
				 l_2 = -60; end
		31280: begin l_1 = -12;
				 l_2 = +60; end
		15485: begin l_1 = -12;
				 l_2 = -60; end
		17843: begin l_1 = +12;
				 l_2 = +61; end
		37114: begin l_1 = +12;
				 l_2 = -61; end
		13747: begin l_1 = -12;
				 l_2 = +61; end
		33018: begin l_1 = -12;
				 l_2 = -61; end
		33638: begin l_1 = +12;
				 l_2 = +62; end
		21319: begin l_1 = +12;
				 l_2 = -62; end
		29542: begin l_1 = -12;
				 l_2 = +62; end
		17223: begin l_1 = -12;
				 l_2 = -62; end
		14367: begin l_1 = +12;
				 l_2 = +63; end
		40590: begin l_1 = +12;
				 l_2 = -63; end
		10271: begin l_1 = -12;
				 l_2 = +63; end
		36494: begin l_1 = -12;
				 l_2 = -63; end
		26686: begin l_1 = +12;
				 l_2 = +64; end
		28271: begin l_1 = +12;
				 l_2 = -64; end
		22590: begin l_1 = -12;
				 l_2 = +64; end
		24175: begin l_1 = -12;
				 l_2 = -64; end
		463: begin l_1 = +12;
				 l_2 = +65; end
		3633: begin l_1 = +12;
				 l_2 = -65; end
		47228: begin l_1 = -12;
				 l_2 = +65; end
		50398: begin l_1 = -12;
				 l_2 = -65; end
		49739: begin l_1 = +12;
				 l_2 = +66; end
		5218: begin l_1 = +12;
				 l_2 = -66; end
		45643: begin l_1 = -12;
				 l_2 = +66; end
		1122: begin l_1 = -12;
				 l_2 = -66; end
		46569: begin l_1 = +12;
				 l_2 = +67; end
		8388: begin l_1 = +12;
				 l_2 = -67; end
		42473: begin l_1 = -12;
				 l_2 = +67; end
		4292: begin l_1 = -12;
				 l_2 = -67; end
		40229: begin l_1 = +12;
				 l_2 = +68; end
		14728: begin l_1 = +12;
				 l_2 = -68; end
		36133: begin l_1 = -12;
				 l_2 = +68; end
		10632: begin l_1 = -12;
				 l_2 = -68; end
		12288: begin l_1 = -13;
				 l_2 = +15; end
		38573: begin l_1 = -13;
				 l_2 = -14; end
		20480: begin l_1 = +13;
				 l_2 = +15; end
		30381: begin l_1 = -13;
				 l_2 = -15; end
		36864: begin l_1 = +13;
				 l_2 = +16; end
		22189: begin l_1 = +13;
				 l_2 = -16; end
		28672: begin l_1 = -13;
				 l_2 = +16; end
		13997: begin l_1 = -13;
				 l_2 = -16; end
		18771: begin l_1 = +13;
				 l_2 = +17; end
		40282: begin l_1 = +13;
				 l_2 = -17; end
		10579: begin l_1 = -13;
				 l_2 = +17; end
		32090: begin l_1 = -13;
				 l_2 = -17; end
		33446: begin l_1 = +13;
				 l_2 = +18; end
		25607: begin l_1 = +13;
				 l_2 = -18; end
		25254: begin l_1 = -13;
				 l_2 = +18; end
		17415: begin l_1 = -13;
				 l_2 = -18; end
		11935: begin l_1 = +13;
				 l_2 = +19; end
		47118: begin l_1 = +13;
				 l_2 = -19; end
		3743: begin l_1 = -13;
				 l_2 = +19; end
		38926: begin l_1 = -13;
				 l_2 = -19; end
		19774: begin l_1 = +13;
				 l_2 = +20; end
		39279: begin l_1 = +13;
				 l_2 = -20; end
		11582: begin l_1 = -13;
				 l_2 = +20; end
		31087: begin l_1 = -13;
				 l_2 = -20; end
		35452: begin l_1 = +13;
				 l_2 = +21; end
		23601: begin l_1 = +13;
				 l_2 = -21; end
		27260: begin l_1 = -13;
				 l_2 = +21; end
		15409: begin l_1 = -13;
				 l_2 = -21; end
		15947: begin l_1 = +13;
				 l_2 = +22; end
		43106: begin l_1 = +13;
				 l_2 = -22; end
		7755: begin l_1 = -13;
				 l_2 = +22; end
		34914: begin l_1 = -13;
				 l_2 = -22; end
		27798: begin l_1 = +13;
				 l_2 = +23; end
		31255: begin l_1 = +13;
				 l_2 = -23; end
		19606: begin l_1 = -13;
				 l_2 = +23; end
		23063: begin l_1 = -13;
				 l_2 = -23; end
		639: begin l_1 = +13;
				 l_2 = +24; end
		7553: begin l_1 = +13;
				 l_2 = -24; end
		43308: begin l_1 = -13;
				 l_2 = +24; end
		50222: begin l_1 = -13;
				 l_2 = -24; end
		48043: begin l_1 = +13;
				 l_2 = +25; end
		11010: begin l_1 = +13;
				 l_2 = -25; end
		39851: begin l_1 = -13;
				 l_2 = +25; end
		2818: begin l_1 = -13;
				 l_2 = -25; end
		41129: begin l_1 = +13;
				 l_2 = +26; end
		17924: begin l_1 = +13;
				 l_2 = -26; end
		32937: begin l_1 = -13;
				 l_2 = +26; end
		9732: begin l_1 = -13;
				 l_2 = -26; end
		27301: begin l_1 = +13;
				 l_2 = +27; end
		31752: begin l_1 = +13;
				 l_2 = -27; end
		19109: begin l_1 = -13;
				 l_2 = +27; end
		23560: begin l_1 = -13;
				 l_2 = -27; end
		50506: begin l_1 = +13;
				 l_2 = +28; end
		8547: begin l_1 = +13;
				 l_2 = -28; end
		42314: begin l_1 = -13;
				 l_2 = +28; end
		355: begin l_1 = -13;
				 l_2 = -28; end
		46055: begin l_1 = +13;
				 l_2 = +29; end
		12998: begin l_1 = +13;
				 l_2 = -29; end
		37863: begin l_1 = -13;
				 l_2 = +29; end
		4806: begin l_1 = -13;
				 l_2 = -29; end
		37153: begin l_1 = +13;
				 l_2 = +30; end
		21900: begin l_1 = +13;
				 l_2 = -30; end
		28961: begin l_1 = -13;
				 l_2 = +30; end
		13708: begin l_1 = -13;
				 l_2 = -30; end
		19349: begin l_1 = +13;
				 l_2 = +31; end
		39704: begin l_1 = +13;
				 l_2 = -31; end
		11157: begin l_1 = -13;
				 l_2 = +31; end
		31512: begin l_1 = -13;
				 l_2 = -31; end
		34602: begin l_1 = +13;
				 l_2 = +32; end
		24451: begin l_1 = +13;
				 l_2 = -32; end
		26410: begin l_1 = -13;
				 l_2 = +32; end
		16259: begin l_1 = -13;
				 l_2 = -32; end
		14247: begin l_1 = +13;
				 l_2 = +33; end
		44806: begin l_1 = +13;
				 l_2 = -33; end
		6055: begin l_1 = -13;
				 l_2 = +33; end
		36614: begin l_1 = -13;
				 l_2 = -33; end
		24398: begin l_1 = +13;
				 l_2 = +34; end
		34655: begin l_1 = +13;
				 l_2 = -34; end
		16206: begin l_1 = -13;
				 l_2 = +34; end
		26463: begin l_1 = -13;
				 l_2 = -34; end
		44700: begin l_1 = +13;
				 l_2 = +35; end
		14353: begin l_1 = +13;
				 l_2 = -35; end
		36508: begin l_1 = -13;
				 l_2 = +35; end
		6161: begin l_1 = -13;
				 l_2 = -35; end
		34443: begin l_1 = +13;
				 l_2 = +36; end
		24610: begin l_1 = +13;
				 l_2 = -36; end
		26251: begin l_1 = -13;
				 l_2 = +36; end
		16418: begin l_1 = -13;
				 l_2 = -36; end
		13929: begin l_1 = +13;
				 l_2 = +37; end
		45124: begin l_1 = +13;
				 l_2 = -37; end
		5737: begin l_1 = -13;
				 l_2 = +37; end
		36932: begin l_1 = -13;
				 l_2 = -37; end
		23762: begin l_1 = +13;
				 l_2 = +38; end
		35291: begin l_1 = +13;
				 l_2 = -38; end
		15570: begin l_1 = -13;
				 l_2 = +38; end
		27099: begin l_1 = -13;
				 l_2 = -38; end
		43428: begin l_1 = +13;
				 l_2 = +39; end
		15625: begin l_1 = +13;
				 l_2 = -39; end
		35236: begin l_1 = -13;
				 l_2 = +39; end
		7433: begin l_1 = -13;
				 l_2 = -39; end
		31899: begin l_1 = +13;
				 l_2 = +40; end
		27154: begin l_1 = +13;
				 l_2 = -40; end
		23707: begin l_1 = -13;
				 l_2 = +40; end
		18962: begin l_1 = -13;
				 l_2 = -40; end
		8841: begin l_1 = +13;
				 l_2 = +41; end
		50212: begin l_1 = +13;
				 l_2 = -41; end
		649: begin l_1 = -13;
				 l_2 = +41; end
		42020: begin l_1 = -13;
				 l_2 = -41; end
		13586: begin l_1 = +13;
				 l_2 = +42; end
		45467: begin l_1 = +13;
				 l_2 = -42; end
		5394: begin l_1 = -13;
				 l_2 = +42; end
		37275: begin l_1 = -13;
				 l_2 = -42; end
		23076: begin l_1 = +13;
				 l_2 = +43; end
		35977: begin l_1 = +13;
				 l_2 = -43; end
		14884: begin l_1 = -13;
				 l_2 = +43; end
		27785: begin l_1 = -13;
				 l_2 = -43; end
		42056: begin l_1 = +13;
				 l_2 = +44; end
		16997: begin l_1 = +13;
				 l_2 = -44; end
		33864: begin l_1 = -13;
				 l_2 = +44; end
		8805: begin l_1 = -13;
				 l_2 = -44; end
		29155: begin l_1 = +13;
				 l_2 = +45; end
		29898: begin l_1 = +13;
				 l_2 = -45; end
		20963: begin l_1 = -13;
				 l_2 = +45; end
		21706: begin l_1 = -13;
				 l_2 = -45; end
		3353: begin l_1 = +13;
				 l_2 = +46; end
		4839: begin l_1 = +13;
				 l_2 = -46; end
		46022: begin l_1 = -13;
				 l_2 = +46; end
		47508: begin l_1 = -13;
				 l_2 = -46; end
		2610: begin l_1 = +13;
				 l_2 = +47; end
		5582: begin l_1 = +13;
				 l_2 = -47; end
		45279: begin l_1 = -13;
				 l_2 = +47; end
		48251: begin l_1 = -13;
				 l_2 = -47; end
		1124: begin l_1 = +13;
				 l_2 = +48; end
		7068: begin l_1 = +13;
				 l_2 = -48; end
		43793: begin l_1 = -13;
				 l_2 = +48; end
		49737: begin l_1 = -13;
				 l_2 = -48; end
		49013: begin l_1 = +13;
				 l_2 = +49; end
		10040: begin l_1 = +13;
				 l_2 = -49; end
		40821: begin l_1 = -13;
				 l_2 = +49; end
		1848: begin l_1 = -13;
				 l_2 = -49; end
		43069: begin l_1 = +13;
				 l_2 = +50; end
		15984: begin l_1 = +13;
				 l_2 = -50; end
		34877: begin l_1 = -13;
				 l_2 = +50; end
		7792: begin l_1 = -13;
				 l_2 = -50; end
		31181: begin l_1 = +13;
				 l_2 = +51; end
		27872: begin l_1 = +13;
				 l_2 = -51; end
		22989: begin l_1 = -13;
				 l_2 = +51; end
		19680: begin l_1 = -13;
				 l_2 = -51; end
		7405: begin l_1 = +13;
				 l_2 = +52; end
		787: begin l_1 = +13;
				 l_2 = -52; end
		50074: begin l_1 = -13;
				 l_2 = +52; end
		43456: begin l_1 = -13;
				 l_2 = -52; end
		10714: begin l_1 = +13;
				 l_2 = +53; end
		48339: begin l_1 = +13;
				 l_2 = -53; end
		2522: begin l_1 = -13;
				 l_2 = +53; end
		40147: begin l_1 = -13;
				 l_2 = -53; end
		17332: begin l_1 = +13;
				 l_2 = +54; end
		41721: begin l_1 = +13;
				 l_2 = -54; end
		9140: begin l_1 = -13;
				 l_2 = +54; end
		33529: begin l_1 = -13;
				 l_2 = -54; end
		30568: begin l_1 = +13;
				 l_2 = +55; end
		28485: begin l_1 = +13;
				 l_2 = -55; end
		22376: begin l_1 = -13;
				 l_2 = +55; end
		20293: begin l_1 = -13;
				 l_2 = -55; end
		6179: begin l_1 = +13;
				 l_2 = +56; end
		2013: begin l_1 = +13;
				 l_2 = -56; end
		48848: begin l_1 = -13;
				 l_2 = +56; end
		44682: begin l_1 = -13;
				 l_2 = -56; end
		8262: begin l_1 = +13;
				 l_2 = +57; end
		50791: begin l_1 = +13;
				 l_2 = -57; end
		70: begin l_1 = -13;
				 l_2 = +57; end
		42599: begin l_1 = -13;
				 l_2 = -57; end
		12428: begin l_1 = +13;
				 l_2 = +58; end
		46625: begin l_1 = +13;
				 l_2 = -58; end
		4236: begin l_1 = -13;
				 l_2 = +58; end
		38433: begin l_1 = -13;
				 l_2 = -58; end
		20760: begin l_1 = +13;
				 l_2 = +59; end
		38293: begin l_1 = +13;
				 l_2 = -59; end
		12568: begin l_1 = -13;
				 l_2 = +59; end
		30101: begin l_1 = -13;
				 l_2 = -59; end
		37424: begin l_1 = +13;
				 l_2 = +60; end
		21629: begin l_1 = +13;
				 l_2 = -60; end
		29232: begin l_1 = -13;
				 l_2 = +60; end
		13437: begin l_1 = -13;
				 l_2 = -60; end
		19891: begin l_1 = +13;
				 l_2 = +61; end
		39162: begin l_1 = +13;
				 l_2 = -61; end
		11699: begin l_1 = -13;
				 l_2 = +61; end
		30970: begin l_1 = -13;
				 l_2 = -61; end
		35686: begin l_1 = +13;
				 l_2 = +62; end
		23367: begin l_1 = +13;
				 l_2 = -62; end
		27494: begin l_1 = -13;
				 l_2 = +62; end
		15175: begin l_1 = -13;
				 l_2 = -62; end
		16415: begin l_1 = +13;
				 l_2 = +63; end
		42638: begin l_1 = +13;
				 l_2 = -63; end
		8223: begin l_1 = -13;
				 l_2 = +63; end
		34446: begin l_1 = -13;
				 l_2 = -63; end
		28734: begin l_1 = +13;
				 l_2 = +64; end
		30319: begin l_1 = +13;
				 l_2 = -64; end
		20542: begin l_1 = -13;
				 l_2 = +64; end
		22127: begin l_1 = -13;
				 l_2 = -64; end
		2511: begin l_1 = +13;
				 l_2 = +65; end
		5681: begin l_1 = +13;
				 l_2 = -65; end
		45180: begin l_1 = -13;
				 l_2 = +65; end
		48350: begin l_1 = -13;
				 l_2 = -65; end
		926: begin l_1 = +13;
				 l_2 = +66; end
		7266: begin l_1 = +13;
				 l_2 = -66; end
		43595: begin l_1 = -13;
				 l_2 = +66; end
		49935: begin l_1 = -13;
				 l_2 = -66; end
		48617: begin l_1 = +13;
				 l_2 = +67; end
		10436: begin l_1 = +13;
				 l_2 = -67; end
		40425: begin l_1 = -13;
				 l_2 = +67; end
		2244: begin l_1 = -13;
				 l_2 = -67; end
		42277: begin l_1 = +13;
				 l_2 = +68; end
		16776: begin l_1 = +13;
				 l_2 = -68; end
		34085: begin l_1 = -13;
				 l_2 = +68; end
		8584: begin l_1 = -13;
				 l_2 = -68; end
		24576: begin l_1 = -14;
				 l_2 = +16; end
		26285: begin l_1 = -14;
				 l_2 = -15; end
		40960: begin l_1 = +14;
				 l_2 = +16; end
		9901: begin l_1 = -14;
				 l_2 = -16; end
		22867: begin l_1 = +14;
				 l_2 = +17; end
		44378: begin l_1 = +14;
				 l_2 = -17; end
		6483: begin l_1 = -14;
				 l_2 = +17; end
		27994: begin l_1 = -14;
				 l_2 = -17; end
		37542: begin l_1 = +14;
				 l_2 = +18; end
		29703: begin l_1 = +14;
				 l_2 = -18; end
		21158: begin l_1 = -14;
				 l_2 = +18; end
		13319: begin l_1 = -14;
				 l_2 = -18; end
		16031: begin l_1 = +14;
				 l_2 = +19; end
		353: begin l_1 = +14;
				 l_2 = -19; end
		50508: begin l_1 = -14;
				 l_2 = +19; end
		34830: begin l_1 = -14;
				 l_2 = -19; end
		23870: begin l_1 = +14;
				 l_2 = +20; end
		43375: begin l_1 = +14;
				 l_2 = -20; end
		7486: begin l_1 = -14;
				 l_2 = +20; end
		26991: begin l_1 = -14;
				 l_2 = -20; end
		39548: begin l_1 = +14;
				 l_2 = +21; end
		27697: begin l_1 = +14;
				 l_2 = -21; end
		23164: begin l_1 = -14;
				 l_2 = +21; end
		11313: begin l_1 = -14;
				 l_2 = -21; end
		20043: begin l_1 = +14;
				 l_2 = +22; end
		47202: begin l_1 = +14;
				 l_2 = -22; end
		3659: begin l_1 = -14;
				 l_2 = +22; end
		30818: begin l_1 = -14;
				 l_2 = -22; end
		31894: begin l_1 = +14;
				 l_2 = +23; end
		35351: begin l_1 = +14;
				 l_2 = -23; end
		15510: begin l_1 = -14;
				 l_2 = +23; end
		18967: begin l_1 = -14;
				 l_2 = -23; end
		4735: begin l_1 = +14;
				 l_2 = +24; end
		11649: begin l_1 = +14;
				 l_2 = -24; end
		39212: begin l_1 = -14;
				 l_2 = +24; end
		46126: begin l_1 = -14;
				 l_2 = -24; end
		1278: begin l_1 = +14;
				 l_2 = +25; end
		15106: begin l_1 = +14;
				 l_2 = -25; end
		35755: begin l_1 = -14;
				 l_2 = +25; end
		49583: begin l_1 = -14;
				 l_2 = -25; end
		45225: begin l_1 = +14;
				 l_2 = +26; end
		22020: begin l_1 = +14;
				 l_2 = -26; end
		28841: begin l_1 = -14;
				 l_2 = +26; end
		5636: begin l_1 = -14;
				 l_2 = -26; end
		31397: begin l_1 = +14;
				 l_2 = +27; end
		35848: begin l_1 = +14;
				 l_2 = -27; end
		15013: begin l_1 = -14;
				 l_2 = +27; end
		19464: begin l_1 = -14;
				 l_2 = -27; end
		3741: begin l_1 = +14;
				 l_2 = +28; end
		12643: begin l_1 = +14;
				 l_2 = -28; end
		38218: begin l_1 = -14;
				 l_2 = +28; end
		47120: begin l_1 = -14;
				 l_2 = -28; end
		50151: begin l_1 = +14;
				 l_2 = +29; end
		17094: begin l_1 = +14;
				 l_2 = -29; end
		33767: begin l_1 = -14;
				 l_2 = +29; end
		710: begin l_1 = -14;
				 l_2 = -29; end
		41249: begin l_1 = +14;
				 l_2 = +30; end
		25996: begin l_1 = +14;
				 l_2 = -30; end
		24865: begin l_1 = -14;
				 l_2 = +30; end
		9612: begin l_1 = -14;
				 l_2 = -30; end
		23445: begin l_1 = +14;
				 l_2 = +31; end
		43800: begin l_1 = +14;
				 l_2 = -31; end
		7061: begin l_1 = -14;
				 l_2 = +31; end
		27416: begin l_1 = -14;
				 l_2 = -31; end
		38698: begin l_1 = +14;
				 l_2 = +32; end
		28547: begin l_1 = +14;
				 l_2 = -32; end
		22314: begin l_1 = -14;
				 l_2 = +32; end
		12163: begin l_1 = -14;
				 l_2 = -32; end
		18343: begin l_1 = +14;
				 l_2 = +33; end
		48902: begin l_1 = +14;
				 l_2 = -33; end
		1959: begin l_1 = -14;
				 l_2 = +33; end
		32518: begin l_1 = -14;
				 l_2 = -33; end
		28494: begin l_1 = +14;
				 l_2 = +34; end
		38751: begin l_1 = +14;
				 l_2 = -34; end
		12110: begin l_1 = -14;
				 l_2 = +34; end
		22367: begin l_1 = -14;
				 l_2 = -34; end
		48796: begin l_1 = +14;
				 l_2 = +35; end
		18449: begin l_1 = +14;
				 l_2 = -35; end
		32412: begin l_1 = -14;
				 l_2 = +35; end
		2065: begin l_1 = -14;
				 l_2 = -35; end
		38539: begin l_1 = +14;
				 l_2 = +36; end
		28706: begin l_1 = +14;
				 l_2 = -36; end
		22155: begin l_1 = -14;
				 l_2 = +36; end
		12322: begin l_1 = -14;
				 l_2 = -36; end
		18025: begin l_1 = +14;
				 l_2 = +37; end
		49220: begin l_1 = +14;
				 l_2 = -37; end
		1641: begin l_1 = -14;
				 l_2 = +37; end
		32836: begin l_1 = -14;
				 l_2 = -37; end
		27858: begin l_1 = +14;
				 l_2 = +38; end
		39387: begin l_1 = +14;
				 l_2 = -38; end
		11474: begin l_1 = -14;
				 l_2 = +38; end
		23003: begin l_1 = -14;
				 l_2 = -38; end
		47524: begin l_1 = +14;
				 l_2 = +39; end
		19721: begin l_1 = +14;
				 l_2 = -39; end
		31140: begin l_1 = -14;
				 l_2 = +39; end
		3337: begin l_1 = -14;
				 l_2 = -39; end
		35995: begin l_1 = +14;
				 l_2 = +40; end
		31250: begin l_1 = +14;
				 l_2 = -40; end
		19611: begin l_1 = -14;
				 l_2 = +40; end
		14866: begin l_1 = -14;
				 l_2 = -40; end
		12937: begin l_1 = +14;
				 l_2 = +41; end
		3447: begin l_1 = +14;
				 l_2 = -41; end
		47414: begin l_1 = -14;
				 l_2 = +41; end
		37924: begin l_1 = -14;
				 l_2 = -41; end
		17682: begin l_1 = +14;
				 l_2 = +42; end
		49563: begin l_1 = +14;
				 l_2 = -42; end
		1298: begin l_1 = -14;
				 l_2 = +42; end
		33179: begin l_1 = -14;
				 l_2 = -42; end
		27172: begin l_1 = +14;
				 l_2 = +43; end
		40073: begin l_1 = +14;
				 l_2 = -43; end
		10788: begin l_1 = -14;
				 l_2 = +43; end
		23689: begin l_1 = -14;
				 l_2 = -43; end
		46152: begin l_1 = +14;
				 l_2 = +44; end
		21093: begin l_1 = +14;
				 l_2 = -44; end
		29768: begin l_1 = -14;
				 l_2 = +44; end
		4709: begin l_1 = -14;
				 l_2 = -44; end
		33251: begin l_1 = +14;
				 l_2 = +45; end
		33994: begin l_1 = +14;
				 l_2 = -45; end
		16867: begin l_1 = -14;
				 l_2 = +45; end
		17610: begin l_1 = -14;
				 l_2 = -45; end
		7449: begin l_1 = +14;
				 l_2 = +46; end
		8935: begin l_1 = +14;
				 l_2 = -46; end
		41926: begin l_1 = -14;
				 l_2 = +46; end
		43412: begin l_1 = -14;
				 l_2 = -46; end
		6706: begin l_1 = +14;
				 l_2 = +47; end
		9678: begin l_1 = +14;
				 l_2 = -47; end
		41183: begin l_1 = -14;
				 l_2 = +47; end
		44155: begin l_1 = -14;
				 l_2 = -47; end
		5220: begin l_1 = +14;
				 l_2 = +48; end
		11164: begin l_1 = +14;
				 l_2 = -48; end
		39697: begin l_1 = -14;
				 l_2 = +48; end
		45641: begin l_1 = -14;
				 l_2 = -48; end
		2248: begin l_1 = +14;
				 l_2 = +49; end
		14136: begin l_1 = +14;
				 l_2 = -49; end
		36725: begin l_1 = -14;
				 l_2 = +49; end
		48613: begin l_1 = -14;
				 l_2 = -49; end
		47165: begin l_1 = +14;
				 l_2 = +50; end
		20080: begin l_1 = +14;
				 l_2 = -50; end
		30781: begin l_1 = -14;
				 l_2 = +50; end
		3696: begin l_1 = -14;
				 l_2 = -50; end
		35277: begin l_1 = +14;
				 l_2 = +51; end
		31968: begin l_1 = +14;
				 l_2 = -51; end
		18893: begin l_1 = -14;
				 l_2 = +51; end
		15584: begin l_1 = -14;
				 l_2 = -51; end
		11501: begin l_1 = +14;
				 l_2 = +52; end
		4883: begin l_1 = +14;
				 l_2 = -52; end
		45978: begin l_1 = -14;
				 l_2 = +52; end
		39360: begin l_1 = -14;
				 l_2 = -52; end
		14810: begin l_1 = +14;
				 l_2 = +53; end
		1574: begin l_1 = +14;
				 l_2 = -53; end
		49287: begin l_1 = -14;
				 l_2 = +53; end
		36051: begin l_1 = -14;
				 l_2 = -53; end
		21428: begin l_1 = +14;
				 l_2 = +54; end
		45817: begin l_1 = +14;
				 l_2 = -54; end
		5044: begin l_1 = -14;
				 l_2 = +54; end
		29433: begin l_1 = -14;
				 l_2 = -54; end
		34664: begin l_1 = +14;
				 l_2 = +55; end
		32581: begin l_1 = +14;
				 l_2 = -55; end
		18280: begin l_1 = -14;
				 l_2 = +55; end
		16197: begin l_1 = -14;
				 l_2 = -55; end
		10275: begin l_1 = +14;
				 l_2 = +56; end
		6109: begin l_1 = +14;
				 l_2 = -56; end
		44752: begin l_1 = -14;
				 l_2 = +56; end
		40586: begin l_1 = -14;
				 l_2 = -56; end
		12358: begin l_1 = +14;
				 l_2 = +57; end
		4026: begin l_1 = +14;
				 l_2 = -57; end
		46835: begin l_1 = -14;
				 l_2 = +57; end
		38503: begin l_1 = -14;
				 l_2 = -57; end
		16524: begin l_1 = +14;
				 l_2 = +58; end
		50721: begin l_1 = +14;
				 l_2 = -58; end
		140: begin l_1 = -14;
				 l_2 = +58; end
		34337: begin l_1 = -14;
				 l_2 = -58; end
		24856: begin l_1 = +14;
				 l_2 = +59; end
		42389: begin l_1 = +14;
				 l_2 = -59; end
		8472: begin l_1 = -14;
				 l_2 = +59; end
		26005: begin l_1 = -14;
				 l_2 = -59; end
		41520: begin l_1 = +14;
				 l_2 = +60; end
		25725: begin l_1 = +14;
				 l_2 = -60; end
		25136: begin l_1 = -14;
				 l_2 = +60; end
		9341: begin l_1 = -14;
				 l_2 = -60; end
		23987: begin l_1 = +14;
				 l_2 = +61; end
		43258: begin l_1 = +14;
				 l_2 = -61; end
		7603: begin l_1 = -14;
				 l_2 = +61; end
		26874: begin l_1 = -14;
				 l_2 = -61; end
		39782: begin l_1 = +14;
				 l_2 = +62; end
		27463: begin l_1 = +14;
				 l_2 = -62; end
		23398: begin l_1 = -14;
				 l_2 = +62; end
		11079: begin l_1 = -14;
				 l_2 = -62; end
		20511: begin l_1 = +14;
				 l_2 = +63; end
		46734: begin l_1 = +14;
				 l_2 = -63; end
		4127: begin l_1 = -14;
				 l_2 = +63; end
		30350: begin l_1 = -14;
				 l_2 = -63; end
		32830: begin l_1 = +14;
				 l_2 = +64; end
		34415: begin l_1 = +14;
				 l_2 = -64; end
		16446: begin l_1 = -14;
				 l_2 = +64; end
		18031: begin l_1 = -14;
				 l_2 = -64; end
		6607: begin l_1 = +14;
				 l_2 = +65; end
		9777: begin l_1 = +14;
				 l_2 = -65; end
		41084: begin l_1 = -14;
				 l_2 = +65; end
		44254: begin l_1 = -14;
				 l_2 = -65; end
		5022: begin l_1 = +14;
				 l_2 = +66; end
		11362: begin l_1 = +14;
				 l_2 = -66; end
		39499: begin l_1 = -14;
				 l_2 = +66; end
		45839: begin l_1 = -14;
				 l_2 = -66; end
		1852: begin l_1 = +14;
				 l_2 = +67; end
		14532: begin l_1 = +14;
				 l_2 = -67; end
		36329: begin l_1 = -14;
				 l_2 = +67; end
		49009: begin l_1 = -14;
				 l_2 = -67; end
		46373: begin l_1 = +14;
				 l_2 = +68; end
		20872: begin l_1 = +14;
				 l_2 = -68; end
		29989: begin l_1 = -14;
				 l_2 = +68; end
		4488: begin l_1 = -14;
				 l_2 = -68; end
		49152: begin l_1 = -15;
				 l_2 = +17; end
		1709: begin l_1 = -15;
				 l_2 = -16; end
		31059: begin l_1 = +15;
				 l_2 = +17; end
		19802: begin l_1 = -15;
				 l_2 = -17; end
		45734: begin l_1 = +15;
				 l_2 = +18; end
		37895: begin l_1 = +15;
				 l_2 = -18; end
		12966: begin l_1 = -15;
				 l_2 = +18; end
		5127: begin l_1 = -15;
				 l_2 = -18; end
		24223: begin l_1 = +15;
				 l_2 = +19; end
		8545: begin l_1 = +15;
				 l_2 = -19; end
		42316: begin l_1 = -15;
				 l_2 = +19; end
		26638: begin l_1 = -15;
				 l_2 = -19; end
		32062: begin l_1 = +15;
				 l_2 = +20; end
		706: begin l_1 = +15;
				 l_2 = -20; end
		50155: begin l_1 = -15;
				 l_2 = +20; end
		18799: begin l_1 = -15;
				 l_2 = -20; end
		47740: begin l_1 = +15;
				 l_2 = +21; end
		35889: begin l_1 = +15;
				 l_2 = -21; end
		14972: begin l_1 = -15;
				 l_2 = +21; end
		3121: begin l_1 = -15;
				 l_2 = -21; end
		28235: begin l_1 = +15;
				 l_2 = +22; end
		4533: begin l_1 = +15;
				 l_2 = -22; end
		46328: begin l_1 = -15;
				 l_2 = +22; end
		22626: begin l_1 = -15;
				 l_2 = -22; end
		40086: begin l_1 = +15;
				 l_2 = +23; end
		43543: begin l_1 = +15;
				 l_2 = -23; end
		7318: begin l_1 = -15;
				 l_2 = +23; end
		10775: begin l_1 = -15;
				 l_2 = -23; end
		12927: begin l_1 = +15;
				 l_2 = +24; end
		19841: begin l_1 = +15;
				 l_2 = -24; end
		31020: begin l_1 = -15;
				 l_2 = +24; end
		37934: begin l_1 = -15;
				 l_2 = -24; end
		9470: begin l_1 = +15;
				 l_2 = +25; end
		23298: begin l_1 = +15;
				 l_2 = -25; end
		27563: begin l_1 = -15;
				 l_2 = +25; end
		41391: begin l_1 = -15;
				 l_2 = -25; end
		2556: begin l_1 = +15;
				 l_2 = +26; end
		30212: begin l_1 = +15;
				 l_2 = -26; end
		20649: begin l_1 = -15;
				 l_2 = +26; end
		48305: begin l_1 = -15;
				 l_2 = -26; end
		39589: begin l_1 = +15;
				 l_2 = +27; end
		44040: begin l_1 = +15;
				 l_2 = -27; end
		6821: begin l_1 = -15;
				 l_2 = +27; end
		11272: begin l_1 = -15;
				 l_2 = -27; end
		11933: begin l_1 = +15;
				 l_2 = +28; end
		20835: begin l_1 = +15;
				 l_2 = -28; end
		30026: begin l_1 = -15;
				 l_2 = +28; end
		38928: begin l_1 = -15;
				 l_2 = -28; end
		7482: begin l_1 = +15;
				 l_2 = +29; end
		25286: begin l_1 = +15;
				 l_2 = -29; end
		25575: begin l_1 = -15;
				 l_2 = +29; end
		43379: begin l_1 = -15;
				 l_2 = -29; end
		49441: begin l_1 = +15;
				 l_2 = +30; end
		34188: begin l_1 = +15;
				 l_2 = -30; end
		16673: begin l_1 = -15;
				 l_2 = +30; end
		1420: begin l_1 = -15;
				 l_2 = -30; end
		31637: begin l_1 = +15;
				 l_2 = +31; end
		1131: begin l_1 = +15;
				 l_2 = -31; end
		49730: begin l_1 = -15;
				 l_2 = +31; end
		19224: begin l_1 = -15;
				 l_2 = -31; end
		46890: begin l_1 = +15;
				 l_2 = +32; end
		36739: begin l_1 = +15;
				 l_2 = -32; end
		14122: begin l_1 = -15;
				 l_2 = +32; end
		3971: begin l_1 = -15;
				 l_2 = -32; end
		26535: begin l_1 = +15;
				 l_2 = +33; end
		6233: begin l_1 = +15;
				 l_2 = -33; end
		44628: begin l_1 = -15;
				 l_2 = +33; end
		24326: begin l_1 = -15;
				 l_2 = -33; end
		36686: begin l_1 = +15;
				 l_2 = +34; end
		46943: begin l_1 = +15;
				 l_2 = -34; end
		3918: begin l_1 = -15;
				 l_2 = +34; end
		14175: begin l_1 = -15;
				 l_2 = -34; end
		6127: begin l_1 = +15;
				 l_2 = +35; end
		26641: begin l_1 = +15;
				 l_2 = -35; end
		24220: begin l_1 = -15;
				 l_2 = +35; end
		44734: begin l_1 = -15;
				 l_2 = -35; end
		46731: begin l_1 = +15;
				 l_2 = +36; end
		36898: begin l_1 = +15;
				 l_2 = -36; end
		13963: begin l_1 = -15;
				 l_2 = +36; end
		4130: begin l_1 = -15;
				 l_2 = -36; end
		26217: begin l_1 = +15;
				 l_2 = +37; end
		6551: begin l_1 = +15;
				 l_2 = -37; end
		44310: begin l_1 = -15;
				 l_2 = +37; end
		24644: begin l_1 = -15;
				 l_2 = -37; end
		36050: begin l_1 = +15;
				 l_2 = +38; end
		47579: begin l_1 = +15;
				 l_2 = -38; end
		3282: begin l_1 = -15;
				 l_2 = +38; end
		14811: begin l_1 = -15;
				 l_2 = -38; end
		4855: begin l_1 = +15;
				 l_2 = +39; end
		27913: begin l_1 = +15;
				 l_2 = -39; end
		22948: begin l_1 = -15;
				 l_2 = +39; end
		46006: begin l_1 = -15;
				 l_2 = -39; end
		44187: begin l_1 = +15;
				 l_2 = +40; end
		39442: begin l_1 = +15;
				 l_2 = -40; end
		11419: begin l_1 = -15;
				 l_2 = +40; end
		6674: begin l_1 = -15;
				 l_2 = -40; end
		21129: begin l_1 = +15;
				 l_2 = +41; end
		11639: begin l_1 = +15;
				 l_2 = -41; end
		39222: begin l_1 = -15;
				 l_2 = +41; end
		29732: begin l_1 = -15;
				 l_2 = -41; end
		25874: begin l_1 = +15;
				 l_2 = +42; end
		6894: begin l_1 = +15;
				 l_2 = -42; end
		43967: begin l_1 = -15;
				 l_2 = +42; end
		24987: begin l_1 = -15;
				 l_2 = -42; end
		35364: begin l_1 = +15;
				 l_2 = +43; end
		48265: begin l_1 = +15;
				 l_2 = -43; end
		2596: begin l_1 = -15;
				 l_2 = +43; end
		15497: begin l_1 = -15;
				 l_2 = -43; end
		3483: begin l_1 = +15;
				 l_2 = +44; end
		29285: begin l_1 = +15;
				 l_2 = -44; end
		21576: begin l_1 = -15;
				 l_2 = +44; end
		47378: begin l_1 = -15;
				 l_2 = -44; end
		41443: begin l_1 = +15;
				 l_2 = +45; end
		42186: begin l_1 = +15;
				 l_2 = -45; end
		8675: begin l_1 = -15;
				 l_2 = +45; end
		9418: begin l_1 = -15;
				 l_2 = -45; end
		15641: begin l_1 = +15;
				 l_2 = +46; end
		17127: begin l_1 = +15;
				 l_2 = -46; end
		33734: begin l_1 = -15;
				 l_2 = +46; end
		35220: begin l_1 = -15;
				 l_2 = -46; end
		14898: begin l_1 = +15;
				 l_2 = +47; end
		17870: begin l_1 = +15;
				 l_2 = -47; end
		32991: begin l_1 = -15;
				 l_2 = +47; end
		35963: begin l_1 = -15;
				 l_2 = -47; end
		13412: begin l_1 = +15;
				 l_2 = +48; end
		19356: begin l_1 = +15;
				 l_2 = -48; end
		31505: begin l_1 = -15;
				 l_2 = +48; end
		37449: begin l_1 = -15;
				 l_2 = -48; end
		10440: begin l_1 = +15;
				 l_2 = +49; end
		22328: begin l_1 = +15;
				 l_2 = -49; end
		28533: begin l_1 = -15;
				 l_2 = +49; end
		40421: begin l_1 = -15;
				 l_2 = -49; end
		4496: begin l_1 = +15;
				 l_2 = +50; end
		28272: begin l_1 = +15;
				 l_2 = -50; end
		22589: begin l_1 = -15;
				 l_2 = +50; end
		46365: begin l_1 = -15;
				 l_2 = -50; end
		43469: begin l_1 = +15;
				 l_2 = +51; end
		40160: begin l_1 = +15;
				 l_2 = -51; end
		10701: begin l_1 = -15;
				 l_2 = +51; end
		7392: begin l_1 = -15;
				 l_2 = -51; end
		19693: begin l_1 = +15;
				 l_2 = +52; end
		13075: begin l_1 = +15;
				 l_2 = -52; end
		37786: begin l_1 = -15;
				 l_2 = +52; end
		31168: begin l_1 = -15;
				 l_2 = -52; end
		23002: begin l_1 = +15;
				 l_2 = +53; end
		9766: begin l_1 = +15;
				 l_2 = -53; end
		41095: begin l_1 = -15;
				 l_2 = +53; end
		27859: begin l_1 = -15;
				 l_2 = -53; end
		29620: begin l_1 = +15;
				 l_2 = +54; end
		3148: begin l_1 = +15;
				 l_2 = -54; end
		47713: begin l_1 = -15;
				 l_2 = +54; end
		21241: begin l_1 = -15;
				 l_2 = -54; end
		42856: begin l_1 = +15;
				 l_2 = +55; end
		40773: begin l_1 = +15;
				 l_2 = -55; end
		10088: begin l_1 = -15;
				 l_2 = +55; end
		8005: begin l_1 = -15;
				 l_2 = -55; end
		18467: begin l_1 = +15;
				 l_2 = +56; end
		14301: begin l_1 = +15;
				 l_2 = -56; end
		36560: begin l_1 = -15;
				 l_2 = +56; end
		32394: begin l_1 = -15;
				 l_2 = -56; end
		20550: begin l_1 = +15;
				 l_2 = +57; end
		12218: begin l_1 = +15;
				 l_2 = -57; end
		38643: begin l_1 = -15;
				 l_2 = +57; end
		30311: begin l_1 = -15;
				 l_2 = -57; end
		24716: begin l_1 = +15;
				 l_2 = +58; end
		8052: begin l_1 = +15;
				 l_2 = -58; end
		42809: begin l_1 = -15;
				 l_2 = +58; end
		26145: begin l_1 = -15;
				 l_2 = -58; end
		33048: begin l_1 = +15;
				 l_2 = +59; end
		50581: begin l_1 = +15;
				 l_2 = -59; end
		280: begin l_1 = -15;
				 l_2 = +59; end
		17813: begin l_1 = -15;
				 l_2 = -59; end
		49712: begin l_1 = +15;
				 l_2 = +60; end
		33917: begin l_1 = +15;
				 l_2 = -60; end
		16944: begin l_1 = -15;
				 l_2 = +60; end
		1149: begin l_1 = -15;
				 l_2 = -60; end
		32179: begin l_1 = +15;
				 l_2 = +61; end
		589: begin l_1 = +15;
				 l_2 = -61; end
		50272: begin l_1 = -15;
				 l_2 = +61; end
		18682: begin l_1 = -15;
				 l_2 = -61; end
		47974: begin l_1 = +15;
				 l_2 = +62; end
		35655: begin l_1 = +15;
				 l_2 = -62; end
		15206: begin l_1 = -15;
				 l_2 = +62; end
		2887: begin l_1 = -15;
				 l_2 = -62; end
		28703: begin l_1 = +15;
				 l_2 = +63; end
		4065: begin l_1 = +15;
				 l_2 = -63; end
		46796: begin l_1 = -15;
				 l_2 = +63; end
		22158: begin l_1 = -15;
				 l_2 = -63; end
		41022: begin l_1 = +15;
				 l_2 = +64; end
		42607: begin l_1 = +15;
				 l_2 = -64; end
		8254: begin l_1 = -15;
				 l_2 = +64; end
		9839: begin l_1 = -15;
				 l_2 = -64; end
		14799: begin l_1 = +15;
				 l_2 = +65; end
		17969: begin l_1 = +15;
				 l_2 = -65; end
		32892: begin l_1 = -15;
				 l_2 = +65; end
		36062: begin l_1 = -15;
				 l_2 = -65; end
		13214: begin l_1 = +15;
				 l_2 = +66; end
		19554: begin l_1 = +15;
				 l_2 = -66; end
		31307: begin l_1 = -15;
				 l_2 = +66; end
		37647: begin l_1 = -15;
				 l_2 = -66; end
		10044: begin l_1 = +15;
				 l_2 = +67; end
		22724: begin l_1 = +15;
				 l_2 = -67; end
		28137: begin l_1 = -15;
				 l_2 = +67; end
		40817: begin l_1 = -15;
				 l_2 = -67; end
		3704: begin l_1 = +15;
				 l_2 = +68; end
		29064: begin l_1 = +15;
				 l_2 = -68; end
		21797: begin l_1 = -15;
				 l_2 = +68; end
		47157: begin l_1 = -15;
				 l_2 = -68; end
		47443: begin l_1 = -16;
				 l_2 = +18; end
		3418: begin l_1 = -16;
				 l_2 = -17; end
		11257: begin l_1 = +16;
				 l_2 = +18; end
		39604: begin l_1 = -16;
				 l_2 = -18; end
		40607: begin l_1 = +16;
				 l_2 = +19; end
		24929: begin l_1 = +16;
				 l_2 = -19; end
		25932: begin l_1 = -16;
				 l_2 = +19; end
		10254: begin l_1 = -16;
				 l_2 = -19; end
		48446: begin l_1 = +16;
				 l_2 = +20; end
		17090: begin l_1 = +16;
				 l_2 = -20; end
		33771: begin l_1 = -16;
				 l_2 = +20; end
		2415: begin l_1 = -16;
				 l_2 = -20; end
		13263: begin l_1 = +16;
				 l_2 = +21; end
		1412: begin l_1 = +16;
				 l_2 = -21; end
		49449: begin l_1 = -16;
				 l_2 = +21; end
		37598: begin l_1 = -16;
				 l_2 = -21; end
		44619: begin l_1 = +16;
				 l_2 = +22; end
		20917: begin l_1 = +16;
				 l_2 = -22; end
		29944: begin l_1 = -16;
				 l_2 = +22; end
		6242: begin l_1 = -16;
				 l_2 = -22; end
		5609: begin l_1 = +16;
				 l_2 = +23; end
		9066: begin l_1 = +16;
				 l_2 = -23; end
		41795: begin l_1 = -16;
				 l_2 = +23; end
		45252: begin l_1 = -16;
				 l_2 = -23; end
		29311: begin l_1 = +16;
				 l_2 = +24; end
		36225: begin l_1 = +16;
				 l_2 = -24; end
		14636: begin l_1 = -16;
				 l_2 = +24; end
		21550: begin l_1 = -16;
				 l_2 = -24; end
		25854: begin l_1 = +16;
				 l_2 = +25; end
		39682: begin l_1 = +16;
				 l_2 = -25; end
		11179: begin l_1 = -16;
				 l_2 = +25; end
		25007: begin l_1 = -16;
				 l_2 = -25; end
		18940: begin l_1 = +16;
				 l_2 = +26; end
		46596: begin l_1 = +16;
				 l_2 = -26; end
		4265: begin l_1 = -16;
				 l_2 = +26; end
		31921: begin l_1 = -16;
				 l_2 = -26; end
		5112: begin l_1 = +16;
				 l_2 = +27; end
		9563: begin l_1 = +16;
				 l_2 = -27; end
		41298: begin l_1 = -16;
				 l_2 = +27; end
		45749: begin l_1 = -16;
				 l_2 = -27; end
		28317: begin l_1 = +16;
				 l_2 = +28; end
		37219: begin l_1 = +16;
				 l_2 = -28; end
		13642: begin l_1 = -16;
				 l_2 = +28; end
		22544: begin l_1 = -16;
				 l_2 = -28; end
		23866: begin l_1 = +16;
				 l_2 = +29; end
		41670: begin l_1 = +16;
				 l_2 = -29; end
		9191: begin l_1 = -16;
				 l_2 = +29; end
		26995: begin l_1 = -16;
				 l_2 = -29; end
		14964: begin l_1 = +16;
				 l_2 = +30; end
		50572: begin l_1 = +16;
				 l_2 = -30; end
		289: begin l_1 = -16;
				 l_2 = +30; end
		35897: begin l_1 = -16;
				 l_2 = -30; end
		48021: begin l_1 = +16;
				 l_2 = +31; end
		17515: begin l_1 = +16;
				 l_2 = -31; end
		33346: begin l_1 = -16;
				 l_2 = +31; end
		2840: begin l_1 = -16;
				 l_2 = -31; end
		12413: begin l_1 = +16;
				 l_2 = +32; end
		2262: begin l_1 = +16;
				 l_2 = -32; end
		48599: begin l_1 = -16;
				 l_2 = +32; end
		38448: begin l_1 = -16;
				 l_2 = -32; end
		42919: begin l_1 = +16;
				 l_2 = +33; end
		22617: begin l_1 = +16;
				 l_2 = -33; end
		28244: begin l_1 = -16;
				 l_2 = +33; end
		7942: begin l_1 = -16;
				 l_2 = -33; end
		2209: begin l_1 = +16;
				 l_2 = +34; end
		12466: begin l_1 = +16;
				 l_2 = -34; end
		38395: begin l_1 = -16;
				 l_2 = +34; end
		48652: begin l_1 = -16;
				 l_2 = -34; end
		22511: begin l_1 = +16;
				 l_2 = +35; end
		43025: begin l_1 = +16;
				 l_2 = -35; end
		7836: begin l_1 = -16;
				 l_2 = +35; end
		28350: begin l_1 = -16;
				 l_2 = -35; end
		12254: begin l_1 = +16;
				 l_2 = +36; end
		2421: begin l_1 = +16;
				 l_2 = -36; end
		48440: begin l_1 = -16;
				 l_2 = +36; end
		38607: begin l_1 = -16;
				 l_2 = -36; end
		42601: begin l_1 = +16;
				 l_2 = +37; end
		22935: begin l_1 = +16;
				 l_2 = -37; end
		27926: begin l_1 = -16;
				 l_2 = +37; end
		8260: begin l_1 = -16;
				 l_2 = -37; end
		1573: begin l_1 = +16;
				 l_2 = +38; end
		13102: begin l_1 = +16;
				 l_2 = -38; end
		37759: begin l_1 = -16;
				 l_2 = +38; end
		49288: begin l_1 = -16;
				 l_2 = -38; end
		21239: begin l_1 = +16;
				 l_2 = +39; end
		44297: begin l_1 = +16;
				 l_2 = -39; end
		6564: begin l_1 = -16;
				 l_2 = +39; end
		29622: begin l_1 = -16;
				 l_2 = -39; end
		9710: begin l_1 = +16;
				 l_2 = +40; end
		4965: begin l_1 = +16;
				 l_2 = -40; end
		45896: begin l_1 = -16;
				 l_2 = +40; end
		41151: begin l_1 = -16;
				 l_2 = -40; end
		37513: begin l_1 = +16;
				 l_2 = +41; end
		28023: begin l_1 = +16;
				 l_2 = -41; end
		22838: begin l_1 = -16;
				 l_2 = +41; end
		13348: begin l_1 = -16;
				 l_2 = -41; end
		42258: begin l_1 = +16;
				 l_2 = +42; end
		23278: begin l_1 = +16;
				 l_2 = -42; end
		27583: begin l_1 = -16;
				 l_2 = +42; end
		8603: begin l_1 = -16;
				 l_2 = -42; end
		887: begin l_1 = +16;
				 l_2 = +43; end
		13788: begin l_1 = +16;
				 l_2 = -43; end
		37073: begin l_1 = -16;
				 l_2 = +43; end
		49974: begin l_1 = -16;
				 l_2 = -43; end
		19867: begin l_1 = +16;
				 l_2 = +44; end
		45669: begin l_1 = +16;
				 l_2 = -44; end
		5192: begin l_1 = -16;
				 l_2 = +44; end
		30994: begin l_1 = -16;
				 l_2 = -44; end
		6966: begin l_1 = +16;
				 l_2 = +45; end
		7709: begin l_1 = +16;
				 l_2 = -45; end
		43152: begin l_1 = -16;
				 l_2 = +45; end
		43895: begin l_1 = -16;
				 l_2 = -45; end
		32025: begin l_1 = +16;
				 l_2 = +46; end
		33511: begin l_1 = +16;
				 l_2 = -46; end
		17350: begin l_1 = -16;
				 l_2 = +46; end
		18836: begin l_1 = -16;
				 l_2 = -46; end
		31282: begin l_1 = +16;
				 l_2 = +47; end
		34254: begin l_1 = +16;
				 l_2 = -47; end
		16607: begin l_1 = -16;
				 l_2 = +47; end
		19579: begin l_1 = -16;
				 l_2 = -47; end
		29796: begin l_1 = +16;
				 l_2 = +48; end
		35740: begin l_1 = +16;
				 l_2 = -48; end
		15121: begin l_1 = -16;
				 l_2 = +48; end
		21065: begin l_1 = -16;
				 l_2 = -48; end
		26824: begin l_1 = +16;
				 l_2 = +49; end
		38712: begin l_1 = +16;
				 l_2 = -49; end
		12149: begin l_1 = -16;
				 l_2 = +49; end
		24037: begin l_1 = -16;
				 l_2 = -49; end
		20880: begin l_1 = +16;
				 l_2 = +50; end
		44656: begin l_1 = +16;
				 l_2 = -50; end
		6205: begin l_1 = -16;
				 l_2 = +50; end
		29981: begin l_1 = -16;
				 l_2 = -50; end
		8992: begin l_1 = +16;
				 l_2 = +51; end
		5683: begin l_1 = +16;
				 l_2 = -51; end
		45178: begin l_1 = -16;
				 l_2 = +51; end
		41869: begin l_1 = -16;
				 l_2 = -51; end
		36077: begin l_1 = +16;
				 l_2 = +52; end
		29459: begin l_1 = +16;
				 l_2 = -52; end
		21402: begin l_1 = -16;
				 l_2 = +52; end
		14784: begin l_1 = -16;
				 l_2 = -52; end
		39386: begin l_1 = +16;
				 l_2 = +53; end
		26150: begin l_1 = +16;
				 l_2 = -53; end
		24711: begin l_1 = -16;
				 l_2 = +53; end
		11475: begin l_1 = -16;
				 l_2 = -53; end
		46004: begin l_1 = +16;
				 l_2 = +54; end
		19532: begin l_1 = +16;
				 l_2 = -54; end
		31329: begin l_1 = -16;
				 l_2 = +54; end
		4857: begin l_1 = -16;
				 l_2 = -54; end
		8379: begin l_1 = +16;
				 l_2 = +55; end
		6296: begin l_1 = +16;
				 l_2 = -55; end
		44565: begin l_1 = -16;
				 l_2 = +55; end
		42482: begin l_1 = -16;
				 l_2 = -55; end
		34851: begin l_1 = +16;
				 l_2 = +56; end
		30685: begin l_1 = +16;
				 l_2 = -56; end
		20176: begin l_1 = -16;
				 l_2 = +56; end
		16010: begin l_1 = -16;
				 l_2 = -56; end
		36934: begin l_1 = +16;
				 l_2 = +57; end
		28602: begin l_1 = +16;
				 l_2 = -57; end
		22259: begin l_1 = -16;
				 l_2 = +57; end
		13927: begin l_1 = -16;
				 l_2 = -57; end
		41100: begin l_1 = +16;
				 l_2 = +58; end
		24436: begin l_1 = +16;
				 l_2 = -58; end
		26425: begin l_1 = -16;
				 l_2 = +58; end
		9761: begin l_1 = -16;
				 l_2 = -58; end
		49432: begin l_1 = +16;
				 l_2 = +59; end
		16104: begin l_1 = +16;
				 l_2 = -59; end
		34757: begin l_1 = -16;
				 l_2 = +59; end
		1429: begin l_1 = -16;
				 l_2 = -59; end
		15235: begin l_1 = +16;
				 l_2 = +60; end
		50301: begin l_1 = +16;
				 l_2 = -60; end
		560: begin l_1 = -16;
				 l_2 = +60; end
		35626: begin l_1 = -16;
				 l_2 = -60; end
		48563: begin l_1 = +16;
				 l_2 = +61; end
		16973: begin l_1 = +16;
				 l_2 = -61; end
		33888: begin l_1 = -16;
				 l_2 = +61; end
		2298: begin l_1 = -16;
				 l_2 = -61; end
		13497: begin l_1 = +16;
				 l_2 = +62; end
		1178: begin l_1 = +16;
				 l_2 = -62; end
		49683: begin l_1 = -16;
				 l_2 = +62; end
		37364: begin l_1 = -16;
				 l_2 = -62; end
		45087: begin l_1 = +16;
				 l_2 = +63; end
		20449: begin l_1 = +16;
				 l_2 = -63; end
		30412: begin l_1 = -16;
				 l_2 = +63; end
		5774: begin l_1 = -16;
				 l_2 = -63; end
		6545: begin l_1 = +16;
				 l_2 = +64; end
		8130: begin l_1 = +16;
				 l_2 = -64; end
		42731: begin l_1 = -16;
				 l_2 = +64; end
		44316: begin l_1 = -16;
				 l_2 = -64; end
		31183: begin l_1 = +16;
				 l_2 = +65; end
		34353: begin l_1 = +16;
				 l_2 = -65; end
		16508: begin l_1 = -16;
				 l_2 = +65; end
		19678: begin l_1 = -16;
				 l_2 = -65; end
		29598: begin l_1 = +16;
				 l_2 = +66; end
		35938: begin l_1 = +16;
				 l_2 = -66; end
		14923: begin l_1 = -16;
				 l_2 = +66; end
		21263: begin l_1 = -16;
				 l_2 = -66; end
		26428: begin l_1 = +16;
				 l_2 = +67; end
		39108: begin l_1 = +16;
				 l_2 = -67; end
		11753: begin l_1 = -16;
				 l_2 = +67; end
		24433: begin l_1 = -16;
				 l_2 = -67; end
		20088: begin l_1 = +16;
				 l_2 = +68; end
		45448: begin l_1 = +16;
				 l_2 = -68; end
		5413: begin l_1 = -16;
				 l_2 = +68; end
		30773: begin l_1 = -16;
				 l_2 = -68; end
		44025: begin l_1 = -17;
				 l_2 = +19; end
		6836: begin l_1 = -17;
				 l_2 = -18; end
		22514: begin l_1 = +17;
				 l_2 = +19; end
		28347: begin l_1 = -17;
				 l_2 = -19; end
		30353: begin l_1 = +17;
				 l_2 = +20; end
		49858: begin l_1 = +17;
				 l_2 = -20; end
		1003: begin l_1 = -17;
				 l_2 = +20; end
		20508: begin l_1 = -17;
				 l_2 = -20; end
		46031: begin l_1 = +17;
				 l_2 = +21; end
		34180: begin l_1 = +17;
				 l_2 = -21; end
		16681: begin l_1 = -17;
				 l_2 = +21; end
		4830: begin l_1 = -17;
				 l_2 = -21; end
		26526: begin l_1 = +17;
				 l_2 = +22; end
		2824: begin l_1 = +17;
				 l_2 = -22; end
		48037: begin l_1 = -17;
				 l_2 = +22; end
		24335: begin l_1 = -17;
				 l_2 = -22; end
		38377: begin l_1 = +17;
				 l_2 = +23; end
		41834: begin l_1 = +17;
				 l_2 = -23; end
		9027: begin l_1 = -17;
				 l_2 = +23; end
		12484: begin l_1 = -17;
				 l_2 = -23; end
		11218: begin l_1 = +17;
				 l_2 = +24; end
		18132: begin l_1 = +17;
				 l_2 = -24; end
		32729: begin l_1 = -17;
				 l_2 = +24; end
		39643: begin l_1 = -17;
				 l_2 = -24; end
		7761: begin l_1 = +17;
				 l_2 = +25; end
		21589: begin l_1 = +17;
				 l_2 = -25; end
		29272: begin l_1 = -17;
				 l_2 = +25; end
		43100: begin l_1 = -17;
				 l_2 = -25; end
		847: begin l_1 = +17;
				 l_2 = +26; end
		28503: begin l_1 = +17;
				 l_2 = -26; end
		22358: begin l_1 = -17;
				 l_2 = +26; end
		50014: begin l_1 = -17;
				 l_2 = -26; end
		37880: begin l_1 = +17;
				 l_2 = +27; end
		42331: begin l_1 = +17;
				 l_2 = -27; end
		8530: begin l_1 = -17;
				 l_2 = +27; end
		12981: begin l_1 = -17;
				 l_2 = -27; end
		10224: begin l_1 = +17;
				 l_2 = +28; end
		19126: begin l_1 = +17;
				 l_2 = -28; end
		31735: begin l_1 = -17;
				 l_2 = +28; end
		40637: begin l_1 = -17;
				 l_2 = -28; end
		5773: begin l_1 = +17;
				 l_2 = +29; end
		23577: begin l_1 = +17;
				 l_2 = -29; end
		27284: begin l_1 = -17;
				 l_2 = +29; end
		45088: begin l_1 = -17;
				 l_2 = -29; end
		47732: begin l_1 = +17;
				 l_2 = +30; end
		32479: begin l_1 = +17;
				 l_2 = -30; end
		18382: begin l_1 = -17;
				 l_2 = +30; end
		3129: begin l_1 = -17;
				 l_2 = -30; end
		29928: begin l_1 = +17;
				 l_2 = +31; end
		50283: begin l_1 = +17;
				 l_2 = -31; end
		578: begin l_1 = -17;
				 l_2 = +31; end
		20933: begin l_1 = -17;
				 l_2 = -31; end
		45181: begin l_1 = +17;
				 l_2 = +32; end
		35030: begin l_1 = +17;
				 l_2 = -32; end
		15831: begin l_1 = -17;
				 l_2 = +32; end
		5680: begin l_1 = -17;
				 l_2 = -32; end
		24826: begin l_1 = +17;
				 l_2 = +33; end
		4524: begin l_1 = +17;
				 l_2 = -33; end
		46337: begin l_1 = -17;
				 l_2 = +33; end
		26035: begin l_1 = -17;
				 l_2 = -33; end
		34977: begin l_1 = +17;
				 l_2 = +34; end
		45234: begin l_1 = +17;
				 l_2 = -34; end
		5627: begin l_1 = -17;
				 l_2 = +34; end
		15884: begin l_1 = -17;
				 l_2 = -34; end
		4418: begin l_1 = +17;
				 l_2 = +35; end
		24932: begin l_1 = +17;
				 l_2 = -35; end
		25929: begin l_1 = -17;
				 l_2 = +35; end
		46443: begin l_1 = -17;
				 l_2 = -35; end
		45022: begin l_1 = +17;
				 l_2 = +36; end
		35189: begin l_1 = +17;
				 l_2 = -36; end
		15672: begin l_1 = -17;
				 l_2 = +36; end
		5839: begin l_1 = -17;
				 l_2 = -36; end
		24508: begin l_1 = +17;
				 l_2 = +37; end
		4842: begin l_1 = +17;
				 l_2 = -37; end
		46019: begin l_1 = -17;
				 l_2 = +37; end
		26353: begin l_1 = -17;
				 l_2 = -37; end
		34341: begin l_1 = +17;
				 l_2 = +38; end
		45870: begin l_1 = +17;
				 l_2 = -38; end
		4991: begin l_1 = -17;
				 l_2 = +38; end
		16520: begin l_1 = -17;
				 l_2 = -38; end
		3146: begin l_1 = +17;
				 l_2 = +39; end
		26204: begin l_1 = +17;
				 l_2 = -39; end
		24657: begin l_1 = -17;
				 l_2 = +39; end
		47715: begin l_1 = -17;
				 l_2 = -39; end
		42478: begin l_1 = +17;
				 l_2 = +40; end
		37733: begin l_1 = +17;
				 l_2 = -40; end
		13128: begin l_1 = -17;
				 l_2 = +40; end
		8383: begin l_1 = -17;
				 l_2 = -40; end
		19420: begin l_1 = +17;
				 l_2 = +41; end
		9930: begin l_1 = +17;
				 l_2 = -41; end
		40931: begin l_1 = -17;
				 l_2 = +41; end
		31441: begin l_1 = -17;
				 l_2 = -41; end
		24165: begin l_1 = +17;
				 l_2 = +42; end
		5185: begin l_1 = +17;
				 l_2 = -42; end
		45676: begin l_1 = -17;
				 l_2 = +42; end
		26696: begin l_1 = -17;
				 l_2 = -42; end
		33655: begin l_1 = +17;
				 l_2 = +43; end
		46556: begin l_1 = +17;
				 l_2 = -43; end
		4305: begin l_1 = -17;
				 l_2 = +43; end
		17206: begin l_1 = -17;
				 l_2 = -43; end
		1774: begin l_1 = +17;
				 l_2 = +44; end
		27576: begin l_1 = +17;
				 l_2 = -44; end
		23285: begin l_1 = -17;
				 l_2 = +44; end
		49087: begin l_1 = -17;
				 l_2 = -44; end
		39734: begin l_1 = +17;
				 l_2 = +45; end
		40477: begin l_1 = +17;
				 l_2 = -45; end
		10384: begin l_1 = -17;
				 l_2 = +45; end
		11127: begin l_1 = -17;
				 l_2 = -45; end
		13932: begin l_1 = +17;
				 l_2 = +46; end
		15418: begin l_1 = +17;
				 l_2 = -46; end
		35443: begin l_1 = -17;
				 l_2 = +46; end
		36929: begin l_1 = -17;
				 l_2 = -46; end
		13189: begin l_1 = +17;
				 l_2 = +47; end
		16161: begin l_1 = +17;
				 l_2 = -47; end
		34700: begin l_1 = -17;
				 l_2 = +47; end
		37672: begin l_1 = -17;
				 l_2 = -47; end
		11703: begin l_1 = +17;
				 l_2 = +48; end
		17647: begin l_1 = +17;
				 l_2 = -48; end
		33214: begin l_1 = -17;
				 l_2 = +48; end
		39158: begin l_1 = -17;
				 l_2 = -48; end
		8731: begin l_1 = +17;
				 l_2 = +49; end
		20619: begin l_1 = +17;
				 l_2 = -49; end
		30242: begin l_1 = -17;
				 l_2 = +49; end
		42130: begin l_1 = -17;
				 l_2 = -49; end
		2787: begin l_1 = +17;
				 l_2 = +50; end
		26563: begin l_1 = +17;
				 l_2 = -50; end
		24298: begin l_1 = -17;
				 l_2 = +50; end
		48074: begin l_1 = -17;
				 l_2 = -50; end
		41760: begin l_1 = +17;
				 l_2 = +51; end
		38451: begin l_1 = +17;
				 l_2 = -51; end
		12410: begin l_1 = -17;
				 l_2 = +51; end
		9101: begin l_1 = -17;
				 l_2 = -51; end
		17984: begin l_1 = +17;
				 l_2 = +52; end
		11366: begin l_1 = +17;
				 l_2 = -52; end
		39495: begin l_1 = -17;
				 l_2 = +52; end
		32877: begin l_1 = -17;
				 l_2 = -52; end
		21293: begin l_1 = +17;
				 l_2 = +53; end
		8057: begin l_1 = +17;
				 l_2 = -53; end
		42804: begin l_1 = -17;
				 l_2 = +53; end
		29568: begin l_1 = -17;
				 l_2 = -53; end
		27911: begin l_1 = +17;
				 l_2 = +54; end
		1439: begin l_1 = +17;
				 l_2 = -54; end
		49422: begin l_1 = -17;
				 l_2 = +54; end
		22950: begin l_1 = -17;
				 l_2 = -54; end
		41147: begin l_1 = +17;
				 l_2 = +55; end
		39064: begin l_1 = +17;
				 l_2 = -55; end
		11797: begin l_1 = -17;
				 l_2 = +55; end
		9714: begin l_1 = -17;
				 l_2 = -55; end
		16758: begin l_1 = +17;
				 l_2 = +56; end
		12592: begin l_1 = +17;
				 l_2 = -56; end
		38269: begin l_1 = -17;
				 l_2 = +56; end
		34103: begin l_1 = -17;
				 l_2 = -56; end
		18841: begin l_1 = +17;
				 l_2 = +57; end
		10509: begin l_1 = +17;
				 l_2 = -57; end
		40352: begin l_1 = -17;
				 l_2 = +57; end
		32020: begin l_1 = -17;
				 l_2 = -57; end
		23007: begin l_1 = +17;
				 l_2 = +58; end
		6343: begin l_1 = +17;
				 l_2 = -58; end
		44518: begin l_1 = -17;
				 l_2 = +58; end
		27854: begin l_1 = -17;
				 l_2 = -58; end
		31339: begin l_1 = +17;
				 l_2 = +59; end
		48872: begin l_1 = +17;
				 l_2 = -59; end
		1989: begin l_1 = -17;
				 l_2 = +59; end
		19522: begin l_1 = -17;
				 l_2 = -59; end
		48003: begin l_1 = +17;
				 l_2 = +60; end
		32208: begin l_1 = +17;
				 l_2 = -60; end
		18653: begin l_1 = -17;
				 l_2 = +60; end
		2858: begin l_1 = -17;
				 l_2 = -60; end
		30470: begin l_1 = +17;
				 l_2 = +61; end
		49741: begin l_1 = +17;
				 l_2 = -61; end
		1120: begin l_1 = -17;
				 l_2 = +61; end
		20391: begin l_1 = -17;
				 l_2 = -61; end
		46265: begin l_1 = +17;
				 l_2 = +62; end
		33946: begin l_1 = +17;
				 l_2 = -62; end
		16915: begin l_1 = -17;
				 l_2 = +62; end
		4596: begin l_1 = -17;
				 l_2 = -62; end
		26994: begin l_1 = +17;
				 l_2 = +63; end
		2356: begin l_1 = +17;
				 l_2 = -63; end
		48505: begin l_1 = -17;
				 l_2 = +63; end
		23867: begin l_1 = -17;
				 l_2 = -63; end
		39313: begin l_1 = +17;
				 l_2 = +64; end
		40898: begin l_1 = +17;
				 l_2 = -64; end
		9963: begin l_1 = -17;
				 l_2 = +64; end
		11548: begin l_1 = -17;
				 l_2 = -64; end
		13090: begin l_1 = +17;
				 l_2 = +65; end
		16260: begin l_1 = +17;
				 l_2 = -65; end
		34601: begin l_1 = -17;
				 l_2 = +65; end
		37771: begin l_1 = -17;
				 l_2 = -65; end
		11505: begin l_1 = +17;
				 l_2 = +66; end
		17845: begin l_1 = +17;
				 l_2 = -66; end
		33016: begin l_1 = -17;
				 l_2 = +66; end
		39356: begin l_1 = -17;
				 l_2 = -66; end
		8335: begin l_1 = +17;
				 l_2 = +67; end
		21015: begin l_1 = +17;
				 l_2 = -67; end
		29846: begin l_1 = -17;
				 l_2 = +67; end
		42526: begin l_1 = -17;
				 l_2 = -67; end
		1995: begin l_1 = +17;
				 l_2 = +68; end
		27355: begin l_1 = +17;
				 l_2 = -68; end
		23506: begin l_1 = -17;
				 l_2 = +68; end
		48866: begin l_1 = -17;
				 l_2 = -68; end
		37189: begin l_1 = -18;
				 l_2 = +20; end
		13672: begin l_1 = -18;
				 l_2 = -19; end
		45028: begin l_1 = +18;
				 l_2 = +20; end
		5833: begin l_1 = -18;
				 l_2 = -20; end
		9845: begin l_1 = +18;
				 l_2 = +21; end
		48855: begin l_1 = +18;
				 l_2 = -21; end
		2006: begin l_1 = -18;
				 l_2 = +21; end
		41016: begin l_1 = -18;
				 l_2 = -21; end
		41201: begin l_1 = +18;
				 l_2 = +22; end
		17499: begin l_1 = +18;
				 l_2 = -22; end
		33362: begin l_1 = -18;
				 l_2 = +22; end
		9660: begin l_1 = -18;
				 l_2 = -22; end
		2191: begin l_1 = +18;
				 l_2 = +23; end
		5648: begin l_1 = +18;
				 l_2 = -23; end
		45213: begin l_1 = -18;
				 l_2 = +23; end
		48670: begin l_1 = -18;
				 l_2 = -23; end
		25893: begin l_1 = +18;
				 l_2 = +24; end
		32807: begin l_1 = +18;
				 l_2 = -24; end
		18054: begin l_1 = -18;
				 l_2 = +24; end
		24968: begin l_1 = -18;
				 l_2 = -24; end
		22436: begin l_1 = +18;
				 l_2 = +25; end
		36264: begin l_1 = +18;
				 l_2 = -25; end
		14597: begin l_1 = -18;
				 l_2 = +25; end
		28425: begin l_1 = -18;
				 l_2 = -25; end
		15522: begin l_1 = +18;
				 l_2 = +26; end
		43178: begin l_1 = +18;
				 l_2 = -26; end
		7683: begin l_1 = -18;
				 l_2 = +26; end
		35339: begin l_1 = -18;
				 l_2 = -26; end
		1694: begin l_1 = +18;
				 l_2 = +27; end
		6145: begin l_1 = +18;
				 l_2 = -27; end
		44716: begin l_1 = -18;
				 l_2 = +27; end
		49167: begin l_1 = -18;
				 l_2 = -27; end
		24899: begin l_1 = +18;
				 l_2 = +28; end
		33801: begin l_1 = +18;
				 l_2 = -28; end
		17060: begin l_1 = -18;
				 l_2 = +28; end
		25962: begin l_1 = -18;
				 l_2 = -28; end
		20448: begin l_1 = +18;
				 l_2 = +29; end
		38252: begin l_1 = +18;
				 l_2 = -29; end
		12609: begin l_1 = -18;
				 l_2 = +29; end
		30413: begin l_1 = -18;
				 l_2 = -29; end
		11546: begin l_1 = +18;
				 l_2 = +30; end
		47154: begin l_1 = +18;
				 l_2 = -30; end
		3707: begin l_1 = -18;
				 l_2 = +30; end
		39315: begin l_1 = -18;
				 l_2 = -30; end
		44603: begin l_1 = +18;
				 l_2 = +31; end
		14097: begin l_1 = +18;
				 l_2 = -31; end
		36764: begin l_1 = -18;
				 l_2 = +31; end
		6258: begin l_1 = -18;
				 l_2 = -31; end
		8995: begin l_1 = +18;
				 l_2 = +32; end
		49705: begin l_1 = +18;
				 l_2 = -32; end
		1156: begin l_1 = -18;
				 l_2 = +32; end
		41866: begin l_1 = -18;
				 l_2 = -32; end
		39501: begin l_1 = +18;
				 l_2 = +33; end
		19199: begin l_1 = +18;
				 l_2 = -33; end
		31662: begin l_1 = -18;
				 l_2 = +33; end
		11360: begin l_1 = -18;
				 l_2 = -33; end
		49652: begin l_1 = +18;
				 l_2 = +34; end
		9048: begin l_1 = +18;
				 l_2 = -34; end
		41813: begin l_1 = -18;
				 l_2 = +34; end
		1209: begin l_1 = -18;
				 l_2 = -34; end
		19093: begin l_1 = +18;
				 l_2 = +35; end
		39607: begin l_1 = +18;
				 l_2 = -35; end
		11254: begin l_1 = -18;
				 l_2 = +35; end
		31768: begin l_1 = -18;
				 l_2 = -35; end
		8836: begin l_1 = +18;
				 l_2 = +36; end
		49864: begin l_1 = +18;
				 l_2 = -36; end
		997: begin l_1 = -18;
				 l_2 = +36; end
		42025: begin l_1 = -18;
				 l_2 = -36; end
		39183: begin l_1 = +18;
				 l_2 = +37; end
		19517: begin l_1 = +18;
				 l_2 = -37; end
		31344: begin l_1 = -18;
				 l_2 = +37; end
		11678: begin l_1 = -18;
				 l_2 = -37; end
		49016: begin l_1 = +18;
				 l_2 = +38; end
		9684: begin l_1 = +18;
				 l_2 = -38; end
		41177: begin l_1 = -18;
				 l_2 = +38; end
		1845: begin l_1 = -18;
				 l_2 = -38; end
		17821: begin l_1 = +18;
				 l_2 = +39; end
		40879: begin l_1 = +18;
				 l_2 = -39; end
		9982: begin l_1 = -18;
				 l_2 = +39; end
		33040: begin l_1 = -18;
				 l_2 = -39; end
		6292: begin l_1 = +18;
				 l_2 = +40; end
		1547: begin l_1 = +18;
				 l_2 = -40; end
		49314: begin l_1 = -18;
				 l_2 = +40; end
		44569: begin l_1 = -18;
				 l_2 = -40; end
		34095: begin l_1 = +18;
				 l_2 = +41; end
		24605: begin l_1 = +18;
				 l_2 = -41; end
		26256: begin l_1 = -18;
				 l_2 = +41; end
		16766: begin l_1 = -18;
				 l_2 = -41; end
		38840: begin l_1 = +18;
				 l_2 = +42; end
		19860: begin l_1 = +18;
				 l_2 = -42; end
		31001: begin l_1 = -18;
				 l_2 = +42; end
		12021: begin l_1 = -18;
				 l_2 = -42; end
		48330: begin l_1 = +18;
				 l_2 = +43; end
		10370: begin l_1 = +18;
				 l_2 = -43; end
		40491: begin l_1 = -18;
				 l_2 = +43; end
		2531: begin l_1 = -18;
				 l_2 = -43; end
		16449: begin l_1 = +18;
				 l_2 = +44; end
		42251: begin l_1 = +18;
				 l_2 = -44; end
		8610: begin l_1 = -18;
				 l_2 = +44; end
		34412: begin l_1 = -18;
				 l_2 = -44; end
		3548: begin l_1 = +18;
				 l_2 = +45; end
		4291: begin l_1 = +18;
				 l_2 = -45; end
		46570: begin l_1 = -18;
				 l_2 = +45; end
		47313: begin l_1 = -18;
				 l_2 = -45; end
		28607: begin l_1 = +18;
				 l_2 = +46; end
		30093: begin l_1 = +18;
				 l_2 = -46; end
		20768: begin l_1 = -18;
				 l_2 = +46; end
		22254: begin l_1 = -18;
				 l_2 = -46; end
		27864: begin l_1 = +18;
				 l_2 = +47; end
		30836: begin l_1 = +18;
				 l_2 = -47; end
		20025: begin l_1 = -18;
				 l_2 = +47; end
		22997: begin l_1 = -18;
				 l_2 = -47; end
		26378: begin l_1 = +18;
				 l_2 = +48; end
		32322: begin l_1 = +18;
				 l_2 = -48; end
		18539: begin l_1 = -18;
				 l_2 = +48; end
		24483: begin l_1 = -18;
				 l_2 = -48; end
		23406: begin l_1 = +18;
				 l_2 = +49; end
		35294: begin l_1 = +18;
				 l_2 = -49; end
		15567: begin l_1 = -18;
				 l_2 = +49; end
		27455: begin l_1 = -18;
				 l_2 = -49; end
		17462: begin l_1 = +18;
				 l_2 = +50; end
		41238: begin l_1 = +18;
				 l_2 = -50; end
		9623: begin l_1 = -18;
				 l_2 = +50; end
		33399: begin l_1 = -18;
				 l_2 = -50; end
		5574: begin l_1 = +18;
				 l_2 = +51; end
		2265: begin l_1 = +18;
				 l_2 = -51; end
		48596: begin l_1 = -18;
				 l_2 = +51; end
		45287: begin l_1 = -18;
				 l_2 = -51; end
		32659: begin l_1 = +18;
				 l_2 = +52; end
		26041: begin l_1 = +18;
				 l_2 = -52; end
		24820: begin l_1 = -18;
				 l_2 = +52; end
		18202: begin l_1 = -18;
				 l_2 = -52; end
		35968: begin l_1 = +18;
				 l_2 = +53; end
		22732: begin l_1 = +18;
				 l_2 = -53; end
		28129: begin l_1 = -18;
				 l_2 = +53; end
		14893: begin l_1 = -18;
				 l_2 = -53; end
		42586: begin l_1 = +18;
				 l_2 = +54; end
		16114: begin l_1 = +18;
				 l_2 = -54; end
		34747: begin l_1 = -18;
				 l_2 = +54; end
		8275: begin l_1 = -18;
				 l_2 = -54; end
		4961: begin l_1 = +18;
				 l_2 = +55; end
		2878: begin l_1 = +18;
				 l_2 = -55; end
		47983: begin l_1 = -18;
				 l_2 = +55; end
		45900: begin l_1 = -18;
				 l_2 = -55; end
		31433: begin l_1 = +18;
				 l_2 = +56; end
		27267: begin l_1 = +18;
				 l_2 = -56; end
		23594: begin l_1 = -18;
				 l_2 = +56; end
		19428: begin l_1 = -18;
				 l_2 = -56; end
		33516: begin l_1 = +18;
				 l_2 = +57; end
		25184: begin l_1 = +18;
				 l_2 = -57; end
		25677: begin l_1 = -18;
				 l_2 = +57; end
		17345: begin l_1 = -18;
				 l_2 = -57; end
		37682: begin l_1 = +18;
				 l_2 = +58; end
		21018: begin l_1 = +18;
				 l_2 = -58; end
		29843: begin l_1 = -18;
				 l_2 = +58; end
		13179: begin l_1 = -18;
				 l_2 = -58; end
		46014: begin l_1 = +18;
				 l_2 = +59; end
		12686: begin l_1 = +18;
				 l_2 = -59; end
		38175: begin l_1 = -18;
				 l_2 = +59; end
		4847: begin l_1 = -18;
				 l_2 = -59; end
		11817: begin l_1 = +18;
				 l_2 = +60; end
		46883: begin l_1 = +18;
				 l_2 = -60; end
		3978: begin l_1 = -18;
				 l_2 = +60; end
		39044: begin l_1 = -18;
				 l_2 = -60; end
		45145: begin l_1 = +18;
				 l_2 = +61; end
		13555: begin l_1 = +18;
				 l_2 = -61; end
		37306: begin l_1 = -18;
				 l_2 = +61; end
		5716: begin l_1 = -18;
				 l_2 = -61; end
		10079: begin l_1 = +18;
				 l_2 = +62; end
		48621: begin l_1 = +18;
				 l_2 = -62; end
		2240: begin l_1 = -18;
				 l_2 = +62; end
		40782: begin l_1 = -18;
				 l_2 = -62; end
		41669: begin l_1 = +18;
				 l_2 = +63; end
		17031: begin l_1 = +18;
				 l_2 = -63; end
		33830: begin l_1 = -18;
				 l_2 = +63; end
		9192: begin l_1 = -18;
				 l_2 = -63; end
		3127: begin l_1 = +18;
				 l_2 = +64; end
		4712: begin l_1 = +18;
				 l_2 = -64; end
		46149: begin l_1 = -18;
				 l_2 = +64; end
		47734: begin l_1 = -18;
				 l_2 = -64; end
		27765: begin l_1 = +18;
				 l_2 = +65; end
		30935: begin l_1 = +18;
				 l_2 = -65; end
		19926: begin l_1 = -18;
				 l_2 = +65; end
		23096: begin l_1 = -18;
				 l_2 = -65; end
		26180: begin l_1 = +18;
				 l_2 = +66; end
		32520: begin l_1 = +18;
				 l_2 = -66; end
		18341: begin l_1 = -18;
				 l_2 = +66; end
		24681: begin l_1 = -18;
				 l_2 = -66; end
		23010: begin l_1 = +18;
				 l_2 = +67; end
		35690: begin l_1 = +18;
				 l_2 = -67; end
		15171: begin l_1 = -18;
				 l_2 = +67; end
		27851: begin l_1 = -18;
				 l_2 = -67; end
		16670: begin l_1 = +18;
				 l_2 = +68; end
		42030: begin l_1 = +18;
				 l_2 = -68; end
		8831: begin l_1 = -18;
				 l_2 = +68; end
		34191: begin l_1 = -18;
				 l_2 = -68; end
		23517: begin l_1 = -19;
				 l_2 = +21; end
		27344: begin l_1 = -19;
				 l_2 = -20; end
		39195: begin l_1 = +19;
				 l_2 = +21; end
		11666: begin l_1 = -19;
				 l_2 = -21; end
		19690: begin l_1 = +19;
				 l_2 = +22; end
		46849: begin l_1 = +19;
				 l_2 = -22; end
		4012: begin l_1 = -19;
				 l_2 = +22; end
		31171: begin l_1 = -19;
				 l_2 = -22; end
		31541: begin l_1 = +19;
				 l_2 = +23; end
		34998: begin l_1 = +19;
				 l_2 = -23; end
		15863: begin l_1 = -19;
				 l_2 = +23; end
		19320: begin l_1 = -19;
				 l_2 = -23; end
		4382: begin l_1 = +19;
				 l_2 = +24; end
		11296: begin l_1 = +19;
				 l_2 = -24; end
		39565: begin l_1 = -19;
				 l_2 = +24; end
		46479: begin l_1 = -19;
				 l_2 = -24; end
		925: begin l_1 = +19;
				 l_2 = +25; end
		14753: begin l_1 = +19;
				 l_2 = -25; end
		36108: begin l_1 = -19;
				 l_2 = +25; end
		49936: begin l_1 = -19;
				 l_2 = -25; end
		44872: begin l_1 = +19;
				 l_2 = +26; end
		21667: begin l_1 = +19;
				 l_2 = -26; end
		29194: begin l_1 = -19;
				 l_2 = +26; end
		5989: begin l_1 = -19;
				 l_2 = -26; end
		31044: begin l_1 = +19;
				 l_2 = +27; end
		35495: begin l_1 = +19;
				 l_2 = -27; end
		15366: begin l_1 = -19;
				 l_2 = +27; end
		19817: begin l_1 = -19;
				 l_2 = -27; end
		3388: begin l_1 = +19;
				 l_2 = +28; end
		12290: begin l_1 = +19;
				 l_2 = -28; end
		38571: begin l_1 = -19;
				 l_2 = +28; end
		47473: begin l_1 = -19;
				 l_2 = -28; end
		49798: begin l_1 = +19;
				 l_2 = +29; end
		16741: begin l_1 = +19;
				 l_2 = -29; end
		34120: begin l_1 = -19;
				 l_2 = +29; end
		1063: begin l_1 = -19;
				 l_2 = -29; end
		40896: begin l_1 = +19;
				 l_2 = +30; end
		25643: begin l_1 = +19;
				 l_2 = -30; end
		25218: begin l_1 = -19;
				 l_2 = +30; end
		9965: begin l_1 = -19;
				 l_2 = -30; end
		23092: begin l_1 = +19;
				 l_2 = +31; end
		43447: begin l_1 = +19;
				 l_2 = -31; end
		7414: begin l_1 = -19;
				 l_2 = +31; end
		27769: begin l_1 = -19;
				 l_2 = -31; end
		38345: begin l_1 = +19;
				 l_2 = +32; end
		28194: begin l_1 = +19;
				 l_2 = -32; end
		22667: begin l_1 = -19;
				 l_2 = +32; end
		12516: begin l_1 = -19;
				 l_2 = -32; end
		17990: begin l_1 = +19;
				 l_2 = +33; end
		48549: begin l_1 = +19;
				 l_2 = -33; end
		2312: begin l_1 = -19;
				 l_2 = +33; end
		32871: begin l_1 = -19;
				 l_2 = -33; end
		28141: begin l_1 = +19;
				 l_2 = +34; end
		38398: begin l_1 = +19;
				 l_2 = -34; end
		12463: begin l_1 = -19;
				 l_2 = +34; end
		22720: begin l_1 = -19;
				 l_2 = -34; end
		48443: begin l_1 = +19;
				 l_2 = +35; end
		18096: begin l_1 = +19;
				 l_2 = -35; end
		32765: begin l_1 = -19;
				 l_2 = +35; end
		2418: begin l_1 = -19;
				 l_2 = -35; end
		38186: begin l_1 = +19;
				 l_2 = +36; end
		28353: begin l_1 = +19;
				 l_2 = -36; end
		22508: begin l_1 = -19;
				 l_2 = +36; end
		12675: begin l_1 = -19;
				 l_2 = -36; end
		17672: begin l_1 = +19;
				 l_2 = +37; end
		48867: begin l_1 = +19;
				 l_2 = -37; end
		1994: begin l_1 = -19;
				 l_2 = +37; end
		33189: begin l_1 = -19;
				 l_2 = -37; end
		27505: begin l_1 = +19;
				 l_2 = +38; end
		39034: begin l_1 = +19;
				 l_2 = -38; end
		11827: begin l_1 = -19;
				 l_2 = +38; end
		23356: begin l_1 = -19;
				 l_2 = -38; end
		47171: begin l_1 = +19;
				 l_2 = +39; end
		19368: begin l_1 = +19;
				 l_2 = -39; end
		31493: begin l_1 = -19;
				 l_2 = +39; end
		3690: begin l_1 = -19;
				 l_2 = -39; end
		35642: begin l_1 = +19;
				 l_2 = +40; end
		30897: begin l_1 = +19;
				 l_2 = -40; end
		19964: begin l_1 = -19;
				 l_2 = +40; end
		15219: begin l_1 = -19;
				 l_2 = -40; end
		12584: begin l_1 = +19;
				 l_2 = +41; end
		3094: begin l_1 = +19;
				 l_2 = -41; end
		47767: begin l_1 = -19;
				 l_2 = +41; end
		38277: begin l_1 = -19;
				 l_2 = -41; end
		17329: begin l_1 = +19;
				 l_2 = +42; end
		49210: begin l_1 = +19;
				 l_2 = -42; end
		1651: begin l_1 = -19;
				 l_2 = +42; end
		33532: begin l_1 = -19;
				 l_2 = -42; end
		26819: begin l_1 = +19;
				 l_2 = +43; end
		39720: begin l_1 = +19;
				 l_2 = -43; end
		11141: begin l_1 = -19;
				 l_2 = +43; end
		24042: begin l_1 = -19;
				 l_2 = -43; end
		45799: begin l_1 = +19;
				 l_2 = +44; end
		20740: begin l_1 = +19;
				 l_2 = -44; end
		30121: begin l_1 = -19;
				 l_2 = +44; end
		5062: begin l_1 = -19;
				 l_2 = -44; end
		32898: begin l_1 = +19;
				 l_2 = +45; end
		33641: begin l_1 = +19;
				 l_2 = -45; end
		17220: begin l_1 = -19;
				 l_2 = +45; end
		17963: begin l_1 = -19;
				 l_2 = -45; end
		7096: begin l_1 = +19;
				 l_2 = +46; end
		8582: begin l_1 = +19;
				 l_2 = -46; end
		42279: begin l_1 = -19;
				 l_2 = +46; end
		43765: begin l_1 = -19;
				 l_2 = -46; end
		6353: begin l_1 = +19;
				 l_2 = +47; end
		9325: begin l_1 = +19;
				 l_2 = -47; end
		41536: begin l_1 = -19;
				 l_2 = +47; end
		44508: begin l_1 = -19;
				 l_2 = -47; end
		4867: begin l_1 = +19;
				 l_2 = +48; end
		10811: begin l_1 = +19;
				 l_2 = -48; end
		40050: begin l_1 = -19;
				 l_2 = +48; end
		45994: begin l_1 = -19;
				 l_2 = -48; end
		1895: begin l_1 = +19;
				 l_2 = +49; end
		13783: begin l_1 = +19;
				 l_2 = -49; end
		37078: begin l_1 = -19;
				 l_2 = +49; end
		48966: begin l_1 = -19;
				 l_2 = -49; end
		46812: begin l_1 = +19;
				 l_2 = +50; end
		19727: begin l_1 = +19;
				 l_2 = -50; end
		31134: begin l_1 = -19;
				 l_2 = +50; end
		4049: begin l_1 = -19;
				 l_2 = -50; end
		34924: begin l_1 = +19;
				 l_2 = +51; end
		31615: begin l_1 = +19;
				 l_2 = -51; end
		19246: begin l_1 = -19;
				 l_2 = +51; end
		15937: begin l_1 = -19;
				 l_2 = -51; end
		11148: begin l_1 = +19;
				 l_2 = +52; end
		4530: begin l_1 = +19;
				 l_2 = -52; end
		46331: begin l_1 = -19;
				 l_2 = +52; end
		39713: begin l_1 = -19;
				 l_2 = -52; end
		14457: begin l_1 = +19;
				 l_2 = +53; end
		1221: begin l_1 = +19;
				 l_2 = -53; end
		49640: begin l_1 = -19;
				 l_2 = +53; end
		36404: begin l_1 = -19;
				 l_2 = -53; end
		21075: begin l_1 = +19;
				 l_2 = +54; end
		45464: begin l_1 = +19;
				 l_2 = -54; end
		5397: begin l_1 = -19;
				 l_2 = +54; end
		29786: begin l_1 = -19;
				 l_2 = -54; end
		34311: begin l_1 = +19;
				 l_2 = +55; end
		32228: begin l_1 = +19;
				 l_2 = -55; end
		18633: begin l_1 = -19;
				 l_2 = +55; end
		16550: begin l_1 = -19;
				 l_2 = -55; end
		9922: begin l_1 = +19;
				 l_2 = +56; end
		5756: begin l_1 = +19;
				 l_2 = -56; end
		45105: begin l_1 = -19;
				 l_2 = +56; end
		40939: begin l_1 = -19;
				 l_2 = -56; end
		12005: begin l_1 = +19;
				 l_2 = +57; end
		3673: begin l_1 = +19;
				 l_2 = -57; end
		47188: begin l_1 = -19;
				 l_2 = +57; end
		38856: begin l_1 = -19;
				 l_2 = -57; end
		16171: begin l_1 = +19;
				 l_2 = +58; end
		50368: begin l_1 = +19;
				 l_2 = -58; end
		493: begin l_1 = -19;
				 l_2 = +58; end
		34690: begin l_1 = -19;
				 l_2 = -58; end
		24503: begin l_1 = +19;
				 l_2 = +59; end
		42036: begin l_1 = +19;
				 l_2 = -59; end
		8825: begin l_1 = -19;
				 l_2 = +59; end
		26358: begin l_1 = -19;
				 l_2 = -59; end
		41167: begin l_1 = +19;
				 l_2 = +60; end
		25372: begin l_1 = +19;
				 l_2 = -60; end
		25489: begin l_1 = -19;
				 l_2 = +60; end
		9694: begin l_1 = -19;
				 l_2 = -60; end
		23634: begin l_1 = +19;
				 l_2 = +61; end
		42905: begin l_1 = +19;
				 l_2 = -61; end
		7956: begin l_1 = -19;
				 l_2 = +61; end
		27227: begin l_1 = -19;
				 l_2 = -61; end
		39429: begin l_1 = +19;
				 l_2 = +62; end
		27110: begin l_1 = +19;
				 l_2 = -62; end
		23751: begin l_1 = -19;
				 l_2 = +62; end
		11432: begin l_1 = -19;
				 l_2 = -62; end
		20158: begin l_1 = +19;
				 l_2 = +63; end
		46381: begin l_1 = +19;
				 l_2 = -63; end
		4480: begin l_1 = -19;
				 l_2 = +63; end
		30703: begin l_1 = -19;
				 l_2 = -63; end
		32477: begin l_1 = +19;
				 l_2 = +64; end
		34062: begin l_1 = +19;
				 l_2 = -64; end
		16799: begin l_1 = -19;
				 l_2 = +64; end
		18384: begin l_1 = -19;
				 l_2 = -64; end
		6254: begin l_1 = +19;
				 l_2 = +65; end
		9424: begin l_1 = +19;
				 l_2 = -65; end
		41437: begin l_1 = -19;
				 l_2 = +65; end
		44607: begin l_1 = -19;
				 l_2 = -65; end
		4669: begin l_1 = +19;
				 l_2 = +66; end
		11009: begin l_1 = +19;
				 l_2 = -66; end
		39852: begin l_1 = -19;
				 l_2 = +66; end
		46192: begin l_1 = -19;
				 l_2 = -66; end
		1499: begin l_1 = +19;
				 l_2 = +67; end
		14179: begin l_1 = +19;
				 l_2 = -67; end
		36682: begin l_1 = -19;
				 l_2 = +67; end
		49362: begin l_1 = -19;
				 l_2 = -67; end
		46020: begin l_1 = +19;
				 l_2 = +68; end
		20519: begin l_1 = +19;
				 l_2 = -68; end
		30342: begin l_1 = -19;
				 l_2 = +68; end
		4841: begin l_1 = -19;
				 l_2 = -68; end
		47034: begin l_1 = -20;
				 l_2 = +22; end
		3827: begin l_1 = -20;
				 l_2 = -21; end
		27529: begin l_1 = +20;
				 l_2 = +22; end
		23332: begin l_1 = -20;
				 l_2 = -22; end
		39380: begin l_1 = +20;
				 l_2 = +23; end
		42837: begin l_1 = +20;
				 l_2 = -23; end
		8024: begin l_1 = -20;
				 l_2 = +23; end
		11481: begin l_1 = -20;
				 l_2 = -23; end
		12221: begin l_1 = +20;
				 l_2 = +24; end
		19135: begin l_1 = +20;
				 l_2 = -24; end
		31726: begin l_1 = -20;
				 l_2 = +24; end
		38640: begin l_1 = -20;
				 l_2 = -24; end
		8764: begin l_1 = +20;
				 l_2 = +25; end
		22592: begin l_1 = +20;
				 l_2 = -25; end
		28269: begin l_1 = -20;
				 l_2 = +25; end
		42097: begin l_1 = -20;
				 l_2 = -25; end
		1850: begin l_1 = +20;
				 l_2 = +26; end
		29506: begin l_1 = +20;
				 l_2 = -26; end
		21355: begin l_1 = -20;
				 l_2 = +26; end
		49011: begin l_1 = -20;
				 l_2 = -26; end
		38883: begin l_1 = +20;
				 l_2 = +27; end
		43334: begin l_1 = +20;
				 l_2 = -27; end
		7527: begin l_1 = -20;
				 l_2 = +27; end
		11978: begin l_1 = -20;
				 l_2 = -27; end
		11227: begin l_1 = +20;
				 l_2 = +28; end
		20129: begin l_1 = +20;
				 l_2 = -28; end
		30732: begin l_1 = -20;
				 l_2 = +28; end
		39634: begin l_1 = -20;
				 l_2 = -28; end
		6776: begin l_1 = +20;
				 l_2 = +29; end
		24580: begin l_1 = +20;
				 l_2 = -29; end
		26281: begin l_1 = -20;
				 l_2 = +29; end
		44085: begin l_1 = -20;
				 l_2 = -29; end
		48735: begin l_1 = +20;
				 l_2 = +30; end
		33482: begin l_1 = +20;
				 l_2 = -30; end
		17379: begin l_1 = -20;
				 l_2 = +30; end
		2126: begin l_1 = -20;
				 l_2 = -30; end
		30931: begin l_1 = +20;
				 l_2 = +31; end
		425: begin l_1 = +20;
				 l_2 = -31; end
		50436: begin l_1 = -20;
				 l_2 = +31; end
		19930: begin l_1 = -20;
				 l_2 = -31; end
		46184: begin l_1 = +20;
				 l_2 = +32; end
		36033: begin l_1 = +20;
				 l_2 = -32; end
		14828: begin l_1 = -20;
				 l_2 = +32; end
		4677: begin l_1 = -20;
				 l_2 = -32; end
		25829: begin l_1 = +20;
				 l_2 = +33; end
		5527: begin l_1 = +20;
				 l_2 = -33; end
		45334: begin l_1 = -20;
				 l_2 = +33; end
		25032: begin l_1 = -20;
				 l_2 = -33; end
		35980: begin l_1 = +20;
				 l_2 = +34; end
		46237: begin l_1 = +20;
				 l_2 = -34; end
		4624: begin l_1 = -20;
				 l_2 = +34; end
		14881: begin l_1 = -20;
				 l_2 = -34; end
		5421: begin l_1 = +20;
				 l_2 = +35; end
		25935: begin l_1 = +20;
				 l_2 = -35; end
		24926: begin l_1 = -20;
				 l_2 = +35; end
		45440: begin l_1 = -20;
				 l_2 = -35; end
		46025: begin l_1 = +20;
				 l_2 = +36; end
		36192: begin l_1 = +20;
				 l_2 = -36; end
		14669: begin l_1 = -20;
				 l_2 = +36; end
		4836: begin l_1 = -20;
				 l_2 = -36; end
		25511: begin l_1 = +20;
				 l_2 = +37; end
		5845: begin l_1 = +20;
				 l_2 = -37; end
		45016: begin l_1 = -20;
				 l_2 = +37; end
		25350: begin l_1 = -20;
				 l_2 = -37; end
		35344: begin l_1 = +20;
				 l_2 = +38; end
		46873: begin l_1 = +20;
				 l_2 = -38; end
		3988: begin l_1 = -20;
				 l_2 = +38; end
		15517: begin l_1 = -20;
				 l_2 = -38; end
		4149: begin l_1 = +20;
				 l_2 = +39; end
		27207: begin l_1 = +20;
				 l_2 = -39; end
		23654: begin l_1 = -20;
				 l_2 = +39; end
		46712: begin l_1 = -20;
				 l_2 = -39; end
		43481: begin l_1 = +20;
				 l_2 = +40; end
		38736: begin l_1 = +20;
				 l_2 = -40; end
		12125: begin l_1 = -20;
				 l_2 = +40; end
		7380: begin l_1 = -20;
				 l_2 = -40; end
		20423: begin l_1 = +20;
				 l_2 = +41; end
		10933: begin l_1 = +20;
				 l_2 = -41; end
		39928: begin l_1 = -20;
				 l_2 = +41; end
		30438: begin l_1 = -20;
				 l_2 = -41; end
		25168: begin l_1 = +20;
				 l_2 = +42; end
		6188: begin l_1 = +20;
				 l_2 = -42; end
		44673: begin l_1 = -20;
				 l_2 = +42; end
		25693: begin l_1 = -20;
				 l_2 = -42; end
		34658: begin l_1 = +20;
				 l_2 = +43; end
		47559: begin l_1 = +20;
				 l_2 = -43; end
		3302: begin l_1 = -20;
				 l_2 = +43; end
		16203: begin l_1 = -20;
				 l_2 = -43; end
		2777: begin l_1 = +20;
				 l_2 = +44; end
		28579: begin l_1 = +20;
				 l_2 = -44; end
		22282: begin l_1 = -20;
				 l_2 = +44; end
		48084: begin l_1 = -20;
				 l_2 = -44; end
		40737: begin l_1 = +20;
				 l_2 = +45; end
		41480: begin l_1 = +20;
				 l_2 = -45; end
		9381: begin l_1 = -20;
				 l_2 = +45; end
		10124: begin l_1 = -20;
				 l_2 = -45; end
		14935: begin l_1 = +20;
				 l_2 = +46; end
		16421: begin l_1 = +20;
				 l_2 = -46; end
		34440: begin l_1 = -20;
				 l_2 = +46; end
		35926: begin l_1 = -20;
				 l_2 = -46; end
		14192: begin l_1 = +20;
				 l_2 = +47; end
		17164: begin l_1 = +20;
				 l_2 = -47; end
		33697: begin l_1 = -20;
				 l_2 = +47; end
		36669: begin l_1 = -20;
				 l_2 = -47; end
		12706: begin l_1 = +20;
				 l_2 = +48; end
		18650: begin l_1 = +20;
				 l_2 = -48; end
		32211: begin l_1 = -20;
				 l_2 = +48; end
		38155: begin l_1 = -20;
				 l_2 = -48; end
		9734: begin l_1 = +20;
				 l_2 = +49; end
		21622: begin l_1 = +20;
				 l_2 = -49; end
		29239: begin l_1 = -20;
				 l_2 = +49; end
		41127: begin l_1 = -20;
				 l_2 = -49; end
		3790: begin l_1 = +20;
				 l_2 = +50; end
		27566: begin l_1 = +20;
				 l_2 = -50; end
		23295: begin l_1 = -20;
				 l_2 = +50; end
		47071: begin l_1 = -20;
				 l_2 = -50; end
		42763: begin l_1 = +20;
				 l_2 = +51; end
		39454: begin l_1 = +20;
				 l_2 = -51; end
		11407: begin l_1 = -20;
				 l_2 = +51; end
		8098: begin l_1 = -20;
				 l_2 = -51; end
		18987: begin l_1 = +20;
				 l_2 = +52; end
		12369: begin l_1 = +20;
				 l_2 = -52; end
		38492: begin l_1 = -20;
				 l_2 = +52; end
		31874: begin l_1 = -20;
				 l_2 = -52; end
		22296: begin l_1 = +20;
				 l_2 = +53; end
		9060: begin l_1 = +20;
				 l_2 = -53; end
		41801: begin l_1 = -20;
				 l_2 = +53; end
		28565: begin l_1 = -20;
				 l_2 = -53; end
		28914: begin l_1 = +20;
				 l_2 = +54; end
		2442: begin l_1 = +20;
				 l_2 = -54; end
		48419: begin l_1 = -20;
				 l_2 = +54; end
		21947: begin l_1 = -20;
				 l_2 = -54; end
		42150: begin l_1 = +20;
				 l_2 = +55; end
		40067: begin l_1 = +20;
				 l_2 = -55; end
		10794: begin l_1 = -20;
				 l_2 = +55; end
		8711: begin l_1 = -20;
				 l_2 = -55; end
		17761: begin l_1 = +20;
				 l_2 = +56; end
		13595: begin l_1 = +20;
				 l_2 = -56; end
		37266: begin l_1 = -20;
				 l_2 = +56; end
		33100: begin l_1 = -20;
				 l_2 = -56; end
		19844: begin l_1 = +20;
				 l_2 = +57; end
		11512: begin l_1 = +20;
				 l_2 = -57; end
		39349: begin l_1 = -20;
				 l_2 = +57; end
		31017: begin l_1 = -20;
				 l_2 = -57; end
		24010: begin l_1 = +20;
				 l_2 = +58; end
		7346: begin l_1 = +20;
				 l_2 = -58; end
		43515: begin l_1 = -20;
				 l_2 = +58; end
		26851: begin l_1 = -20;
				 l_2 = -58; end
		32342: begin l_1 = +20;
				 l_2 = +59; end
		49875: begin l_1 = +20;
				 l_2 = -59; end
		986: begin l_1 = -20;
				 l_2 = +59; end
		18519: begin l_1 = -20;
				 l_2 = -59; end
		49006: begin l_1 = +20;
				 l_2 = +60; end
		33211: begin l_1 = +20;
				 l_2 = -60; end
		17650: begin l_1 = -20;
				 l_2 = +60; end
		1855: begin l_1 = -20;
				 l_2 = -60; end
		31473: begin l_1 = +20;
				 l_2 = +61; end
		50744: begin l_1 = +20;
				 l_2 = -61; end
		117: begin l_1 = -20;
				 l_2 = +61; end
		19388: begin l_1 = -20;
				 l_2 = -61; end
		47268: begin l_1 = +20;
				 l_2 = +62; end
		34949: begin l_1 = +20;
				 l_2 = -62; end
		15912: begin l_1 = -20;
				 l_2 = +62; end
		3593: begin l_1 = -20;
				 l_2 = -62; end
		27997: begin l_1 = +20;
				 l_2 = +63; end
		3359: begin l_1 = +20;
				 l_2 = -63; end
		47502: begin l_1 = -20;
				 l_2 = +63; end
		22864: begin l_1 = -20;
				 l_2 = -63; end
		40316: begin l_1 = +20;
				 l_2 = +64; end
		41901: begin l_1 = +20;
				 l_2 = -64; end
		8960: begin l_1 = -20;
				 l_2 = +64; end
		10545: begin l_1 = -20;
				 l_2 = -64; end
		14093: begin l_1 = +20;
				 l_2 = +65; end
		17263: begin l_1 = +20;
				 l_2 = -65; end
		33598: begin l_1 = -20;
				 l_2 = +65; end
		36768: begin l_1 = -20;
				 l_2 = -65; end
		12508: begin l_1 = +20;
				 l_2 = +66; end
		18848: begin l_1 = +20;
				 l_2 = -66; end
		32013: begin l_1 = -20;
				 l_2 = +66; end
		38353: begin l_1 = -20;
				 l_2 = -66; end
		9338: begin l_1 = +20;
				 l_2 = +67; end
		22018: begin l_1 = +20;
				 l_2 = -67; end
		28843: begin l_1 = -20;
				 l_2 = +67; end
		41523: begin l_1 = -20;
				 l_2 = -67; end
		2998: begin l_1 = +20;
				 l_2 = +68; end
		28358: begin l_1 = +20;
				 l_2 = -68; end
		22503: begin l_1 = -20;
				 l_2 = +68; end
		47863: begin l_1 = -20;
				 l_2 = -68; end
		43207: begin l_1 = -21;
				 l_2 = +23; end
		7654: begin l_1 = -21;
				 l_2 = -22; end
		4197: begin l_1 = +21;
				 l_2 = +23; end
		46664: begin l_1 = -21;
				 l_2 = -23; end
		27899: begin l_1 = +21;
				 l_2 = +24; end
		34813: begin l_1 = +21;
				 l_2 = -24; end
		16048: begin l_1 = -21;
				 l_2 = +24; end
		22962: begin l_1 = -21;
				 l_2 = -24; end
		24442: begin l_1 = +21;
				 l_2 = +25; end
		38270: begin l_1 = +21;
				 l_2 = -25; end
		12591: begin l_1 = -21;
				 l_2 = +25; end
		26419: begin l_1 = -21;
				 l_2 = -25; end
		17528: begin l_1 = +21;
				 l_2 = +26; end
		45184: begin l_1 = +21;
				 l_2 = -26; end
		5677: begin l_1 = -21;
				 l_2 = +26; end
		33333: begin l_1 = -21;
				 l_2 = -26; end
		3700: begin l_1 = +21;
				 l_2 = +27; end
		8151: begin l_1 = +21;
				 l_2 = -27; end
		42710: begin l_1 = -21;
				 l_2 = +27; end
		47161: begin l_1 = -21;
				 l_2 = -27; end
		26905: begin l_1 = +21;
				 l_2 = +28; end
		35807: begin l_1 = +21;
				 l_2 = -28; end
		15054: begin l_1 = -21;
				 l_2 = +28; end
		23956: begin l_1 = -21;
				 l_2 = -28; end
		22454: begin l_1 = +21;
				 l_2 = +29; end
		40258: begin l_1 = +21;
				 l_2 = -29; end
		10603: begin l_1 = -21;
				 l_2 = +29; end
		28407: begin l_1 = -21;
				 l_2 = -29; end
		13552: begin l_1 = +21;
				 l_2 = +30; end
		49160: begin l_1 = +21;
				 l_2 = -30; end
		1701: begin l_1 = -21;
				 l_2 = +30; end
		37309: begin l_1 = -21;
				 l_2 = -30; end
		46609: begin l_1 = +21;
				 l_2 = +31; end
		16103: begin l_1 = +21;
				 l_2 = -31; end
		34758: begin l_1 = -21;
				 l_2 = +31; end
		4252: begin l_1 = -21;
				 l_2 = -31; end
		11001: begin l_1 = +21;
				 l_2 = +32; end
		850: begin l_1 = +21;
				 l_2 = -32; end
		50011: begin l_1 = -21;
				 l_2 = +32; end
		39860: begin l_1 = -21;
				 l_2 = -32; end
		41507: begin l_1 = +21;
				 l_2 = +33; end
		21205: begin l_1 = +21;
				 l_2 = -33; end
		29656: begin l_1 = -21;
				 l_2 = +33; end
		9354: begin l_1 = -21;
				 l_2 = -33; end
		797: begin l_1 = +21;
				 l_2 = +34; end
		11054: begin l_1 = +21;
				 l_2 = -34; end
		39807: begin l_1 = -21;
				 l_2 = +34; end
		50064: begin l_1 = -21;
				 l_2 = -34; end
		21099: begin l_1 = +21;
				 l_2 = +35; end
		41613: begin l_1 = +21;
				 l_2 = -35; end
		9248: begin l_1 = -21;
				 l_2 = +35; end
		29762: begin l_1 = -21;
				 l_2 = -35; end
		10842: begin l_1 = +21;
				 l_2 = +36; end
		1009: begin l_1 = +21;
				 l_2 = -36; end
		49852: begin l_1 = -21;
				 l_2 = +36; end
		40019: begin l_1 = -21;
				 l_2 = -36; end
		41189: begin l_1 = +21;
				 l_2 = +37; end
		21523: begin l_1 = +21;
				 l_2 = -37; end
		29338: begin l_1 = -21;
				 l_2 = +37; end
		9672: begin l_1 = -21;
				 l_2 = -37; end
		161: begin l_1 = +21;
				 l_2 = +38; end
		11690: begin l_1 = +21;
				 l_2 = -38; end
		39171: begin l_1 = -21;
				 l_2 = +38; end
		50700: begin l_1 = -21;
				 l_2 = -38; end
		19827: begin l_1 = +21;
				 l_2 = +39; end
		42885: begin l_1 = +21;
				 l_2 = -39; end
		7976: begin l_1 = -21;
				 l_2 = +39; end
		31034: begin l_1 = -21;
				 l_2 = -39; end
		8298: begin l_1 = +21;
				 l_2 = +40; end
		3553: begin l_1 = +21;
				 l_2 = -40; end
		47308: begin l_1 = -21;
				 l_2 = +40; end
		42563: begin l_1 = -21;
				 l_2 = -40; end
		36101: begin l_1 = +21;
				 l_2 = +41; end
		26611: begin l_1 = +21;
				 l_2 = -41; end
		24250: begin l_1 = -21;
				 l_2 = +41; end
		14760: begin l_1 = -21;
				 l_2 = -41; end
		40846: begin l_1 = +21;
				 l_2 = +42; end
		21866: begin l_1 = +21;
				 l_2 = -42; end
		28995: begin l_1 = -21;
				 l_2 = +42; end
		10015: begin l_1 = -21;
				 l_2 = -42; end
		50336: begin l_1 = +21;
				 l_2 = +43; end
		12376: begin l_1 = +21;
				 l_2 = -43; end
		38485: begin l_1 = -21;
				 l_2 = +43; end
		525: begin l_1 = -21;
				 l_2 = -43; end
		18455: begin l_1 = +21;
				 l_2 = +44; end
		44257: begin l_1 = +21;
				 l_2 = -44; end
		6604: begin l_1 = -21;
				 l_2 = +44; end
		32406: begin l_1 = -21;
				 l_2 = -44; end
		5554: begin l_1 = +21;
				 l_2 = +45; end
		6297: begin l_1 = +21;
				 l_2 = -45; end
		44564: begin l_1 = -21;
				 l_2 = +45; end
		45307: begin l_1 = -21;
				 l_2 = -45; end
		30613: begin l_1 = +21;
				 l_2 = +46; end
		32099: begin l_1 = +21;
				 l_2 = -46; end
		18762: begin l_1 = -21;
				 l_2 = +46; end
		20248: begin l_1 = -21;
				 l_2 = -46; end
		29870: begin l_1 = +21;
				 l_2 = +47; end
		32842: begin l_1 = +21;
				 l_2 = -47; end
		18019: begin l_1 = -21;
				 l_2 = +47; end
		20991: begin l_1 = -21;
				 l_2 = -47; end
		28384: begin l_1 = +21;
				 l_2 = +48; end
		34328: begin l_1 = +21;
				 l_2 = -48; end
		16533: begin l_1 = -21;
				 l_2 = +48; end
		22477: begin l_1 = -21;
				 l_2 = -48; end
		25412: begin l_1 = +21;
				 l_2 = +49; end
		37300: begin l_1 = +21;
				 l_2 = -49; end
		13561: begin l_1 = -21;
				 l_2 = +49; end
		25449: begin l_1 = -21;
				 l_2 = -49; end
		19468: begin l_1 = +21;
				 l_2 = +50; end
		43244: begin l_1 = +21;
				 l_2 = -50; end
		7617: begin l_1 = -21;
				 l_2 = +50; end
		31393: begin l_1 = -21;
				 l_2 = -50; end
		7580: begin l_1 = +21;
				 l_2 = +51; end
		4271: begin l_1 = +21;
				 l_2 = -51; end
		46590: begin l_1 = -21;
				 l_2 = +51; end
		43281: begin l_1 = -21;
				 l_2 = -51; end
		34665: begin l_1 = +21;
				 l_2 = +52; end
		28047: begin l_1 = +21;
				 l_2 = -52; end
		22814: begin l_1 = -21;
				 l_2 = +52; end
		16196: begin l_1 = -21;
				 l_2 = -52; end
		37974: begin l_1 = +21;
				 l_2 = +53; end
		24738: begin l_1 = +21;
				 l_2 = -53; end
		26123: begin l_1 = -21;
				 l_2 = +53; end
		12887: begin l_1 = -21;
				 l_2 = -53; end
		44592: begin l_1 = +21;
				 l_2 = +54; end
		18120: begin l_1 = +21;
				 l_2 = -54; end
		32741: begin l_1 = -21;
				 l_2 = +54; end
		6269: begin l_1 = -21;
				 l_2 = -54; end
		6967: begin l_1 = +21;
				 l_2 = +55; end
		4884: begin l_1 = +21;
				 l_2 = -55; end
		45977: begin l_1 = -21;
				 l_2 = +55; end
		43894: begin l_1 = -21;
				 l_2 = -55; end
		33439: begin l_1 = +21;
				 l_2 = +56; end
		29273: begin l_1 = +21;
				 l_2 = -56; end
		21588: begin l_1 = -21;
				 l_2 = +56; end
		17422: begin l_1 = -21;
				 l_2 = -56; end
		35522: begin l_1 = +21;
				 l_2 = +57; end
		27190: begin l_1 = +21;
				 l_2 = -57; end
		23671: begin l_1 = -21;
				 l_2 = +57; end
		15339: begin l_1 = -21;
				 l_2 = -57; end
		39688: begin l_1 = +21;
				 l_2 = +58; end
		23024: begin l_1 = +21;
				 l_2 = -58; end
		27837: begin l_1 = -21;
				 l_2 = +58; end
		11173: begin l_1 = -21;
				 l_2 = -58; end
		48020: begin l_1 = +21;
				 l_2 = +59; end
		14692: begin l_1 = +21;
				 l_2 = -59; end
		36169: begin l_1 = -21;
				 l_2 = +59; end
		2841: begin l_1 = -21;
				 l_2 = -59; end
		13823: begin l_1 = +21;
				 l_2 = +60; end
		48889: begin l_1 = +21;
				 l_2 = -60; end
		1972: begin l_1 = -21;
				 l_2 = +60; end
		37038: begin l_1 = -21;
				 l_2 = -60; end
		47151: begin l_1 = +21;
				 l_2 = +61; end
		15561: begin l_1 = +21;
				 l_2 = -61; end
		35300: begin l_1 = -21;
				 l_2 = +61; end
		3710: begin l_1 = -21;
				 l_2 = -61; end
		12085: begin l_1 = +21;
				 l_2 = +62; end
		50627: begin l_1 = +21;
				 l_2 = -62; end
		234: begin l_1 = -21;
				 l_2 = +62; end
		38776: begin l_1 = -21;
				 l_2 = -62; end
		43675: begin l_1 = +21;
				 l_2 = +63; end
		19037: begin l_1 = +21;
				 l_2 = -63; end
		31824: begin l_1 = -21;
				 l_2 = +63; end
		7186: begin l_1 = -21;
				 l_2 = -63; end
		5133: begin l_1 = +21;
				 l_2 = +64; end
		6718: begin l_1 = +21;
				 l_2 = -64; end
		44143: begin l_1 = -21;
				 l_2 = +64; end
		45728: begin l_1 = -21;
				 l_2 = -64; end
		29771: begin l_1 = +21;
				 l_2 = +65; end
		32941: begin l_1 = +21;
				 l_2 = -65; end
		17920: begin l_1 = -21;
				 l_2 = +65; end
		21090: begin l_1 = -21;
				 l_2 = -65; end
		28186: begin l_1 = +21;
				 l_2 = +66; end
		34526: begin l_1 = +21;
				 l_2 = -66; end
		16335: begin l_1 = -21;
				 l_2 = +66; end
		22675: begin l_1 = -21;
				 l_2 = -66; end
		25016: begin l_1 = +21;
				 l_2 = +67; end
		37696: begin l_1 = +21;
				 l_2 = -67; end
		13165: begin l_1 = -21;
				 l_2 = +67; end
		25845: begin l_1 = -21;
				 l_2 = -67; end
		18676: begin l_1 = +21;
				 l_2 = +68; end
		44036: begin l_1 = +21;
				 l_2 = -68; end
		6825: begin l_1 = -21;
				 l_2 = +68; end
		32185: begin l_1 = -21;
				 l_2 = -68; end
		35553: begin l_1 = -22;
				 l_2 = +24; end
		15308: begin l_1 = -22;
				 l_2 = -23; end
		8394: begin l_1 = +22;
				 l_2 = +24; end
		42467: begin l_1 = -22;
				 l_2 = -24; end
		4937: begin l_1 = +22;
				 l_2 = +25; end
		18765: begin l_1 = +22;
				 l_2 = -25; end
		32096: begin l_1 = -22;
				 l_2 = +25; end
		45924: begin l_1 = -22;
				 l_2 = -25; end
		48884: begin l_1 = +22;
				 l_2 = +26; end
		25679: begin l_1 = +22;
				 l_2 = -26; end
		25182: begin l_1 = -22;
				 l_2 = +26; end
		1977: begin l_1 = -22;
				 l_2 = -26; end
		35056: begin l_1 = +22;
				 l_2 = +27; end
		39507: begin l_1 = +22;
				 l_2 = -27; end
		11354: begin l_1 = -22;
				 l_2 = +27; end
		15805: begin l_1 = -22;
				 l_2 = -27; end
		7400: begin l_1 = +22;
				 l_2 = +28; end
		16302: begin l_1 = +22;
				 l_2 = -28; end
		34559: begin l_1 = -22;
				 l_2 = +28; end
		43461: begin l_1 = -22;
				 l_2 = -28; end
		2949: begin l_1 = +22;
				 l_2 = +29; end
		20753: begin l_1 = +22;
				 l_2 = -29; end
		30108: begin l_1 = -22;
				 l_2 = +29; end
		47912: begin l_1 = -22;
				 l_2 = -29; end
		44908: begin l_1 = +22;
				 l_2 = +30; end
		29655: begin l_1 = +22;
				 l_2 = -30; end
		21206: begin l_1 = -22;
				 l_2 = +30; end
		5953: begin l_1 = -22;
				 l_2 = -30; end
		27104: begin l_1 = +22;
				 l_2 = +31; end
		47459: begin l_1 = +22;
				 l_2 = -31; end
		3402: begin l_1 = -22;
				 l_2 = +31; end
		23757: begin l_1 = -22;
				 l_2 = -31; end
		42357: begin l_1 = +22;
				 l_2 = +32; end
		32206: begin l_1 = +22;
				 l_2 = -32; end
		18655: begin l_1 = -22;
				 l_2 = +32; end
		8504: begin l_1 = -22;
				 l_2 = -32; end
		22002: begin l_1 = +22;
				 l_2 = +33; end
		1700: begin l_1 = +22;
				 l_2 = -33; end
		49161: begin l_1 = -22;
				 l_2 = +33; end
		28859: begin l_1 = -22;
				 l_2 = -33; end
		32153: begin l_1 = +22;
				 l_2 = +34; end
		42410: begin l_1 = +22;
				 l_2 = -34; end
		8451: begin l_1 = -22;
				 l_2 = +34; end
		18708: begin l_1 = -22;
				 l_2 = -34; end
		1594: begin l_1 = +22;
				 l_2 = +35; end
		22108: begin l_1 = +22;
				 l_2 = -35; end
		28753: begin l_1 = -22;
				 l_2 = +35; end
		49267: begin l_1 = -22;
				 l_2 = -35; end
		42198: begin l_1 = +22;
				 l_2 = +36; end
		32365: begin l_1 = +22;
				 l_2 = -36; end
		18496: begin l_1 = -22;
				 l_2 = +36; end
		8663: begin l_1 = -22;
				 l_2 = -36; end
		21684: begin l_1 = +22;
				 l_2 = +37; end
		2018: begin l_1 = +22;
				 l_2 = -37; end
		48843: begin l_1 = -22;
				 l_2 = +37; end
		29177: begin l_1 = -22;
				 l_2 = -37; end
		31517: begin l_1 = +22;
				 l_2 = +38; end
		43046: begin l_1 = +22;
				 l_2 = -38; end
		7815: begin l_1 = -22;
				 l_2 = +38; end
		19344: begin l_1 = -22;
				 l_2 = -38; end
		322: begin l_1 = +22;
				 l_2 = +39; end
		23380: begin l_1 = +22;
				 l_2 = -39; end
		27481: begin l_1 = -22;
				 l_2 = +39; end
		50539: begin l_1 = -22;
				 l_2 = -39; end
		39654: begin l_1 = +22;
				 l_2 = +40; end
		34909: begin l_1 = +22;
				 l_2 = -40; end
		15952: begin l_1 = -22;
				 l_2 = +40; end
		11207: begin l_1 = -22;
				 l_2 = -40; end
		16596: begin l_1 = +22;
				 l_2 = +41; end
		7106: begin l_1 = +22;
				 l_2 = -41; end
		43755: begin l_1 = -22;
				 l_2 = +41; end
		34265: begin l_1 = -22;
				 l_2 = -41; end
		21341: begin l_1 = +22;
				 l_2 = +42; end
		2361: begin l_1 = +22;
				 l_2 = -42; end
		48500: begin l_1 = -22;
				 l_2 = +42; end
		29520: begin l_1 = -22;
				 l_2 = -42; end
		30831: begin l_1 = +22;
				 l_2 = +43; end
		43732: begin l_1 = +22;
				 l_2 = -43; end
		7129: begin l_1 = -22;
				 l_2 = +43; end
		20030: begin l_1 = -22;
				 l_2 = -43; end
		49811: begin l_1 = +22;
				 l_2 = +44; end
		24752: begin l_1 = +22;
				 l_2 = -44; end
		26109: begin l_1 = -22;
				 l_2 = +44; end
		1050: begin l_1 = -22;
				 l_2 = -44; end
		36910: begin l_1 = +22;
				 l_2 = +45; end
		37653: begin l_1 = +22;
				 l_2 = -45; end
		13208: begin l_1 = -22;
				 l_2 = +45; end
		13951: begin l_1 = -22;
				 l_2 = -45; end
		11108: begin l_1 = +22;
				 l_2 = +46; end
		12594: begin l_1 = +22;
				 l_2 = -46; end
		38267: begin l_1 = -22;
				 l_2 = +46; end
		39753: begin l_1 = -22;
				 l_2 = -46; end
		10365: begin l_1 = +22;
				 l_2 = +47; end
		13337: begin l_1 = +22;
				 l_2 = -47; end
		37524: begin l_1 = -22;
				 l_2 = +47; end
		40496: begin l_1 = -22;
				 l_2 = -47; end
		8879: begin l_1 = +22;
				 l_2 = +48; end
		14823: begin l_1 = +22;
				 l_2 = -48; end
		36038: begin l_1 = -22;
				 l_2 = +48; end
		41982: begin l_1 = -22;
				 l_2 = -48; end
		5907: begin l_1 = +22;
				 l_2 = +49; end
		17795: begin l_1 = +22;
				 l_2 = -49; end
		33066: begin l_1 = -22;
				 l_2 = +49; end
		44954: begin l_1 = -22;
				 l_2 = -49; end
		50824: begin l_1 = +22;
				 l_2 = +50; end
		23739: begin l_1 = +22;
				 l_2 = -50; end
		27122: begin l_1 = -22;
				 l_2 = +50; end
		37: begin l_1 = -22;
				 l_2 = -50; end
		38936: begin l_1 = +22;
				 l_2 = +51; end
		35627: begin l_1 = +22;
				 l_2 = -51; end
		15234: begin l_1 = -22;
				 l_2 = +51; end
		11925: begin l_1 = -22;
				 l_2 = -51; end
		15160: begin l_1 = +22;
				 l_2 = +52; end
		8542: begin l_1 = +22;
				 l_2 = -52; end
		42319: begin l_1 = -22;
				 l_2 = +52; end
		35701: begin l_1 = -22;
				 l_2 = -52; end
		18469: begin l_1 = +22;
				 l_2 = +53; end
		5233: begin l_1 = +22;
				 l_2 = -53; end
		45628: begin l_1 = -22;
				 l_2 = +53; end
		32392: begin l_1 = -22;
				 l_2 = -53; end
		25087: begin l_1 = +22;
				 l_2 = +54; end
		49476: begin l_1 = +22;
				 l_2 = -54; end
		1385: begin l_1 = -22;
				 l_2 = +54; end
		25774: begin l_1 = -22;
				 l_2 = -54; end
		38323: begin l_1 = +22;
				 l_2 = +55; end
		36240: begin l_1 = +22;
				 l_2 = -55; end
		14621: begin l_1 = -22;
				 l_2 = +55; end
		12538: begin l_1 = -22;
				 l_2 = -55; end
		13934: begin l_1 = +22;
				 l_2 = +56; end
		9768: begin l_1 = +22;
				 l_2 = -56; end
		41093: begin l_1 = -22;
				 l_2 = +56; end
		36927: begin l_1 = -22;
				 l_2 = -56; end
		16017: begin l_1 = +22;
				 l_2 = +57; end
		7685: begin l_1 = +22;
				 l_2 = -57; end
		43176: begin l_1 = -22;
				 l_2 = +57; end
		34844: begin l_1 = -22;
				 l_2 = -57; end
		20183: begin l_1 = +22;
				 l_2 = +58; end
		3519: begin l_1 = +22;
				 l_2 = -58; end
		47342: begin l_1 = -22;
				 l_2 = +58; end
		30678: begin l_1 = -22;
				 l_2 = -58; end
		28515: begin l_1 = +22;
				 l_2 = +59; end
		46048: begin l_1 = +22;
				 l_2 = -59; end
		4813: begin l_1 = -22;
				 l_2 = +59; end
		22346: begin l_1 = -22;
				 l_2 = -59; end
		45179: begin l_1 = +22;
				 l_2 = +60; end
		29384: begin l_1 = +22;
				 l_2 = -60; end
		21477: begin l_1 = -22;
				 l_2 = +60; end
		5682: begin l_1 = -22;
				 l_2 = -60; end
		27646: begin l_1 = +22;
				 l_2 = +61; end
		46917: begin l_1 = +22;
				 l_2 = -61; end
		3944: begin l_1 = -22;
				 l_2 = +61; end
		23215: begin l_1 = -22;
				 l_2 = -61; end
		43441: begin l_1 = +22;
				 l_2 = +62; end
		31122: begin l_1 = +22;
				 l_2 = -62; end
		19739: begin l_1 = -22;
				 l_2 = +62; end
		7420: begin l_1 = -22;
				 l_2 = -62; end
		24170: begin l_1 = +22;
				 l_2 = +63; end
		50393: begin l_1 = +22;
				 l_2 = -63; end
		468: begin l_1 = -22;
				 l_2 = +63; end
		26691: begin l_1 = -22;
				 l_2 = -63; end
		36489: begin l_1 = +22;
				 l_2 = +64; end
		38074: begin l_1 = +22;
				 l_2 = -64; end
		12787: begin l_1 = -22;
				 l_2 = +64; end
		14372: begin l_1 = -22;
				 l_2 = -64; end
		10266: begin l_1 = +22;
				 l_2 = +65; end
		13436: begin l_1 = +22;
				 l_2 = -65; end
		37425: begin l_1 = -22;
				 l_2 = +65; end
		40595: begin l_1 = -22;
				 l_2 = -65; end
		8681: begin l_1 = +22;
				 l_2 = +66; end
		15021: begin l_1 = +22;
				 l_2 = -66; end
		35840: begin l_1 = -22;
				 l_2 = +66; end
		42180: begin l_1 = -22;
				 l_2 = -66; end
		5511: begin l_1 = +22;
				 l_2 = +67; end
		18191: begin l_1 = +22;
				 l_2 = -67; end
		32670: begin l_1 = -22;
				 l_2 = +67; end
		45350: begin l_1 = -22;
				 l_2 = -67; end
		50032: begin l_1 = +22;
				 l_2 = +68; end
		24531: begin l_1 = +22;
				 l_2 = -68; end
		26330: begin l_1 = -22;
				 l_2 = +68; end
		829: begin l_1 = -22;
				 l_2 = -68; end
		20245: begin l_1 = -23;
				 l_2 = +25; end
		30616: begin l_1 = -23;
				 l_2 = -24; end
		16788: begin l_1 = +23;
				 l_2 = +25; end
		34073: begin l_1 = -23;
				 l_2 = -25; end
		9874: begin l_1 = +23;
				 l_2 = +26; end
		37530: begin l_1 = +23;
				 l_2 = -26; end
		13331: begin l_1 = -23;
				 l_2 = +26; end
		40987: begin l_1 = -23;
				 l_2 = -26; end
		46907: begin l_1 = +23;
				 l_2 = +27; end
		497: begin l_1 = +23;
				 l_2 = -27; end
		50364: begin l_1 = -23;
				 l_2 = +27; end
		3954: begin l_1 = -23;
				 l_2 = -27; end
		19251: begin l_1 = +23;
				 l_2 = +28; end
		28153: begin l_1 = +23;
				 l_2 = -28; end
		22708: begin l_1 = -23;
				 l_2 = +28; end
		31610: begin l_1 = -23;
				 l_2 = -28; end
		14800: begin l_1 = +23;
				 l_2 = +29; end
		32604: begin l_1 = +23;
				 l_2 = -29; end
		18257: begin l_1 = -23;
				 l_2 = +29; end
		36061: begin l_1 = -23;
				 l_2 = -29; end
		5898: begin l_1 = +23;
				 l_2 = +30; end
		41506: begin l_1 = +23;
				 l_2 = -30; end
		9355: begin l_1 = -23;
				 l_2 = +30; end
		44963: begin l_1 = -23;
				 l_2 = -30; end
		38955: begin l_1 = +23;
				 l_2 = +31; end
		8449: begin l_1 = +23;
				 l_2 = -31; end
		42412: begin l_1 = -23;
				 l_2 = +31; end
		11906: begin l_1 = -23;
				 l_2 = -31; end
		3347: begin l_1 = +23;
				 l_2 = +32; end
		44057: begin l_1 = +23;
				 l_2 = -32; end
		6804: begin l_1 = -23;
				 l_2 = +32; end
		47514: begin l_1 = -23;
				 l_2 = -32; end
		33853: begin l_1 = +23;
				 l_2 = +33; end
		13551: begin l_1 = +23;
				 l_2 = -33; end
		37310: begin l_1 = -23;
				 l_2 = +33; end
		17008: begin l_1 = -23;
				 l_2 = -33; end
		44004: begin l_1 = +23;
				 l_2 = +34; end
		3400: begin l_1 = +23;
				 l_2 = -34; end
		47461: begin l_1 = -23;
				 l_2 = +34; end
		6857: begin l_1 = -23;
				 l_2 = -34; end
		13445: begin l_1 = +23;
				 l_2 = +35; end
		33959: begin l_1 = +23;
				 l_2 = -35; end
		16902: begin l_1 = -23;
				 l_2 = +35; end
		37416: begin l_1 = -23;
				 l_2 = -35; end
		3188: begin l_1 = +23;
				 l_2 = +36; end
		44216: begin l_1 = +23;
				 l_2 = -36; end
		6645: begin l_1 = -23;
				 l_2 = +36; end
		47673: begin l_1 = -23;
				 l_2 = -36; end
		33535: begin l_1 = +23;
				 l_2 = +37; end
		13869: begin l_1 = +23;
				 l_2 = -37; end
		36992: begin l_1 = -23;
				 l_2 = +37; end
		17326: begin l_1 = -23;
				 l_2 = -37; end
		43368: begin l_1 = +23;
				 l_2 = +38; end
		4036: begin l_1 = +23;
				 l_2 = -38; end
		46825: begin l_1 = -23;
				 l_2 = +38; end
		7493: begin l_1 = -23;
				 l_2 = -38; end
		12173: begin l_1 = +23;
				 l_2 = +39; end
		35231: begin l_1 = +23;
				 l_2 = -39; end
		15630: begin l_1 = -23;
				 l_2 = +39; end
		38688: begin l_1 = -23;
				 l_2 = -39; end
		644: begin l_1 = +23;
				 l_2 = +40; end
		46760: begin l_1 = +23;
				 l_2 = -40; end
		4101: begin l_1 = -23;
				 l_2 = +40; end
		50217: begin l_1 = -23;
				 l_2 = -40; end
		28447: begin l_1 = +23;
				 l_2 = +41; end
		18957: begin l_1 = +23;
				 l_2 = -41; end
		31904: begin l_1 = -23;
				 l_2 = +41; end
		22414: begin l_1 = -23;
				 l_2 = -41; end
		33192: begin l_1 = +23;
				 l_2 = +42; end
		14212: begin l_1 = +23;
				 l_2 = -42; end
		36649: begin l_1 = -23;
				 l_2 = +42; end
		17669: begin l_1 = -23;
				 l_2 = -42; end
		42682: begin l_1 = +23;
				 l_2 = +43; end
		4722: begin l_1 = +23;
				 l_2 = -43; end
		46139: begin l_1 = -23;
				 l_2 = +43; end
		8179: begin l_1 = -23;
				 l_2 = -43; end
		10801: begin l_1 = +23;
				 l_2 = +44; end
		36603: begin l_1 = +23;
				 l_2 = -44; end
		14258: begin l_1 = -23;
				 l_2 = +44; end
		40060: begin l_1 = -23;
				 l_2 = -44; end
		48761: begin l_1 = +23;
				 l_2 = +45; end
		49504: begin l_1 = +23;
				 l_2 = -45; end
		1357: begin l_1 = -23;
				 l_2 = +45; end
		2100: begin l_1 = -23;
				 l_2 = -45; end
		22959: begin l_1 = +23;
				 l_2 = +46; end
		24445: begin l_1 = +23;
				 l_2 = -46; end
		26416: begin l_1 = -23;
				 l_2 = +46; end
		27902: begin l_1 = -23;
				 l_2 = -46; end
		22216: begin l_1 = +23;
				 l_2 = +47; end
		25188: begin l_1 = +23;
				 l_2 = -47; end
		25673: begin l_1 = -23;
				 l_2 = +47; end
		28645: begin l_1 = -23;
				 l_2 = -47; end
		20730: begin l_1 = +23;
				 l_2 = +48; end
		26674: begin l_1 = +23;
				 l_2 = -48; end
		24187: begin l_1 = -23;
				 l_2 = +48; end
		30131: begin l_1 = -23;
				 l_2 = -48; end
		17758: begin l_1 = +23;
				 l_2 = +49; end
		29646: begin l_1 = +23;
				 l_2 = -49; end
		21215: begin l_1 = -23;
				 l_2 = +49; end
		33103: begin l_1 = -23;
				 l_2 = -49; end
		11814: begin l_1 = +23;
				 l_2 = +50; end
		35590: begin l_1 = +23;
				 l_2 = -50; end
		15271: begin l_1 = -23;
				 l_2 = +50; end
		39047: begin l_1 = -23;
				 l_2 = -50; end
		50787: begin l_1 = +23;
				 l_2 = +51; end
		47478: begin l_1 = +23;
				 l_2 = -51; end
		3383: begin l_1 = -23;
				 l_2 = +51; end
		74: begin l_1 = -23;
				 l_2 = -51; end
		27011: begin l_1 = +23;
				 l_2 = +52; end
		20393: begin l_1 = +23;
				 l_2 = -52; end
		30468: begin l_1 = -23;
				 l_2 = +52; end
		23850: begin l_1 = -23;
				 l_2 = -52; end
		30320: begin l_1 = +23;
				 l_2 = +53; end
		17084: begin l_1 = +23;
				 l_2 = -53; end
		33777: begin l_1 = -23;
				 l_2 = +53; end
		20541: begin l_1 = -23;
				 l_2 = -53; end
		36938: begin l_1 = +23;
				 l_2 = +54; end
		10466: begin l_1 = +23;
				 l_2 = -54; end
		40395: begin l_1 = -23;
				 l_2 = +54; end
		13923: begin l_1 = -23;
				 l_2 = -54; end
		50174: begin l_1 = +23;
				 l_2 = +55; end
		48091: begin l_1 = +23;
				 l_2 = -55; end
		2770: begin l_1 = -23;
				 l_2 = +55; end
		687: begin l_1 = -23;
				 l_2 = -55; end
		25785: begin l_1 = +23;
				 l_2 = +56; end
		21619: begin l_1 = +23;
				 l_2 = -56; end
		29242: begin l_1 = -23;
				 l_2 = +56; end
		25076: begin l_1 = -23;
				 l_2 = -56; end
		27868: begin l_1 = +23;
				 l_2 = +57; end
		19536: begin l_1 = +23;
				 l_2 = -57; end
		31325: begin l_1 = -23;
				 l_2 = +57; end
		22993: begin l_1 = -23;
				 l_2 = -57; end
		32034: begin l_1 = +23;
				 l_2 = +58; end
		15370: begin l_1 = +23;
				 l_2 = -58; end
		35491: begin l_1 = -23;
				 l_2 = +58; end
		18827: begin l_1 = -23;
				 l_2 = -58; end
		40366: begin l_1 = +23;
				 l_2 = +59; end
		7038: begin l_1 = +23;
				 l_2 = -59; end
		43823: begin l_1 = -23;
				 l_2 = +59; end
		10495: begin l_1 = -23;
				 l_2 = -59; end
		6169: begin l_1 = +23;
				 l_2 = +60; end
		41235: begin l_1 = +23;
				 l_2 = -60; end
		9626: begin l_1 = -23;
				 l_2 = +60; end
		44692: begin l_1 = -23;
				 l_2 = -60; end
		39497: begin l_1 = +23;
				 l_2 = +61; end
		7907: begin l_1 = +23;
				 l_2 = -61; end
		42954: begin l_1 = -23;
				 l_2 = +61; end
		11364: begin l_1 = -23;
				 l_2 = -61; end
		4431: begin l_1 = +23;
				 l_2 = +62; end
		42973: begin l_1 = +23;
				 l_2 = -62; end
		7888: begin l_1 = -23;
				 l_2 = +62; end
		46430: begin l_1 = -23;
				 l_2 = -62; end
		36021: begin l_1 = +23;
				 l_2 = +63; end
		11383: begin l_1 = +23;
				 l_2 = -63; end
		39478: begin l_1 = -23;
				 l_2 = +63; end
		14840: begin l_1 = -23;
				 l_2 = -63; end
		48340: begin l_1 = +23;
				 l_2 = +64; end
		49925: begin l_1 = +23;
				 l_2 = -64; end
		936: begin l_1 = -23;
				 l_2 = +64; end
		2521: begin l_1 = -23;
				 l_2 = -64; end
		22117: begin l_1 = +23;
				 l_2 = +65; end
		25287: begin l_1 = +23;
				 l_2 = -65; end
		25574: begin l_1 = -23;
				 l_2 = +65; end
		28744: begin l_1 = -23;
				 l_2 = -65; end
		20532: begin l_1 = +23;
				 l_2 = +66; end
		26872: begin l_1 = +23;
				 l_2 = -66; end
		23989: begin l_1 = -23;
				 l_2 = +66; end
		30329: begin l_1 = -23;
				 l_2 = -66; end
		17362: begin l_1 = +23;
				 l_2 = +67; end
		30042: begin l_1 = +23;
				 l_2 = -67; end
		20819: begin l_1 = -23;
				 l_2 = +67; end
		33499: begin l_1 = -23;
				 l_2 = -67; end
		11022: begin l_1 = +23;
				 l_2 = +68; end
		36382: begin l_1 = +23;
				 l_2 = -68; end
		14479: begin l_1 = -23;
				 l_2 = +68; end
		39839: begin l_1 = -23;
				 l_2 = -68; end
		40490: begin l_1 = -24;
				 l_2 = +26; end
		10371: begin l_1 = -24;
				 l_2 = -25; end
		33576: begin l_1 = +24;
				 l_2 = +26; end
		17285: begin l_1 = -24;
				 l_2 = -26; end
		19748: begin l_1 = +24;
				 l_2 = +27; end
		24199: begin l_1 = +24;
				 l_2 = -27; end
		26662: begin l_1 = -24;
				 l_2 = +27; end
		31113: begin l_1 = -24;
				 l_2 = -27; end
		42953: begin l_1 = +24;
				 l_2 = +28; end
		994: begin l_1 = +24;
				 l_2 = -28; end
		49867: begin l_1 = -24;
				 l_2 = +28; end
		7908: begin l_1 = -24;
				 l_2 = -28; end
		38502: begin l_1 = +24;
				 l_2 = +29; end
		5445: begin l_1 = +24;
				 l_2 = -29; end
		45416: begin l_1 = -24;
				 l_2 = +29; end
		12359: begin l_1 = -24;
				 l_2 = -29; end
		29600: begin l_1 = +24;
				 l_2 = +30; end
		14347: begin l_1 = +24;
				 l_2 = -30; end
		36514: begin l_1 = -24;
				 l_2 = +30; end
		21261: begin l_1 = -24;
				 l_2 = -30; end
		11796: begin l_1 = +24;
				 l_2 = +31; end
		32151: begin l_1 = +24;
				 l_2 = -31; end
		18710: begin l_1 = -24;
				 l_2 = +31; end
		39065: begin l_1 = -24;
				 l_2 = -31; end
		27049: begin l_1 = +24;
				 l_2 = +32; end
		16898: begin l_1 = +24;
				 l_2 = -32; end
		33963: begin l_1 = -24;
				 l_2 = +32; end
		23812: begin l_1 = -24;
				 l_2 = -32; end
		6694: begin l_1 = +24;
				 l_2 = +33; end
		37253: begin l_1 = +24;
				 l_2 = -33; end
		13608: begin l_1 = -24;
				 l_2 = +33; end
		44167: begin l_1 = -24;
				 l_2 = -33; end
		16845: begin l_1 = +24;
				 l_2 = +34; end
		27102: begin l_1 = +24;
				 l_2 = -34; end
		23759: begin l_1 = -24;
				 l_2 = +34; end
		34016: begin l_1 = -24;
				 l_2 = -34; end
		37147: begin l_1 = +24;
				 l_2 = +35; end
		6800: begin l_1 = +24;
				 l_2 = -35; end
		44061: begin l_1 = -24;
				 l_2 = +35; end
		13714: begin l_1 = -24;
				 l_2 = -35; end
		26890: begin l_1 = +24;
				 l_2 = +36; end
		17057: begin l_1 = +24;
				 l_2 = -36; end
		33804: begin l_1 = -24;
				 l_2 = +36; end
		23971: begin l_1 = -24;
				 l_2 = -36; end
		6376: begin l_1 = +24;
				 l_2 = +37; end
		37571: begin l_1 = +24;
				 l_2 = -37; end
		13290: begin l_1 = -24;
				 l_2 = +37; end
		44485: begin l_1 = -24;
				 l_2 = -37; end
		16209: begin l_1 = +24;
				 l_2 = +38; end
		27738: begin l_1 = +24;
				 l_2 = -38; end
		23123: begin l_1 = -24;
				 l_2 = +38; end
		34652: begin l_1 = -24;
				 l_2 = -38; end
		35875: begin l_1 = +24;
				 l_2 = +39; end
		8072: begin l_1 = +24;
				 l_2 = -39; end
		42789: begin l_1 = -24;
				 l_2 = +39; end
		14986: begin l_1 = -24;
				 l_2 = -39; end
		24346: begin l_1 = +24;
				 l_2 = +40; end
		19601: begin l_1 = +24;
				 l_2 = -40; end
		31260: begin l_1 = -24;
				 l_2 = +40; end
		26515: begin l_1 = -24;
				 l_2 = -40; end
		1288: begin l_1 = +24;
				 l_2 = +41; end
		42659: begin l_1 = +24;
				 l_2 = -41; end
		8202: begin l_1 = -24;
				 l_2 = +41; end
		49573: begin l_1 = -24;
				 l_2 = -41; end
		6033: begin l_1 = +24;
				 l_2 = +42; end
		37914: begin l_1 = +24;
				 l_2 = -42; end
		12947: begin l_1 = -24;
				 l_2 = +42; end
		44828: begin l_1 = -24;
				 l_2 = -42; end
		15523: begin l_1 = +24;
				 l_2 = +43; end
		28424: begin l_1 = +24;
				 l_2 = -43; end
		22437: begin l_1 = -24;
				 l_2 = +43; end
		35338: begin l_1 = -24;
				 l_2 = -43; end
		34503: begin l_1 = +24;
				 l_2 = +44; end
		9444: begin l_1 = +24;
				 l_2 = -44; end
		41417: begin l_1 = -24;
				 l_2 = +44; end
		16358: begin l_1 = -24;
				 l_2 = -44; end
		21602: begin l_1 = +24;
				 l_2 = +45; end
		22345: begin l_1 = +24;
				 l_2 = -45; end
		28516: begin l_1 = -24;
				 l_2 = +45; end
		29259: begin l_1 = -24;
				 l_2 = -45; end
		46661: begin l_1 = +24;
				 l_2 = +46; end
		48147: begin l_1 = +24;
				 l_2 = -46; end
		2714: begin l_1 = -24;
				 l_2 = +46; end
		4200: begin l_1 = -24;
				 l_2 = -46; end
		45918: begin l_1 = +24;
				 l_2 = +47; end
		48890: begin l_1 = +24;
				 l_2 = -47; end
		1971: begin l_1 = -24;
				 l_2 = +47; end
		4943: begin l_1 = -24;
				 l_2 = -47; end
		44432: begin l_1 = +24;
				 l_2 = +48; end
		50376: begin l_1 = +24;
				 l_2 = -48; end
		485: begin l_1 = -24;
				 l_2 = +48; end
		6429: begin l_1 = -24;
				 l_2 = -48; end
		41460: begin l_1 = +24;
				 l_2 = +49; end
		2487: begin l_1 = +24;
				 l_2 = -49; end
		48374: begin l_1 = -24;
				 l_2 = +49; end
		9401: begin l_1 = -24;
				 l_2 = -49; end
		35516: begin l_1 = +24;
				 l_2 = +50; end
		8431: begin l_1 = +24;
				 l_2 = -50; end
		42430: begin l_1 = -24;
				 l_2 = +50; end
		15345: begin l_1 = -24;
				 l_2 = -50; end
		23628: begin l_1 = +24;
				 l_2 = +51; end
		20319: begin l_1 = +24;
				 l_2 = -51; end
		30542: begin l_1 = -24;
				 l_2 = +51; end
		27233: begin l_1 = -24;
				 l_2 = -51; end
		50713: begin l_1 = +24;
				 l_2 = +52; end
		44095: begin l_1 = +24;
				 l_2 = -52; end
		6766: begin l_1 = -24;
				 l_2 = +52; end
		148: begin l_1 = -24;
				 l_2 = -52; end
		3161: begin l_1 = +24;
				 l_2 = +53; end
		40786: begin l_1 = +24;
				 l_2 = -53; end
		10075: begin l_1 = -24;
				 l_2 = +53; end
		47700: begin l_1 = -24;
				 l_2 = -53; end
		9779: begin l_1 = +24;
				 l_2 = +54; end
		34168: begin l_1 = +24;
				 l_2 = -54; end
		16693: begin l_1 = -24;
				 l_2 = +54; end
		41082: begin l_1 = -24;
				 l_2 = -54; end
		23015: begin l_1 = +24;
				 l_2 = +55; end
		20932: begin l_1 = +24;
				 l_2 = -55; end
		29929: begin l_1 = -24;
				 l_2 = +55; end
		27846: begin l_1 = -24;
				 l_2 = -55; end
		49487: begin l_1 = +24;
				 l_2 = +56; end
		45321: begin l_1 = +24;
				 l_2 = -56; end
		5540: begin l_1 = -24;
				 l_2 = +56; end
		1374: begin l_1 = -24;
				 l_2 = -56; end
		709: begin l_1 = +24;
				 l_2 = +57; end
		43238: begin l_1 = +24;
				 l_2 = -57; end
		7623: begin l_1 = -24;
				 l_2 = +57; end
		50152: begin l_1 = -24;
				 l_2 = -57; end
		4875: begin l_1 = +24;
				 l_2 = +58; end
		39072: begin l_1 = +24;
				 l_2 = -58; end
		11789: begin l_1 = -24;
				 l_2 = +58; end
		45986: begin l_1 = -24;
				 l_2 = -58; end
		13207: begin l_1 = +24;
				 l_2 = +59; end
		30740: begin l_1 = +24;
				 l_2 = -59; end
		20121: begin l_1 = -24;
				 l_2 = +59; end
		37654: begin l_1 = -24;
				 l_2 = -59; end
		29871: begin l_1 = +24;
				 l_2 = +60; end
		14076: begin l_1 = +24;
				 l_2 = -60; end
		36785: begin l_1 = -24;
				 l_2 = +60; end
		20990: begin l_1 = -24;
				 l_2 = -60; end
		12338: begin l_1 = +24;
				 l_2 = +61; end
		31609: begin l_1 = +24;
				 l_2 = -61; end
		19252: begin l_1 = -24;
				 l_2 = +61; end
		38523: begin l_1 = -24;
				 l_2 = -61; end
		28133: begin l_1 = +24;
				 l_2 = +62; end
		15814: begin l_1 = +24;
				 l_2 = -62; end
		35047: begin l_1 = -24;
				 l_2 = +62; end
		22728: begin l_1 = -24;
				 l_2 = -62; end
		8862: begin l_1 = +24;
				 l_2 = +63; end
		35085: begin l_1 = +24;
				 l_2 = -63; end
		15776: begin l_1 = -24;
				 l_2 = +63; end
		41999: begin l_1 = -24;
				 l_2 = -63; end
		21181: begin l_1 = +24;
				 l_2 = +64; end
		22766: begin l_1 = +24;
				 l_2 = -64; end
		28095: begin l_1 = -24;
				 l_2 = +64; end
		29680: begin l_1 = -24;
				 l_2 = -64; end
		45819: begin l_1 = +24;
				 l_2 = +65; end
		48989: begin l_1 = +24;
				 l_2 = -65; end
		1872: begin l_1 = -24;
				 l_2 = +65; end
		5042: begin l_1 = -24;
				 l_2 = -65; end
		44234: begin l_1 = +24;
				 l_2 = +66; end
		50574: begin l_1 = +24;
				 l_2 = -66; end
		287: begin l_1 = -24;
				 l_2 = +66; end
		6627: begin l_1 = -24;
				 l_2 = -66; end
		41064: begin l_1 = +24;
				 l_2 = +67; end
		2883: begin l_1 = +24;
				 l_2 = -67; end
		47978: begin l_1 = -24;
				 l_2 = +67; end
		9797: begin l_1 = -24;
				 l_2 = -67; end
		34724: begin l_1 = +24;
				 l_2 = +68; end
		9223: begin l_1 = +24;
				 l_2 = -68; end
		41638: begin l_1 = -24;
				 l_2 = +68; end
		16137: begin l_1 = -24;
				 l_2 = -68; end
		30119: begin l_1 = -25;
				 l_2 = +27; end
		20742: begin l_1 = -25;
				 l_2 = -26; end
		16291: begin l_1 = +25;
				 l_2 = +27; end
		34570: begin l_1 = -25;
				 l_2 = -27; end
		39496: begin l_1 = +25;
				 l_2 = +28; end
		48398: begin l_1 = +25;
				 l_2 = -28; end
		2463: begin l_1 = -25;
				 l_2 = +28; end
		11365: begin l_1 = -25;
				 l_2 = -28; end
		35045: begin l_1 = +25;
				 l_2 = +29; end
		1988: begin l_1 = +25;
				 l_2 = -29; end
		48873: begin l_1 = -25;
				 l_2 = +29; end
		15816: begin l_1 = -25;
				 l_2 = -29; end
		26143: begin l_1 = +25;
				 l_2 = +30; end
		10890: begin l_1 = +25;
				 l_2 = -30; end
		39971: begin l_1 = -25;
				 l_2 = +30; end
		24718: begin l_1 = -25;
				 l_2 = -30; end
		8339: begin l_1 = +25;
				 l_2 = +31; end
		28694: begin l_1 = +25;
				 l_2 = -31; end
		22167: begin l_1 = -25;
				 l_2 = +31; end
		42522: begin l_1 = -25;
				 l_2 = -31; end
		23592: begin l_1 = +25;
				 l_2 = +32; end
		13441: begin l_1 = +25;
				 l_2 = -32; end
		37420: begin l_1 = -25;
				 l_2 = +32; end
		27269: begin l_1 = -25;
				 l_2 = -32; end
		3237: begin l_1 = +25;
				 l_2 = +33; end
		33796: begin l_1 = +25;
				 l_2 = -33; end
		17065: begin l_1 = -25;
				 l_2 = +33; end
		47624: begin l_1 = -25;
				 l_2 = -33; end
		13388: begin l_1 = +25;
				 l_2 = +34; end
		23645: begin l_1 = +25;
				 l_2 = -34; end
		27216: begin l_1 = -25;
				 l_2 = +34; end
		37473: begin l_1 = -25;
				 l_2 = -34; end
		33690: begin l_1 = +25;
				 l_2 = +35; end
		3343: begin l_1 = +25;
				 l_2 = -35; end
		47518: begin l_1 = -25;
				 l_2 = +35; end
		17171: begin l_1 = -25;
				 l_2 = -35; end
		23433: begin l_1 = +25;
				 l_2 = +36; end
		13600: begin l_1 = +25;
				 l_2 = -36; end
		37261: begin l_1 = -25;
				 l_2 = +36; end
		27428: begin l_1 = -25;
				 l_2 = -36; end
		2919: begin l_1 = +25;
				 l_2 = +37; end
		34114: begin l_1 = +25;
				 l_2 = -37; end
		16747: begin l_1 = -25;
				 l_2 = +37; end
		47942: begin l_1 = -25;
				 l_2 = -37; end
		12752: begin l_1 = +25;
				 l_2 = +38; end
		24281: begin l_1 = +25;
				 l_2 = -38; end
		26580: begin l_1 = -25;
				 l_2 = +38; end
		38109: begin l_1 = -25;
				 l_2 = -38; end
		32418: begin l_1 = +25;
				 l_2 = +39; end
		4615: begin l_1 = +25;
				 l_2 = -39; end
		46246: begin l_1 = -25;
				 l_2 = +39; end
		18443: begin l_1 = -25;
				 l_2 = -39; end
		20889: begin l_1 = +25;
				 l_2 = +40; end
		16144: begin l_1 = +25;
				 l_2 = -40; end
		34717: begin l_1 = -25;
				 l_2 = +40; end
		29972: begin l_1 = -25;
				 l_2 = -40; end
		48692: begin l_1 = +25;
				 l_2 = +41; end
		39202: begin l_1 = +25;
				 l_2 = -41; end
		11659: begin l_1 = -25;
				 l_2 = +41; end
		2169: begin l_1 = -25;
				 l_2 = -41; end
		2576: begin l_1 = +25;
				 l_2 = +42; end
		34457: begin l_1 = +25;
				 l_2 = -42; end
		16404: begin l_1 = -25;
				 l_2 = +42; end
		48285: begin l_1 = -25;
				 l_2 = -42; end
		12066: begin l_1 = +25;
				 l_2 = +43; end
		24967: begin l_1 = +25;
				 l_2 = -43; end
		25894: begin l_1 = -25;
				 l_2 = +43; end
		38795: begin l_1 = -25;
				 l_2 = -43; end
		31046: begin l_1 = +25;
				 l_2 = +44; end
		5987: begin l_1 = +25;
				 l_2 = -44; end
		44874: begin l_1 = -25;
				 l_2 = +44; end
		19815: begin l_1 = -25;
				 l_2 = -44; end
		18145: begin l_1 = +25;
				 l_2 = +45; end
		18888: begin l_1 = +25;
				 l_2 = -45; end
		31973: begin l_1 = -25;
				 l_2 = +45; end
		32716: begin l_1 = -25;
				 l_2 = -45; end
		43204: begin l_1 = +25;
				 l_2 = +46; end
		44690: begin l_1 = +25;
				 l_2 = -46; end
		6171: begin l_1 = -25;
				 l_2 = +46; end
		7657: begin l_1 = -25;
				 l_2 = -46; end
		42461: begin l_1 = +25;
				 l_2 = +47; end
		45433: begin l_1 = +25;
				 l_2 = -47; end
		5428: begin l_1 = -25;
				 l_2 = +47; end
		8400: begin l_1 = -25;
				 l_2 = -47; end
		40975: begin l_1 = +25;
				 l_2 = +48; end
		46919: begin l_1 = +25;
				 l_2 = -48; end
		3942: begin l_1 = -25;
				 l_2 = +48; end
		9886: begin l_1 = -25;
				 l_2 = -48; end
		38003: begin l_1 = +25;
				 l_2 = +49; end
		49891: begin l_1 = +25;
				 l_2 = -49; end
		970: begin l_1 = -25;
				 l_2 = +49; end
		12858: begin l_1 = -25;
				 l_2 = -49; end
		32059: begin l_1 = +25;
				 l_2 = +50; end
		4974: begin l_1 = +25;
				 l_2 = -50; end
		45887: begin l_1 = -25;
				 l_2 = +50; end
		18802: begin l_1 = -25;
				 l_2 = -50; end
		20171: begin l_1 = +25;
				 l_2 = +51; end
		16862: begin l_1 = +25;
				 l_2 = -51; end
		33999: begin l_1 = -25;
				 l_2 = +51; end
		30690: begin l_1 = -25;
				 l_2 = -51; end
		47256: begin l_1 = +25;
				 l_2 = +52; end
		40638: begin l_1 = +25;
				 l_2 = -52; end
		10223: begin l_1 = -25;
				 l_2 = +52; end
		3605: begin l_1 = -25;
				 l_2 = -52; end
		50565: begin l_1 = +25;
				 l_2 = +53; end
		37329: begin l_1 = +25;
				 l_2 = -53; end
		13532: begin l_1 = -25;
				 l_2 = +53; end
		296: begin l_1 = -25;
				 l_2 = -53; end
		6322: begin l_1 = +25;
				 l_2 = +54; end
		30711: begin l_1 = +25;
				 l_2 = -54; end
		20150: begin l_1 = -25;
				 l_2 = +54; end
		44539: begin l_1 = -25;
				 l_2 = -54; end
		19558: begin l_1 = +25;
				 l_2 = +55; end
		17475: begin l_1 = +25;
				 l_2 = -55; end
		33386: begin l_1 = -25;
				 l_2 = +55; end
		31303: begin l_1 = -25;
				 l_2 = -55; end
		46030: begin l_1 = +25;
				 l_2 = +56; end
		41864: begin l_1 = +25;
				 l_2 = -56; end
		8997: begin l_1 = -25;
				 l_2 = +56; end
		4831: begin l_1 = -25;
				 l_2 = -56; end
		48113: begin l_1 = +25;
				 l_2 = +57; end
		39781: begin l_1 = +25;
				 l_2 = -57; end
		11080: begin l_1 = -25;
				 l_2 = +57; end
		2748: begin l_1 = -25;
				 l_2 = -57; end
		1418: begin l_1 = +25;
				 l_2 = +58; end
		35615: begin l_1 = +25;
				 l_2 = -58; end
		15246: begin l_1 = -25;
				 l_2 = +58; end
		49443: begin l_1 = -25;
				 l_2 = -58; end
		9750: begin l_1 = +25;
				 l_2 = +59; end
		27283: begin l_1 = +25;
				 l_2 = -59; end
		23578: begin l_1 = -25;
				 l_2 = +59; end
		41111: begin l_1 = -25;
				 l_2 = -59; end
		26414: begin l_1 = +25;
				 l_2 = +60; end
		10619: begin l_1 = +25;
				 l_2 = -60; end
		40242: begin l_1 = -25;
				 l_2 = +60; end
		24447: begin l_1 = -25;
				 l_2 = -60; end
		8881: begin l_1 = +25;
				 l_2 = +61; end
		28152: begin l_1 = +25;
				 l_2 = -61; end
		22709: begin l_1 = -25;
				 l_2 = +61; end
		41980: begin l_1 = -25;
				 l_2 = -61; end
		24676: begin l_1 = +25;
				 l_2 = +62; end
		12357: begin l_1 = +25;
				 l_2 = -62; end
		38504: begin l_1 = -25;
				 l_2 = +62; end
		26185: begin l_1 = -25;
				 l_2 = -62; end
		5405: begin l_1 = +25;
				 l_2 = +63; end
		31628: begin l_1 = +25;
				 l_2 = -63; end
		19233: begin l_1 = -25;
				 l_2 = +63; end
		45456: begin l_1 = -25;
				 l_2 = -63; end
		17724: begin l_1 = +25;
				 l_2 = +64; end
		19309: begin l_1 = +25;
				 l_2 = -64; end
		31552: begin l_1 = -25;
				 l_2 = +64; end
		33137: begin l_1 = -25;
				 l_2 = -64; end
		42362: begin l_1 = +25;
				 l_2 = +65; end
		45532: begin l_1 = +25;
				 l_2 = -65; end
		5329: begin l_1 = -25;
				 l_2 = +65; end
		8499: begin l_1 = -25;
				 l_2 = -65; end
		40777: begin l_1 = +25;
				 l_2 = +66; end
		47117: begin l_1 = +25;
				 l_2 = -66; end
		3744: begin l_1 = -25;
				 l_2 = +66; end
		10084: begin l_1 = -25;
				 l_2 = -66; end
		37607: begin l_1 = +25;
				 l_2 = +67; end
		50287: begin l_1 = +25;
				 l_2 = -67; end
		574: begin l_1 = -25;
				 l_2 = +67; end
		13254: begin l_1 = -25;
				 l_2 = -67; end
		31267: begin l_1 = +25;
				 l_2 = +68; end
		5766: begin l_1 = +25;
				 l_2 = -68; end
		45095: begin l_1 = -25;
				 l_2 = +68; end
		19594: begin l_1 = -25;
				 l_2 = -68; end
		9377: begin l_1 = -26;
				 l_2 = +28; end
		41484: begin l_1 = -26;
				 l_2 = -27; end
		32582: begin l_1 = +26;
				 l_2 = +28; end
		18279: begin l_1 = -26;
				 l_2 = -28; end
		28131: begin l_1 = +26;
				 l_2 = +29; end
		45935: begin l_1 = +26;
				 l_2 = -29; end
		4926: begin l_1 = -26;
				 l_2 = +29; end
		22730: begin l_1 = -26;
				 l_2 = -29; end
		19229: begin l_1 = +26;
				 l_2 = +30; end
		3976: begin l_1 = +26;
				 l_2 = -30; end
		46885: begin l_1 = -26;
				 l_2 = +30; end
		31632: begin l_1 = -26;
				 l_2 = -30; end
		1425: begin l_1 = +26;
				 l_2 = +31; end
		21780: begin l_1 = +26;
				 l_2 = -31; end
		29081: begin l_1 = -26;
				 l_2 = +31; end
		49436: begin l_1 = -26;
				 l_2 = -31; end
		16678: begin l_1 = +26;
				 l_2 = +32; end
		6527: begin l_1 = +26;
				 l_2 = -32; end
		44334: begin l_1 = -26;
				 l_2 = +32; end
		34183: begin l_1 = -26;
				 l_2 = -32; end
		47184: begin l_1 = +26;
				 l_2 = +33; end
		26882: begin l_1 = +26;
				 l_2 = -33; end
		23979: begin l_1 = -26;
				 l_2 = +33; end
		3677: begin l_1 = -26;
				 l_2 = -33; end
		6474: begin l_1 = +26;
				 l_2 = +34; end
		16731: begin l_1 = +26;
				 l_2 = -34; end
		34130: begin l_1 = -26;
				 l_2 = +34; end
		44387: begin l_1 = -26;
				 l_2 = -34; end
		26776: begin l_1 = +26;
				 l_2 = +35; end
		47290: begin l_1 = +26;
				 l_2 = -35; end
		3571: begin l_1 = -26;
				 l_2 = +35; end
		24085: begin l_1 = -26;
				 l_2 = -35; end
		16519: begin l_1 = +26;
				 l_2 = +36; end
		6686: begin l_1 = +26;
				 l_2 = -36; end
		44175: begin l_1 = -26;
				 l_2 = +36; end
		34342: begin l_1 = -26;
				 l_2 = -36; end
		46866: begin l_1 = +26;
				 l_2 = +37; end
		27200: begin l_1 = +26;
				 l_2 = -37; end
		23661: begin l_1 = -26;
				 l_2 = +37; end
		3995: begin l_1 = -26;
				 l_2 = -37; end
		5838: begin l_1 = +26;
				 l_2 = +38; end
		17367: begin l_1 = +26;
				 l_2 = -38; end
		33494: begin l_1 = -26;
				 l_2 = +38; end
		45023: begin l_1 = -26;
				 l_2 = -38; end
		25504: begin l_1 = +26;
				 l_2 = +39; end
		48562: begin l_1 = +26;
				 l_2 = -39; end
		2299: begin l_1 = -26;
				 l_2 = +39; end
		25357: begin l_1 = -26;
				 l_2 = -39; end
		13975: begin l_1 = +26;
				 l_2 = +40; end
		9230: begin l_1 = +26;
				 l_2 = -40; end
		41631: begin l_1 = -26;
				 l_2 = +40; end
		36886: begin l_1 = -26;
				 l_2 = -40; end
		41778: begin l_1 = +26;
				 l_2 = +41; end
		32288: begin l_1 = +26;
				 l_2 = -41; end
		18573: begin l_1 = -26;
				 l_2 = +41; end
		9083: begin l_1 = -26;
				 l_2 = -41; end
		46523: begin l_1 = +26;
				 l_2 = +42; end
		27543: begin l_1 = +26;
				 l_2 = -42; end
		23318: begin l_1 = -26;
				 l_2 = +42; end
		4338: begin l_1 = -26;
				 l_2 = -42; end
		5152: begin l_1 = +26;
				 l_2 = +43; end
		18053: begin l_1 = +26;
				 l_2 = -43; end
		32808: begin l_1 = -26;
				 l_2 = +43; end
		45709: begin l_1 = -26;
				 l_2 = -43; end
		24132: begin l_1 = +26;
				 l_2 = +44; end
		49934: begin l_1 = +26;
				 l_2 = -44; end
		927: begin l_1 = -26;
				 l_2 = +44; end
		26729: begin l_1 = -26;
				 l_2 = -44; end
		11231: begin l_1 = +26;
				 l_2 = +45; end
		11974: begin l_1 = +26;
				 l_2 = -45; end
		38887: begin l_1 = -26;
				 l_2 = +45; end
		39630: begin l_1 = -26;
				 l_2 = -45; end
		36290: begin l_1 = +26;
				 l_2 = +46; end
		37776: begin l_1 = +26;
				 l_2 = -46; end
		13085: begin l_1 = -26;
				 l_2 = +46; end
		14571: begin l_1 = -26;
				 l_2 = -46; end
		35547: begin l_1 = +26;
				 l_2 = +47; end
		38519: begin l_1 = +26;
				 l_2 = -47; end
		12342: begin l_1 = -26;
				 l_2 = +47; end
		15314: begin l_1 = -26;
				 l_2 = -47; end
		34061: begin l_1 = +26;
				 l_2 = +48; end
		40005: begin l_1 = +26;
				 l_2 = -48; end
		10856: begin l_1 = -26;
				 l_2 = +48; end
		16800: begin l_1 = -26;
				 l_2 = -48; end
		31089: begin l_1 = +26;
				 l_2 = +49; end
		42977: begin l_1 = +26;
				 l_2 = -49; end
		7884: begin l_1 = -26;
				 l_2 = +49; end
		19772: begin l_1 = -26;
				 l_2 = -49; end
		25145: begin l_1 = +26;
				 l_2 = +50; end
		48921: begin l_1 = +26;
				 l_2 = -50; end
		1940: begin l_1 = -26;
				 l_2 = +50; end
		25716: begin l_1 = -26;
				 l_2 = -50; end
		13257: begin l_1 = +26;
				 l_2 = +51; end
		9948: begin l_1 = +26;
				 l_2 = -51; end
		40913: begin l_1 = -26;
				 l_2 = +51; end
		37604: begin l_1 = -26;
				 l_2 = -51; end
		40342: begin l_1 = +26;
				 l_2 = +52; end
		33724: begin l_1 = +26;
				 l_2 = -52; end
		17137: begin l_1 = -26;
				 l_2 = +52; end
		10519: begin l_1 = -26;
				 l_2 = -52; end
		43651: begin l_1 = +26;
				 l_2 = +53; end
		30415: begin l_1 = +26;
				 l_2 = -53; end
		20446: begin l_1 = -26;
				 l_2 = +53; end
		7210: begin l_1 = -26;
				 l_2 = -53; end
		50269: begin l_1 = +26;
				 l_2 = +54; end
		23797: begin l_1 = +26;
				 l_2 = -54; end
		27064: begin l_1 = -26;
				 l_2 = +54; end
		592: begin l_1 = -26;
				 l_2 = -54; end
		12644: begin l_1 = +26;
				 l_2 = +55; end
		10561: begin l_1 = +26;
				 l_2 = -55; end
		40300: begin l_1 = -26;
				 l_2 = +55; end
		38217: begin l_1 = -26;
				 l_2 = -55; end
		39116: begin l_1 = +26;
				 l_2 = +56; end
		34950: begin l_1 = +26;
				 l_2 = -56; end
		15911: begin l_1 = -26;
				 l_2 = +56; end
		11745: begin l_1 = -26;
				 l_2 = -56; end
		41199: begin l_1 = +26;
				 l_2 = +57; end
		32867: begin l_1 = +26;
				 l_2 = -57; end
		17994: begin l_1 = -26;
				 l_2 = +57; end
		9662: begin l_1 = -26;
				 l_2 = -57; end
		45365: begin l_1 = +26;
				 l_2 = +58; end
		28701: begin l_1 = +26;
				 l_2 = -58; end
		22160: begin l_1 = -26;
				 l_2 = +58; end
		5496: begin l_1 = -26;
				 l_2 = -58; end
		2836: begin l_1 = +26;
				 l_2 = +59; end
		20369: begin l_1 = +26;
				 l_2 = -59; end
		30492: begin l_1 = -26;
				 l_2 = +59; end
		48025: begin l_1 = -26;
				 l_2 = -59; end
		19500: begin l_1 = +26;
				 l_2 = +60; end
		3705: begin l_1 = +26;
				 l_2 = -60; end
		47156: begin l_1 = -26;
				 l_2 = +60; end
		31361: begin l_1 = -26;
				 l_2 = -60; end
		1967: begin l_1 = +26;
				 l_2 = +61; end
		21238: begin l_1 = +26;
				 l_2 = -61; end
		29623: begin l_1 = -26;
				 l_2 = +61; end
		48894: begin l_1 = -26;
				 l_2 = -61; end
		17762: begin l_1 = +26;
				 l_2 = +62; end
		5443: begin l_1 = +26;
				 l_2 = -62; end
		45418: begin l_1 = -26;
				 l_2 = +62; end
		33099: begin l_1 = -26;
				 l_2 = -62; end
		49352: begin l_1 = +26;
				 l_2 = +63; end
		24714: begin l_1 = +26;
				 l_2 = -63; end
		26147: begin l_1 = -26;
				 l_2 = +63; end
		1509: begin l_1 = -26;
				 l_2 = -63; end
		10810: begin l_1 = +26;
				 l_2 = +64; end
		12395: begin l_1 = +26;
				 l_2 = -64; end
		38466: begin l_1 = -26;
				 l_2 = +64; end
		40051: begin l_1 = -26;
				 l_2 = -64; end
		35448: begin l_1 = +26;
				 l_2 = +65; end
		38618: begin l_1 = +26;
				 l_2 = -65; end
		12243: begin l_1 = -26;
				 l_2 = +65; end
		15413: begin l_1 = -26;
				 l_2 = -65; end
		33863: begin l_1 = +26;
				 l_2 = +66; end
		40203: begin l_1 = +26;
				 l_2 = -66; end
		10658: begin l_1 = -26;
				 l_2 = +66; end
		16998: begin l_1 = -26;
				 l_2 = -66; end
		30693: begin l_1 = +26;
				 l_2 = +67; end
		43373: begin l_1 = +26;
				 l_2 = -67; end
		7488: begin l_1 = -26;
				 l_2 = +67; end
		20168: begin l_1 = -26;
				 l_2 = -67; end
		24353: begin l_1 = +26;
				 l_2 = +68; end
		49713: begin l_1 = +26;
				 l_2 = -68; end
		1148: begin l_1 = -26;
				 l_2 = +68; end
		26508: begin l_1 = -26;
				 l_2 = -68; end
		18754: begin l_1 = -27;
				 l_2 = +29; end
		32107: begin l_1 = -27;
				 l_2 = -28; end
		14303: begin l_1 = +27;
				 l_2 = +29; end
		36558: begin l_1 = -27;
				 l_2 = -29; end
		5401: begin l_1 = +27;
				 l_2 = +30; end
		41009: begin l_1 = +27;
				 l_2 = -30; end
		9852: begin l_1 = -27;
				 l_2 = +30; end
		45460: begin l_1 = -27;
				 l_2 = -30; end
		38458: begin l_1 = +27;
				 l_2 = +31; end
		7952: begin l_1 = +27;
				 l_2 = -31; end
		42909: begin l_1 = -27;
				 l_2 = +31; end
		12403: begin l_1 = -27;
				 l_2 = -31; end
		2850: begin l_1 = +27;
				 l_2 = +32; end
		43560: begin l_1 = +27;
				 l_2 = -32; end
		7301: begin l_1 = -27;
				 l_2 = +32; end
		48011: begin l_1 = -27;
				 l_2 = -32; end
		33356: begin l_1 = +27;
				 l_2 = +33; end
		13054: begin l_1 = +27;
				 l_2 = -33; end
		37807: begin l_1 = -27;
				 l_2 = +33; end
		17505: begin l_1 = -27;
				 l_2 = -33; end
		43507: begin l_1 = +27;
				 l_2 = +34; end
		2903: begin l_1 = +27;
				 l_2 = -34; end
		47958: begin l_1 = -27;
				 l_2 = +34; end
		7354: begin l_1 = -27;
				 l_2 = -34; end
		12948: begin l_1 = +27;
				 l_2 = +35; end
		33462: begin l_1 = +27;
				 l_2 = -35; end
		17399: begin l_1 = -27;
				 l_2 = +35; end
		37913: begin l_1 = -27;
				 l_2 = -35; end
		2691: begin l_1 = +27;
				 l_2 = +36; end
		43719: begin l_1 = +27;
				 l_2 = -36; end
		7142: begin l_1 = -27;
				 l_2 = +36; end
		48170: begin l_1 = -27;
				 l_2 = -36; end
		33038: begin l_1 = +27;
				 l_2 = +37; end
		13372: begin l_1 = +27;
				 l_2 = -37; end
		37489: begin l_1 = -27;
				 l_2 = +37; end
		17823: begin l_1 = -27;
				 l_2 = -37; end
		42871: begin l_1 = +27;
				 l_2 = +38; end
		3539: begin l_1 = +27;
				 l_2 = -38; end
		47322: begin l_1 = -27;
				 l_2 = +38; end
		7990: begin l_1 = -27;
				 l_2 = -38; end
		11676: begin l_1 = +27;
				 l_2 = +39; end
		34734: begin l_1 = +27;
				 l_2 = -39; end
		16127: begin l_1 = -27;
				 l_2 = +39; end
		39185: begin l_1 = -27;
				 l_2 = -39; end
		147: begin l_1 = +27;
				 l_2 = +40; end
		46263: begin l_1 = +27;
				 l_2 = -40; end
		4598: begin l_1 = -27;
				 l_2 = +40; end
		50714: begin l_1 = -27;
				 l_2 = -40; end
		27950: begin l_1 = +27;
				 l_2 = +41; end
		18460: begin l_1 = +27;
				 l_2 = -41; end
		32401: begin l_1 = -27;
				 l_2 = +41; end
		22911: begin l_1 = -27;
				 l_2 = -41; end
		32695: begin l_1 = +27;
				 l_2 = +42; end
		13715: begin l_1 = +27;
				 l_2 = -42; end
		37146: begin l_1 = -27;
				 l_2 = +42; end
		18166: begin l_1 = -27;
				 l_2 = -42; end
		42185: begin l_1 = +27;
				 l_2 = +43; end
		4225: begin l_1 = +27;
				 l_2 = -43; end
		46636: begin l_1 = -27;
				 l_2 = +43; end
		8676: begin l_1 = -27;
				 l_2 = -43; end
		10304: begin l_1 = +27;
				 l_2 = +44; end
		36106: begin l_1 = +27;
				 l_2 = -44; end
		14755: begin l_1 = -27;
				 l_2 = +44; end
		40557: begin l_1 = -27;
				 l_2 = -44; end
		48264: begin l_1 = +27;
				 l_2 = +45; end
		49007: begin l_1 = +27;
				 l_2 = -45; end
		1854: begin l_1 = -27;
				 l_2 = +45; end
		2597: begin l_1 = -27;
				 l_2 = -45; end
		22462: begin l_1 = +27;
				 l_2 = +46; end
		23948: begin l_1 = +27;
				 l_2 = -46; end
		26913: begin l_1 = -27;
				 l_2 = +46; end
		28399: begin l_1 = -27;
				 l_2 = -46; end
		21719: begin l_1 = +27;
				 l_2 = +47; end
		24691: begin l_1 = +27;
				 l_2 = -47; end
		26170: begin l_1 = -27;
				 l_2 = +47; end
		29142: begin l_1 = -27;
				 l_2 = -47; end
		20233: begin l_1 = +27;
				 l_2 = +48; end
		26177: begin l_1 = +27;
				 l_2 = -48; end
		24684: begin l_1 = -27;
				 l_2 = +48; end
		30628: begin l_1 = -27;
				 l_2 = -48; end
		17261: begin l_1 = +27;
				 l_2 = +49; end
		29149: begin l_1 = +27;
				 l_2 = -49; end
		21712: begin l_1 = -27;
				 l_2 = +49; end
		33600: begin l_1 = -27;
				 l_2 = -49; end
		11317: begin l_1 = +27;
				 l_2 = +50; end
		35093: begin l_1 = +27;
				 l_2 = -50; end
		15768: begin l_1 = -27;
				 l_2 = +50; end
		39544: begin l_1 = -27;
				 l_2 = -50; end
		50290: begin l_1 = +27;
				 l_2 = +51; end
		46981: begin l_1 = +27;
				 l_2 = -51; end
		3880: begin l_1 = -27;
				 l_2 = +51; end
		571: begin l_1 = -27;
				 l_2 = -51; end
		26514: begin l_1 = +27;
				 l_2 = +52; end
		19896: begin l_1 = +27;
				 l_2 = -52; end
		30965: begin l_1 = -27;
				 l_2 = +52; end
		24347: begin l_1 = -27;
				 l_2 = -52; end
		29823: begin l_1 = +27;
				 l_2 = +53; end
		16587: begin l_1 = +27;
				 l_2 = -53; end
		34274: begin l_1 = -27;
				 l_2 = +53; end
		21038: begin l_1 = -27;
				 l_2 = -53; end
		36441: begin l_1 = +27;
				 l_2 = +54; end
		9969: begin l_1 = +27;
				 l_2 = -54; end
		40892: begin l_1 = -27;
				 l_2 = +54; end
		14420: begin l_1 = -27;
				 l_2 = -54; end
		49677: begin l_1 = +27;
				 l_2 = +55; end
		47594: begin l_1 = +27;
				 l_2 = -55; end
		3267: begin l_1 = -27;
				 l_2 = +55; end
		1184: begin l_1 = -27;
				 l_2 = -55; end
		25288: begin l_1 = +27;
				 l_2 = +56; end
		21122: begin l_1 = +27;
				 l_2 = -56; end
		29739: begin l_1 = -27;
				 l_2 = +56; end
		25573: begin l_1 = -27;
				 l_2 = -56; end
		27371: begin l_1 = +27;
				 l_2 = +57; end
		19039: begin l_1 = +27;
				 l_2 = -57; end
		31822: begin l_1 = -27;
				 l_2 = +57; end
		23490: begin l_1 = -27;
				 l_2 = -57; end
		31537: begin l_1 = +27;
				 l_2 = +58; end
		14873: begin l_1 = +27;
				 l_2 = -58; end
		35988: begin l_1 = -27;
				 l_2 = +58; end
		19324: begin l_1 = -27;
				 l_2 = -58; end
		39869: begin l_1 = +27;
				 l_2 = +59; end
		6541: begin l_1 = +27;
				 l_2 = -59; end
		44320: begin l_1 = -27;
				 l_2 = +59; end
		10992: begin l_1 = -27;
				 l_2 = -59; end
		5672: begin l_1 = +27;
				 l_2 = +60; end
		40738: begin l_1 = +27;
				 l_2 = -60; end
		10123: begin l_1 = -27;
				 l_2 = +60; end
		45189: begin l_1 = -27;
				 l_2 = -60; end
		39000: begin l_1 = +27;
				 l_2 = +61; end
		7410: begin l_1 = +27;
				 l_2 = -61; end
		43451: begin l_1 = -27;
				 l_2 = +61; end
		11861: begin l_1 = -27;
				 l_2 = -61; end
		3934: begin l_1 = +27;
				 l_2 = +62; end
		42476: begin l_1 = +27;
				 l_2 = -62; end
		8385: begin l_1 = -27;
				 l_2 = +62; end
		46927: begin l_1 = -27;
				 l_2 = -62; end
		35524: begin l_1 = +27;
				 l_2 = +63; end
		10886: begin l_1 = +27;
				 l_2 = -63; end
		39975: begin l_1 = -27;
				 l_2 = +63; end
		15337: begin l_1 = -27;
				 l_2 = -63; end
		47843: begin l_1 = +27;
				 l_2 = +64; end
		49428: begin l_1 = +27;
				 l_2 = -64; end
		1433: begin l_1 = -27;
				 l_2 = +64; end
		3018: begin l_1 = -27;
				 l_2 = -64; end
		21620: begin l_1 = +27;
				 l_2 = +65; end
		24790: begin l_1 = +27;
				 l_2 = -65; end
		26071: begin l_1 = -27;
				 l_2 = +65; end
		29241: begin l_1 = -27;
				 l_2 = -65; end
		20035: begin l_1 = +27;
				 l_2 = +66; end
		26375: begin l_1 = +27;
				 l_2 = -66; end
		24486: begin l_1 = -27;
				 l_2 = +66; end
		30826: begin l_1 = -27;
				 l_2 = -66; end
		16865: begin l_1 = +27;
				 l_2 = +67; end
		29545: begin l_1 = +27;
				 l_2 = -67; end
		21316: begin l_1 = -27;
				 l_2 = +67; end
		33996: begin l_1 = -27;
				 l_2 = -67; end
		10525: begin l_1 = +27;
				 l_2 = +68; end
		35885: begin l_1 = +27;
				 l_2 = -68; end
		14976: begin l_1 = -27;
				 l_2 = +68; end
		40336: begin l_1 = -27;
				 l_2 = -68; end
		37508: begin l_1 = -28;
				 l_2 = +30; end
		13353: begin l_1 = -28;
				 l_2 = -29; end
		28606: begin l_1 = +28;
				 l_2 = +30; end
		22255: begin l_1 = -28;
				 l_2 = -30; end
		10802: begin l_1 = +28;
				 l_2 = +31; end
		31157: begin l_1 = +28;
				 l_2 = -31; end
		19704: begin l_1 = -28;
				 l_2 = +31; end
		40059: begin l_1 = -28;
				 l_2 = -31; end
		26055: begin l_1 = +28;
				 l_2 = +32; end
		15904: begin l_1 = +28;
				 l_2 = -32; end
		34957: begin l_1 = -28;
				 l_2 = +32; end
		24806: begin l_1 = -28;
				 l_2 = -32; end
		5700: begin l_1 = +28;
				 l_2 = +33; end
		36259: begin l_1 = +28;
				 l_2 = -33; end
		14602: begin l_1 = -28;
				 l_2 = +33; end
		45161: begin l_1 = -28;
				 l_2 = -33; end
		15851: begin l_1 = +28;
				 l_2 = +34; end
		26108: begin l_1 = +28;
				 l_2 = -34; end
		24753: begin l_1 = -28;
				 l_2 = +34; end
		35010: begin l_1 = -28;
				 l_2 = -34; end
		36153: begin l_1 = +28;
				 l_2 = +35; end
		5806: begin l_1 = +28;
				 l_2 = -35; end
		45055: begin l_1 = -28;
				 l_2 = +35; end
		14708: begin l_1 = -28;
				 l_2 = -35; end
		25896: begin l_1 = +28;
				 l_2 = +36; end
		16063: begin l_1 = +28;
				 l_2 = -36; end
		34798: begin l_1 = -28;
				 l_2 = +36; end
		24965: begin l_1 = -28;
				 l_2 = -36; end
		5382: begin l_1 = +28;
				 l_2 = +37; end
		36577: begin l_1 = +28;
				 l_2 = -37; end
		14284: begin l_1 = -28;
				 l_2 = +37; end
		45479: begin l_1 = -28;
				 l_2 = -37; end
		15215: begin l_1 = +28;
				 l_2 = +38; end
		26744: begin l_1 = +28;
				 l_2 = -38; end
		24117: begin l_1 = -28;
				 l_2 = +38; end
		35646: begin l_1 = -28;
				 l_2 = -38; end
		34881: begin l_1 = +28;
				 l_2 = +39; end
		7078: begin l_1 = +28;
				 l_2 = -39; end
		43783: begin l_1 = -28;
				 l_2 = +39; end
		15980: begin l_1 = -28;
				 l_2 = -39; end
		23352: begin l_1 = +28;
				 l_2 = +40; end
		18607: begin l_1 = +28;
				 l_2 = -40; end
		32254: begin l_1 = -28;
				 l_2 = +40; end
		27509: begin l_1 = -28;
				 l_2 = -40; end
		294: begin l_1 = +28;
				 l_2 = +41; end
		41665: begin l_1 = +28;
				 l_2 = -41; end
		9196: begin l_1 = -28;
				 l_2 = +41; end
		50567: begin l_1 = -28;
				 l_2 = -41; end
		5039: begin l_1 = +28;
				 l_2 = +42; end
		36920: begin l_1 = +28;
				 l_2 = -42; end
		13941: begin l_1 = -28;
				 l_2 = +42; end
		45822: begin l_1 = -28;
				 l_2 = -42; end
		14529: begin l_1 = +28;
				 l_2 = +43; end
		27430: begin l_1 = +28;
				 l_2 = -43; end
		23431: begin l_1 = -28;
				 l_2 = +43; end
		36332: begin l_1 = -28;
				 l_2 = -43; end
		33509: begin l_1 = +28;
				 l_2 = +44; end
		8450: begin l_1 = +28;
				 l_2 = -44; end
		42411: begin l_1 = -28;
				 l_2 = +44; end
		17352: begin l_1 = -28;
				 l_2 = -44; end
		20608: begin l_1 = +28;
				 l_2 = +45; end
		21351: begin l_1 = +28;
				 l_2 = -45; end
		29510: begin l_1 = -28;
				 l_2 = +45; end
		30253: begin l_1 = -28;
				 l_2 = -45; end
		45667: begin l_1 = +28;
				 l_2 = +46; end
		47153: begin l_1 = +28;
				 l_2 = -46; end
		3708: begin l_1 = -28;
				 l_2 = +46; end
		5194: begin l_1 = -28;
				 l_2 = -46; end
		44924: begin l_1 = +28;
				 l_2 = +47; end
		47896: begin l_1 = +28;
				 l_2 = -47; end
		2965: begin l_1 = -28;
				 l_2 = +47; end
		5937: begin l_1 = -28;
				 l_2 = -47; end
		43438: begin l_1 = +28;
				 l_2 = +48; end
		49382: begin l_1 = +28;
				 l_2 = -48; end
		1479: begin l_1 = -28;
				 l_2 = +48; end
		7423: begin l_1 = -28;
				 l_2 = -48; end
		40466: begin l_1 = +28;
				 l_2 = +49; end
		1493: begin l_1 = +28;
				 l_2 = -49; end
		49368: begin l_1 = -28;
				 l_2 = +49; end
		10395: begin l_1 = -28;
				 l_2 = -49; end
		34522: begin l_1 = +28;
				 l_2 = +50; end
		7437: begin l_1 = +28;
				 l_2 = -50; end
		43424: begin l_1 = -28;
				 l_2 = +50; end
		16339: begin l_1 = -28;
				 l_2 = -50; end
		22634: begin l_1 = +28;
				 l_2 = +51; end
		19325: begin l_1 = +28;
				 l_2 = -51; end
		31536: begin l_1 = -28;
				 l_2 = +51; end
		28227: begin l_1 = -28;
				 l_2 = -51; end
		49719: begin l_1 = +28;
				 l_2 = +52; end
		43101: begin l_1 = +28;
				 l_2 = -52; end
		7760: begin l_1 = -28;
				 l_2 = +52; end
		1142: begin l_1 = -28;
				 l_2 = -52; end
		2167: begin l_1 = +28;
				 l_2 = +53; end
		39792: begin l_1 = +28;
				 l_2 = -53; end
		11069: begin l_1 = -28;
				 l_2 = +53; end
		48694: begin l_1 = -28;
				 l_2 = -53; end
		8785: begin l_1 = +28;
				 l_2 = +54; end
		33174: begin l_1 = +28;
				 l_2 = -54; end
		17687: begin l_1 = -28;
				 l_2 = +54; end
		42076: begin l_1 = -28;
				 l_2 = -54; end
		22021: begin l_1 = +28;
				 l_2 = +55; end
		19938: begin l_1 = +28;
				 l_2 = -55; end
		30923: begin l_1 = -28;
				 l_2 = +55; end
		28840: begin l_1 = -28;
				 l_2 = -55; end
		48493: begin l_1 = +28;
				 l_2 = +56; end
		44327: begin l_1 = +28;
				 l_2 = -56; end
		6534: begin l_1 = -28;
				 l_2 = +56; end
		2368: begin l_1 = -28;
				 l_2 = -56; end
		50576: begin l_1 = +28;
				 l_2 = +57; end
		42244: begin l_1 = +28;
				 l_2 = -57; end
		8617: begin l_1 = -28;
				 l_2 = +57; end
		285: begin l_1 = -28;
				 l_2 = -57; end
		3881: begin l_1 = +28;
				 l_2 = +58; end
		38078: begin l_1 = +28;
				 l_2 = -58; end
		12783: begin l_1 = -28;
				 l_2 = +58; end
		46980: begin l_1 = -28;
				 l_2 = -58; end
		12213: begin l_1 = +28;
				 l_2 = +59; end
		29746: begin l_1 = +28;
				 l_2 = -59; end
		21115: begin l_1 = -28;
				 l_2 = +59; end
		38648: begin l_1 = -28;
				 l_2 = -59; end
		28877: begin l_1 = +28;
				 l_2 = +60; end
		13082: begin l_1 = +28;
				 l_2 = -60; end
		37779: begin l_1 = -28;
				 l_2 = +60; end
		21984: begin l_1 = -28;
				 l_2 = -60; end
		11344: begin l_1 = +28;
				 l_2 = +61; end
		30615: begin l_1 = +28;
				 l_2 = -61; end
		20246: begin l_1 = -28;
				 l_2 = +61; end
		39517: begin l_1 = -28;
				 l_2 = -61; end
		27139: begin l_1 = +28;
				 l_2 = +62; end
		14820: begin l_1 = +28;
				 l_2 = -62; end
		36041: begin l_1 = -28;
				 l_2 = +62; end
		23722: begin l_1 = -28;
				 l_2 = -62; end
		7868: begin l_1 = +28;
				 l_2 = +63; end
		34091: begin l_1 = +28;
				 l_2 = -63; end
		16770: begin l_1 = -28;
				 l_2 = +63; end
		42993: begin l_1 = -28;
				 l_2 = -63; end
		20187: begin l_1 = +28;
				 l_2 = +64; end
		21772: begin l_1 = +28;
				 l_2 = -64; end
		29089: begin l_1 = -28;
				 l_2 = +64; end
		30674: begin l_1 = -28;
				 l_2 = -64; end
		44825: begin l_1 = +28;
				 l_2 = +65; end
		47995: begin l_1 = +28;
				 l_2 = -65; end
		2866: begin l_1 = -28;
				 l_2 = +65; end
		6036: begin l_1 = -28;
				 l_2 = -65; end
		43240: begin l_1 = +28;
				 l_2 = +66; end
		49580: begin l_1 = +28;
				 l_2 = -66; end
		1281: begin l_1 = -28;
				 l_2 = +66; end
		7621: begin l_1 = -28;
				 l_2 = -66; end
		40070: begin l_1 = +28;
				 l_2 = +67; end
		1889: begin l_1 = +28;
				 l_2 = -67; end
		48972: begin l_1 = -28;
				 l_2 = +67; end
		10791: begin l_1 = -28;
				 l_2 = -67; end
		33730: begin l_1 = +28;
				 l_2 = +68; end
		8229: begin l_1 = +28;
				 l_2 = -68; end
		42632: begin l_1 = -28;
				 l_2 = +68; end
		17131: begin l_1 = -28;
				 l_2 = -68; end
		24155: begin l_1 = -29;
				 l_2 = +31; end
		26706: begin l_1 = -29;
				 l_2 = -30; end
		6351: begin l_1 = +29;
				 l_2 = +31; end
		44510: begin l_1 = -29;
				 l_2 = -31; end
		21604: begin l_1 = +29;
				 l_2 = +32; end
		11453: begin l_1 = +29;
				 l_2 = -32; end
		39408: begin l_1 = -29;
				 l_2 = +32; end
		29257: begin l_1 = -29;
				 l_2 = -32; end
		1249: begin l_1 = +29;
				 l_2 = +33; end
		31808: begin l_1 = +29;
				 l_2 = -33; end
		19053: begin l_1 = -29;
				 l_2 = +33; end
		49612: begin l_1 = -29;
				 l_2 = -33; end
		11400: begin l_1 = +29;
				 l_2 = +34; end
		21657: begin l_1 = +29;
				 l_2 = -34; end
		29204: begin l_1 = -29;
				 l_2 = +34; end
		39461: begin l_1 = -29;
				 l_2 = -34; end
		31702: begin l_1 = +29;
				 l_2 = +35; end
		1355: begin l_1 = +29;
				 l_2 = -35; end
		49506: begin l_1 = -29;
				 l_2 = +35; end
		19159: begin l_1 = -29;
				 l_2 = -35; end
		21445: begin l_1 = +29;
				 l_2 = +36; end
		11612: begin l_1 = +29;
				 l_2 = -36; end
		39249: begin l_1 = -29;
				 l_2 = +36; end
		29416: begin l_1 = -29;
				 l_2 = -36; end
		931: begin l_1 = +29;
				 l_2 = +37; end
		32126: begin l_1 = +29;
				 l_2 = -37; end
		18735: begin l_1 = -29;
				 l_2 = +37; end
		49930: begin l_1 = -29;
				 l_2 = -37; end
		10764: begin l_1 = +29;
				 l_2 = +38; end
		22293: begin l_1 = +29;
				 l_2 = -38; end
		28568: begin l_1 = -29;
				 l_2 = +38; end
		40097: begin l_1 = -29;
				 l_2 = -38; end
		30430: begin l_1 = +29;
				 l_2 = +39; end
		2627: begin l_1 = +29;
				 l_2 = -39; end
		48234: begin l_1 = -29;
				 l_2 = +39; end
		20431: begin l_1 = -29;
				 l_2 = -39; end
		18901: begin l_1 = +29;
				 l_2 = +40; end
		14156: begin l_1 = +29;
				 l_2 = -40; end
		36705: begin l_1 = -29;
				 l_2 = +40; end
		31960: begin l_1 = -29;
				 l_2 = -40; end
		46704: begin l_1 = +29;
				 l_2 = +41; end
		37214: begin l_1 = +29;
				 l_2 = -41; end
		13647: begin l_1 = -29;
				 l_2 = +41; end
		4157: begin l_1 = -29;
				 l_2 = -41; end
		588: begin l_1 = +29;
				 l_2 = +42; end
		32469: begin l_1 = +29;
				 l_2 = -42; end
		18392: begin l_1 = -29;
				 l_2 = +42; end
		50273: begin l_1 = -29;
				 l_2 = -42; end
		10078: begin l_1 = +29;
				 l_2 = +43; end
		22979: begin l_1 = +29;
				 l_2 = -43; end
		27882: begin l_1 = -29;
				 l_2 = +43; end
		40783: begin l_1 = -29;
				 l_2 = -43; end
		29058: begin l_1 = +29;
				 l_2 = +44; end
		3999: begin l_1 = +29;
				 l_2 = -44; end
		46862: begin l_1 = -29;
				 l_2 = +44; end
		21803: begin l_1 = -29;
				 l_2 = -44; end
		16157: begin l_1 = +29;
				 l_2 = +45; end
		16900: begin l_1 = +29;
				 l_2 = -45; end
		33961: begin l_1 = -29;
				 l_2 = +45; end
		34704: begin l_1 = -29;
				 l_2 = -45; end
		41216: begin l_1 = +29;
				 l_2 = +46; end
		42702: begin l_1 = +29;
				 l_2 = -46; end
		8159: begin l_1 = -29;
				 l_2 = +46; end
		9645: begin l_1 = -29;
				 l_2 = -46; end
		40473: begin l_1 = +29;
				 l_2 = +47; end
		43445: begin l_1 = +29;
				 l_2 = -47; end
		7416: begin l_1 = -29;
				 l_2 = +47; end
		10388: begin l_1 = -29;
				 l_2 = -47; end
		38987: begin l_1 = +29;
				 l_2 = +48; end
		44931: begin l_1 = +29;
				 l_2 = -48; end
		5930: begin l_1 = -29;
				 l_2 = +48; end
		11874: begin l_1 = -29;
				 l_2 = -48; end
		36015: begin l_1 = +29;
				 l_2 = +49; end
		47903: begin l_1 = +29;
				 l_2 = -49; end
		2958: begin l_1 = -29;
				 l_2 = +49; end
		14846: begin l_1 = -29;
				 l_2 = -49; end
		30071: begin l_1 = +29;
				 l_2 = +50; end
		2986: begin l_1 = +29;
				 l_2 = -50; end
		47875: begin l_1 = -29;
				 l_2 = +50; end
		20790: begin l_1 = -29;
				 l_2 = -50; end
		18183: begin l_1 = +29;
				 l_2 = +51; end
		14874: begin l_1 = +29;
				 l_2 = -51; end
		35987: begin l_1 = -29;
				 l_2 = +51; end
		32678: begin l_1 = -29;
				 l_2 = -51; end
		45268: begin l_1 = +29;
				 l_2 = +52; end
		38650: begin l_1 = +29;
				 l_2 = -52; end
		12211: begin l_1 = -29;
				 l_2 = +52; end
		5593: begin l_1 = -29;
				 l_2 = -52; end
		48577: begin l_1 = +29;
				 l_2 = +53; end
		35341: begin l_1 = +29;
				 l_2 = -53; end
		15520: begin l_1 = -29;
				 l_2 = +53; end
		2284: begin l_1 = -29;
				 l_2 = -53; end
		4334: begin l_1 = +29;
				 l_2 = +54; end
		28723: begin l_1 = +29;
				 l_2 = -54; end
		22138: begin l_1 = -29;
				 l_2 = +54; end
		46527: begin l_1 = -29;
				 l_2 = -54; end
		17570: begin l_1 = +29;
				 l_2 = +55; end
		15487: begin l_1 = +29;
				 l_2 = -55; end
		35374: begin l_1 = -29;
				 l_2 = +55; end
		33291: begin l_1 = -29;
				 l_2 = -55; end
		44042: begin l_1 = +29;
				 l_2 = +56; end
		39876: begin l_1 = +29;
				 l_2 = -56; end
		10985: begin l_1 = -29;
				 l_2 = +56; end
		6819: begin l_1 = -29;
				 l_2 = -56; end
		46125: begin l_1 = +29;
				 l_2 = +57; end
		37793: begin l_1 = +29;
				 l_2 = -57; end
		13068: begin l_1 = -29;
				 l_2 = +57; end
		4736: begin l_1 = -29;
				 l_2 = -57; end
		50291: begin l_1 = +29;
				 l_2 = +58; end
		33627: begin l_1 = +29;
				 l_2 = -58; end
		17234: begin l_1 = -29;
				 l_2 = +58; end
		570: begin l_1 = -29;
				 l_2 = -58; end
		7762: begin l_1 = +29;
				 l_2 = +59; end
		25295: begin l_1 = +29;
				 l_2 = -59; end
		25566: begin l_1 = -29;
				 l_2 = +59; end
		43099: begin l_1 = -29;
				 l_2 = -59; end
		24426: begin l_1 = +29;
				 l_2 = +60; end
		8631: begin l_1 = +29;
				 l_2 = -60; end
		42230: begin l_1 = -29;
				 l_2 = +60; end
		26435: begin l_1 = -29;
				 l_2 = -60; end
		6893: begin l_1 = +29;
				 l_2 = +61; end
		26164: begin l_1 = +29;
				 l_2 = -61; end
		24697: begin l_1 = -29;
				 l_2 = +61; end
		43968: begin l_1 = -29;
				 l_2 = -61; end
		22688: begin l_1 = +29;
				 l_2 = +62; end
		10369: begin l_1 = +29;
				 l_2 = -62; end
		40492: begin l_1 = -29;
				 l_2 = +62; end
		28173: begin l_1 = -29;
				 l_2 = -62; end
		3417: begin l_1 = +29;
				 l_2 = +63; end
		29640: begin l_1 = +29;
				 l_2 = -63; end
		21221: begin l_1 = -29;
				 l_2 = +63; end
		47444: begin l_1 = -29;
				 l_2 = -63; end
		15736: begin l_1 = +29;
				 l_2 = +64; end
		17321: begin l_1 = +29;
				 l_2 = -64; end
		33540: begin l_1 = -29;
				 l_2 = +64; end
		35125: begin l_1 = -29;
				 l_2 = -64; end
		40374: begin l_1 = +29;
				 l_2 = +65; end
		43544: begin l_1 = +29;
				 l_2 = -65; end
		7317: begin l_1 = -29;
				 l_2 = +65; end
		10487: begin l_1 = -29;
				 l_2 = -65; end
		38789: begin l_1 = +29;
				 l_2 = +66; end
		45129: begin l_1 = +29;
				 l_2 = -66; end
		5732: begin l_1 = -29;
				 l_2 = +66; end
		12072: begin l_1 = -29;
				 l_2 = -66; end
		35619: begin l_1 = +29;
				 l_2 = +67; end
		48299: begin l_1 = +29;
				 l_2 = -67; end
		2562: begin l_1 = -29;
				 l_2 = +67; end
		15242: begin l_1 = -29;
				 l_2 = -67; end
		29279: begin l_1 = +29;
				 l_2 = +68; end
		3778: begin l_1 = +29;
				 l_2 = -68; end
		47083: begin l_1 = -29;
				 l_2 = +68; end
		21582: begin l_1 = -29;
				 l_2 = -68; end
		48310: begin l_1 = -30;
				 l_2 = +32; end
		2551: begin l_1 = -30;
				 l_2 = -31; end
		12702: begin l_1 = +30;
				 l_2 = +32; end
		38159: begin l_1 = -30;
				 l_2 = -32; end
		43208: begin l_1 = +30;
				 l_2 = +33; end
		22906: begin l_1 = +30;
				 l_2 = -33; end
		27955: begin l_1 = -30;
				 l_2 = +33; end
		7653: begin l_1 = -30;
				 l_2 = -33; end
		2498: begin l_1 = +30;
				 l_2 = +34; end
		12755: begin l_1 = +30;
				 l_2 = -34; end
		38106: begin l_1 = -30;
				 l_2 = +34; end
		48363: begin l_1 = -30;
				 l_2 = -34; end
		22800: begin l_1 = +30;
				 l_2 = +35; end
		43314: begin l_1 = +30;
				 l_2 = -35; end
		7547: begin l_1 = -30;
				 l_2 = +35; end
		28061: begin l_1 = -30;
				 l_2 = -35; end
		12543: begin l_1 = +30;
				 l_2 = +36; end
		2710: begin l_1 = +30;
				 l_2 = -36; end
		48151: begin l_1 = -30;
				 l_2 = +36; end
		38318: begin l_1 = -30;
				 l_2 = -36; end
		42890: begin l_1 = +30;
				 l_2 = +37; end
		23224: begin l_1 = +30;
				 l_2 = -37; end
		27637: begin l_1 = -30;
				 l_2 = +37; end
		7971: begin l_1 = -30;
				 l_2 = -37; end
		1862: begin l_1 = +30;
				 l_2 = +38; end
		13391: begin l_1 = +30;
				 l_2 = -38; end
		37470: begin l_1 = -30;
				 l_2 = +38; end
		48999: begin l_1 = -30;
				 l_2 = -38; end
		21528: begin l_1 = +30;
				 l_2 = +39; end
		44586: begin l_1 = +30;
				 l_2 = -39; end
		6275: begin l_1 = -30;
				 l_2 = +39; end
		29333: begin l_1 = -30;
				 l_2 = -39; end
		9999: begin l_1 = +30;
				 l_2 = +40; end
		5254: begin l_1 = +30;
				 l_2 = -40; end
		45607: begin l_1 = -30;
				 l_2 = +40; end
		40862: begin l_1 = -30;
				 l_2 = -40; end
		37802: begin l_1 = +30;
				 l_2 = +41; end
		28312: begin l_1 = +30;
				 l_2 = -41; end
		22549: begin l_1 = -30;
				 l_2 = +41; end
		13059: begin l_1 = -30;
				 l_2 = -41; end
		42547: begin l_1 = +30;
				 l_2 = +42; end
		23567: begin l_1 = +30;
				 l_2 = -42; end
		27294: begin l_1 = -30;
				 l_2 = +42; end
		8314: begin l_1 = -30;
				 l_2 = -42; end
		1176: begin l_1 = +30;
				 l_2 = +43; end
		14077: begin l_1 = +30;
				 l_2 = -43; end
		36784: begin l_1 = -30;
				 l_2 = +43; end
		49685: begin l_1 = -30;
				 l_2 = -43; end
		20156: begin l_1 = +30;
				 l_2 = +44; end
		45958: begin l_1 = +30;
				 l_2 = -44; end
		4903: begin l_1 = -30;
				 l_2 = +44; end
		30705: begin l_1 = -30;
				 l_2 = -44; end
		7255: begin l_1 = +30;
				 l_2 = +45; end
		7998: begin l_1 = +30;
				 l_2 = -45; end
		42863: begin l_1 = -30;
				 l_2 = +45; end
		43606: begin l_1 = -30;
				 l_2 = -45; end
		32314: begin l_1 = +30;
				 l_2 = +46; end
		33800: begin l_1 = +30;
				 l_2 = -46; end
		17061: begin l_1 = -30;
				 l_2 = +46; end
		18547: begin l_1 = -30;
				 l_2 = -46; end
		31571: begin l_1 = +30;
				 l_2 = +47; end
		34543: begin l_1 = +30;
				 l_2 = -47; end
		16318: begin l_1 = -30;
				 l_2 = +47; end
		19290: begin l_1 = -30;
				 l_2 = -47; end
		30085: begin l_1 = +30;
				 l_2 = +48; end
		36029: begin l_1 = +30;
				 l_2 = -48; end
		14832: begin l_1 = -30;
				 l_2 = +48; end
		20776: begin l_1 = -30;
				 l_2 = -48; end
		27113: begin l_1 = +30;
				 l_2 = +49; end
		39001: begin l_1 = +30;
				 l_2 = -49; end
		11860: begin l_1 = -30;
				 l_2 = +49; end
		23748: begin l_1 = -30;
				 l_2 = -49; end
		21169: begin l_1 = +30;
				 l_2 = +50; end
		44945: begin l_1 = +30;
				 l_2 = -50; end
		5916: begin l_1 = -30;
				 l_2 = +50; end
		29692: begin l_1 = -30;
				 l_2 = -50; end
		9281: begin l_1 = +30;
				 l_2 = +51; end
		5972: begin l_1 = +30;
				 l_2 = -51; end
		44889: begin l_1 = -30;
				 l_2 = +51; end
		41580: begin l_1 = -30;
				 l_2 = -51; end
		36366: begin l_1 = +30;
				 l_2 = +52; end
		29748: begin l_1 = +30;
				 l_2 = -52; end
		21113: begin l_1 = -30;
				 l_2 = +52; end
		14495: begin l_1 = -30;
				 l_2 = -52; end
		39675: begin l_1 = +30;
				 l_2 = +53; end
		26439: begin l_1 = +30;
				 l_2 = -53; end
		24422: begin l_1 = -30;
				 l_2 = +53; end
		11186: begin l_1 = -30;
				 l_2 = -53; end
		46293: begin l_1 = +30;
				 l_2 = +54; end
		19821: begin l_1 = +30;
				 l_2 = -54; end
		31040: begin l_1 = -30;
				 l_2 = +54; end
		4568: begin l_1 = -30;
				 l_2 = -54; end
		8668: begin l_1 = +30;
				 l_2 = +55; end
		6585: begin l_1 = +30;
				 l_2 = -55; end
		44276: begin l_1 = -30;
				 l_2 = +55; end
		42193: begin l_1 = -30;
				 l_2 = -55; end
		35140: begin l_1 = +30;
				 l_2 = +56; end
		30974: begin l_1 = +30;
				 l_2 = -56; end
		19887: begin l_1 = -30;
				 l_2 = +56; end
		15721: begin l_1 = -30;
				 l_2 = -56; end
		37223: begin l_1 = +30;
				 l_2 = +57; end
		28891: begin l_1 = +30;
				 l_2 = -57; end
		21970: begin l_1 = -30;
				 l_2 = +57; end
		13638: begin l_1 = -30;
				 l_2 = -57; end
		41389: begin l_1 = +30;
				 l_2 = +58; end
		24725: begin l_1 = +30;
				 l_2 = -58; end
		26136: begin l_1 = -30;
				 l_2 = +58; end
		9472: begin l_1 = -30;
				 l_2 = -58; end
		49721: begin l_1 = +30;
				 l_2 = +59; end
		16393: begin l_1 = +30;
				 l_2 = -59; end
		34468: begin l_1 = -30;
				 l_2 = +59; end
		1140: begin l_1 = -30;
				 l_2 = -59; end
		15524: begin l_1 = +30;
				 l_2 = +60; end
		50590: begin l_1 = +30;
				 l_2 = -60; end
		271: begin l_1 = -30;
				 l_2 = +60; end
		35337: begin l_1 = -30;
				 l_2 = -60; end
		48852: begin l_1 = +30;
				 l_2 = +61; end
		17262: begin l_1 = +30;
				 l_2 = -61; end
		33599: begin l_1 = -30;
				 l_2 = +61; end
		2009: begin l_1 = -30;
				 l_2 = -61; end
		13786: begin l_1 = +30;
				 l_2 = +62; end
		1467: begin l_1 = +30;
				 l_2 = -62; end
		49394: begin l_1 = -30;
				 l_2 = +62; end
		37075: begin l_1 = -30;
				 l_2 = -62; end
		45376: begin l_1 = +30;
				 l_2 = +63; end
		20738: begin l_1 = +30;
				 l_2 = -63; end
		30123: begin l_1 = -30;
				 l_2 = +63; end
		5485: begin l_1 = -30;
				 l_2 = -63; end
		6834: begin l_1 = +30;
				 l_2 = +64; end
		8419: begin l_1 = +30;
				 l_2 = -64; end
		42442: begin l_1 = -30;
				 l_2 = +64; end
		44027: begin l_1 = -30;
				 l_2 = -64; end
		31472: begin l_1 = +30;
				 l_2 = +65; end
		34642: begin l_1 = +30;
				 l_2 = -65; end
		16219: begin l_1 = -30;
				 l_2 = +65; end
		19389: begin l_1 = -30;
				 l_2 = -65; end
		29887: begin l_1 = +30;
				 l_2 = +66; end
		36227: begin l_1 = +30;
				 l_2 = -66; end
		14634: begin l_1 = -30;
				 l_2 = +66; end
		20974: begin l_1 = -30;
				 l_2 = -66; end
		26717: begin l_1 = +30;
				 l_2 = +67; end
		39397: begin l_1 = +30;
				 l_2 = -67; end
		11464: begin l_1 = -30;
				 l_2 = +67; end
		24144: begin l_1 = -30;
				 l_2 = -67; end
		20377: begin l_1 = +30;
				 l_2 = +68; end
		45737: begin l_1 = +30;
				 l_2 = -68; end
		5124: begin l_1 = -30;
				 l_2 = +68; end
		30484: begin l_1 = -30;
				 l_2 = -68; end
		45759: begin l_1 = -31;
				 l_2 = +33; end
		5102: begin l_1 = -31;
				 l_2 = -32; end
		25404: begin l_1 = +31;
				 l_2 = +33; end
		25457: begin l_1 = -31;
				 l_2 = -33; end
		35555: begin l_1 = +31;
				 l_2 = +34; end
		45812: begin l_1 = +31;
				 l_2 = -34; end
		5049: begin l_1 = -31;
				 l_2 = +34; end
		15306: begin l_1 = -31;
				 l_2 = -34; end
		4996: begin l_1 = +31;
				 l_2 = +35; end
		25510: begin l_1 = +31;
				 l_2 = -35; end
		25351: begin l_1 = -31;
				 l_2 = +35; end
		45865: begin l_1 = -31;
				 l_2 = -35; end
		45600: begin l_1 = +31;
				 l_2 = +36; end
		35767: begin l_1 = +31;
				 l_2 = -36; end
		15094: begin l_1 = -31;
				 l_2 = +36; end
		5261: begin l_1 = -31;
				 l_2 = -36; end
		25086: begin l_1 = +31;
				 l_2 = +37; end
		5420: begin l_1 = +31;
				 l_2 = -37; end
		45441: begin l_1 = -31;
				 l_2 = +37; end
		25775: begin l_1 = -31;
				 l_2 = -37; end
		34919: begin l_1 = +31;
				 l_2 = +38; end
		46448: begin l_1 = +31;
				 l_2 = -38; end
		4413: begin l_1 = -31;
				 l_2 = +38; end
		15942: begin l_1 = -31;
				 l_2 = -38; end
		3724: begin l_1 = +31;
				 l_2 = +39; end
		26782: begin l_1 = +31;
				 l_2 = -39; end
		24079: begin l_1 = -31;
				 l_2 = +39; end
		47137: begin l_1 = -31;
				 l_2 = -39; end
		43056: begin l_1 = +31;
				 l_2 = +40; end
		38311: begin l_1 = +31;
				 l_2 = -40; end
		12550: begin l_1 = -31;
				 l_2 = +40; end
		7805: begin l_1 = -31;
				 l_2 = -40; end
		19998: begin l_1 = +31;
				 l_2 = +41; end
		10508: begin l_1 = +31;
				 l_2 = -41; end
		40353: begin l_1 = -31;
				 l_2 = +41; end
		30863: begin l_1 = -31;
				 l_2 = -41; end
		24743: begin l_1 = +31;
				 l_2 = +42; end
		5763: begin l_1 = +31;
				 l_2 = -42; end
		45098: begin l_1 = -31;
				 l_2 = +42; end
		26118: begin l_1 = -31;
				 l_2 = -42; end
		34233: begin l_1 = +31;
				 l_2 = +43; end
		47134: begin l_1 = +31;
				 l_2 = -43; end
		3727: begin l_1 = -31;
				 l_2 = +43; end
		16628: begin l_1 = -31;
				 l_2 = -43; end
		2352: begin l_1 = +31;
				 l_2 = +44; end
		28154: begin l_1 = +31;
				 l_2 = -44; end
		22707: begin l_1 = -31;
				 l_2 = +44; end
		48509: begin l_1 = -31;
				 l_2 = -44; end
		40312: begin l_1 = +31;
				 l_2 = +45; end
		41055: begin l_1 = +31;
				 l_2 = -45; end
		9806: begin l_1 = -31;
				 l_2 = +45; end
		10549: begin l_1 = -31;
				 l_2 = -45; end
		14510: begin l_1 = +31;
				 l_2 = +46; end
		15996: begin l_1 = +31;
				 l_2 = -46; end
		34865: begin l_1 = -31;
				 l_2 = +46; end
		36351: begin l_1 = -31;
				 l_2 = -46; end
		13767: begin l_1 = +31;
				 l_2 = +47; end
		16739: begin l_1 = +31;
				 l_2 = -47; end
		34122: begin l_1 = -31;
				 l_2 = +47; end
		37094: begin l_1 = -31;
				 l_2 = -47; end
		12281: begin l_1 = +31;
				 l_2 = +48; end
		18225: begin l_1 = +31;
				 l_2 = -48; end
		32636: begin l_1 = -31;
				 l_2 = +48; end
		38580: begin l_1 = -31;
				 l_2 = -48; end
		9309: begin l_1 = +31;
				 l_2 = +49; end
		21197: begin l_1 = +31;
				 l_2 = -49; end
		29664: begin l_1 = -31;
				 l_2 = +49; end
		41552: begin l_1 = -31;
				 l_2 = -49; end
		3365: begin l_1 = +31;
				 l_2 = +50; end
		27141: begin l_1 = +31;
				 l_2 = -50; end
		23720: begin l_1 = -31;
				 l_2 = +50; end
		47496: begin l_1 = -31;
				 l_2 = -50; end
		42338: begin l_1 = +31;
				 l_2 = +51; end
		39029: begin l_1 = +31;
				 l_2 = -51; end
		11832: begin l_1 = -31;
				 l_2 = +51; end
		8523: begin l_1 = -31;
				 l_2 = -51; end
		18562: begin l_1 = +31;
				 l_2 = +52; end
		11944: begin l_1 = +31;
				 l_2 = -52; end
		38917: begin l_1 = -31;
				 l_2 = +52; end
		32299: begin l_1 = -31;
				 l_2 = -52; end
		21871: begin l_1 = +31;
				 l_2 = +53; end
		8635: begin l_1 = +31;
				 l_2 = -53; end
		42226: begin l_1 = -31;
				 l_2 = +53; end
		28990: begin l_1 = -31;
				 l_2 = -53; end
		28489: begin l_1 = +31;
				 l_2 = +54; end
		2017: begin l_1 = +31;
				 l_2 = -54; end
		48844: begin l_1 = -31;
				 l_2 = +54; end
		22372: begin l_1 = -31;
				 l_2 = -54; end
		41725: begin l_1 = +31;
				 l_2 = +55; end
		39642: begin l_1 = +31;
				 l_2 = -55; end
		11219: begin l_1 = -31;
				 l_2 = +55; end
		9136: begin l_1 = -31;
				 l_2 = -55; end
		17336: begin l_1 = +31;
				 l_2 = +56; end
		13170: begin l_1 = +31;
				 l_2 = -56; end
		37691: begin l_1 = -31;
				 l_2 = +56; end
		33525: begin l_1 = -31;
				 l_2 = -56; end
		19419: begin l_1 = +31;
				 l_2 = +57; end
		11087: begin l_1 = +31;
				 l_2 = -57; end
		39774: begin l_1 = -31;
				 l_2 = +57; end
		31442: begin l_1 = -31;
				 l_2 = -57; end
		23585: begin l_1 = +31;
				 l_2 = +58; end
		6921: begin l_1 = +31;
				 l_2 = -58; end
		43940: begin l_1 = -31;
				 l_2 = +58; end
		27276: begin l_1 = -31;
				 l_2 = -58; end
		31917: begin l_1 = +31;
				 l_2 = +59; end
		49450: begin l_1 = +31;
				 l_2 = -59; end
		1411: begin l_1 = -31;
				 l_2 = +59; end
		18944: begin l_1 = -31;
				 l_2 = -59; end
		48581: begin l_1 = +31;
				 l_2 = +60; end
		32786: begin l_1 = +31;
				 l_2 = -60; end
		18075: begin l_1 = -31;
				 l_2 = +60; end
		2280: begin l_1 = -31;
				 l_2 = -60; end
		31048: begin l_1 = +31;
				 l_2 = +61; end
		50319: begin l_1 = +31;
				 l_2 = -61; end
		542: begin l_1 = -31;
				 l_2 = +61; end
		19813: begin l_1 = -31;
				 l_2 = -61; end
		46843: begin l_1 = +31;
				 l_2 = +62; end
		34524: begin l_1 = +31;
				 l_2 = -62; end
		16337: begin l_1 = -31;
				 l_2 = +62; end
		4018: begin l_1 = -31;
				 l_2 = -62; end
		27572: begin l_1 = +31;
				 l_2 = +63; end
		2934: begin l_1 = +31;
				 l_2 = -63; end
		47927: begin l_1 = -31;
				 l_2 = +63; end
		23289: begin l_1 = -31;
				 l_2 = -63; end
		39891: begin l_1 = +31;
				 l_2 = +64; end
		41476: begin l_1 = +31;
				 l_2 = -64; end
		9385: begin l_1 = -31;
				 l_2 = +64; end
		10970: begin l_1 = -31;
				 l_2 = -64; end
		13668: begin l_1 = +31;
				 l_2 = +65; end
		16838: begin l_1 = +31;
				 l_2 = -65; end
		34023: begin l_1 = -31;
				 l_2 = +65; end
		37193: begin l_1 = -31;
				 l_2 = -65; end
		12083: begin l_1 = +31;
				 l_2 = +66; end
		18423: begin l_1 = +31;
				 l_2 = -66; end
		32438: begin l_1 = -31;
				 l_2 = +66; end
		38778: begin l_1 = -31;
				 l_2 = -66; end
		8913: begin l_1 = +31;
				 l_2 = +67; end
		21593: begin l_1 = +31;
				 l_2 = -67; end
		29268: begin l_1 = -31;
				 l_2 = +67; end
		41948: begin l_1 = -31;
				 l_2 = -67; end
		2573: begin l_1 = +31;
				 l_2 = +68; end
		27933: begin l_1 = +31;
				 l_2 = -68; end
		22928: begin l_1 = -31;
				 l_2 = +68; end
		48288: begin l_1 = -31;
				 l_2 = -68; end
		40657: begin l_1 = -32;
				 l_2 = +34; end
		10204: begin l_1 = -32;
				 l_2 = -33; end
		50808: begin l_1 = +32;
				 l_2 = +34; end
		53: begin l_1 = -32;
				 l_2 = -34; end
		20249: begin l_1 = +32;
				 l_2 = +35; end
		40763: begin l_1 = +32;
				 l_2 = -35; end
		10098: begin l_1 = -32;
				 l_2 = +35; end
		30612: begin l_1 = -32;
				 l_2 = -35; end
		9992: begin l_1 = +32;
				 l_2 = +36; end
		159: begin l_1 = +32;
				 l_2 = -36; end
		50702: begin l_1 = -32;
				 l_2 = +36; end
		40869: begin l_1 = -32;
				 l_2 = -36; end
		40339: begin l_1 = +32;
				 l_2 = +37; end
		20673: begin l_1 = +32;
				 l_2 = -37; end
		30188: begin l_1 = -32;
				 l_2 = +37; end
		10522: begin l_1 = -32;
				 l_2 = -37; end
		50172: begin l_1 = +32;
				 l_2 = +38; end
		10840: begin l_1 = +32;
				 l_2 = -38; end
		40021: begin l_1 = -32;
				 l_2 = +38; end
		689: begin l_1 = -32;
				 l_2 = -38; end
		18977: begin l_1 = +32;
				 l_2 = +39; end
		42035: begin l_1 = +32;
				 l_2 = -39; end
		8826: begin l_1 = -32;
				 l_2 = +39; end
		31884: begin l_1 = -32;
				 l_2 = -39; end
		7448: begin l_1 = +32;
				 l_2 = +40; end
		2703: begin l_1 = +32;
				 l_2 = -40; end
		48158: begin l_1 = -32;
				 l_2 = +40; end
		43413: begin l_1 = -32;
				 l_2 = -40; end
		35251: begin l_1 = +32;
				 l_2 = +41; end
		25761: begin l_1 = +32;
				 l_2 = -41; end
		25100: begin l_1 = -32;
				 l_2 = +41; end
		15610: begin l_1 = -32;
				 l_2 = -41; end
		39996: begin l_1 = +32;
				 l_2 = +42; end
		21016: begin l_1 = +32;
				 l_2 = -42; end
		29845: begin l_1 = -32;
				 l_2 = +42; end
		10865: begin l_1 = -32;
				 l_2 = -42; end
		49486: begin l_1 = +32;
				 l_2 = +43; end
		11526: begin l_1 = +32;
				 l_2 = -43; end
		39335: begin l_1 = -32;
				 l_2 = +43; end
		1375: begin l_1 = -32;
				 l_2 = -43; end
		17605: begin l_1 = +32;
				 l_2 = +44; end
		43407: begin l_1 = +32;
				 l_2 = -44; end
		7454: begin l_1 = -32;
				 l_2 = +44; end
		33256: begin l_1 = -32;
				 l_2 = -44; end
		4704: begin l_1 = +32;
				 l_2 = +45; end
		5447: begin l_1 = +32;
				 l_2 = -45; end
		45414: begin l_1 = -32;
				 l_2 = +45; end
		46157: begin l_1 = -32;
				 l_2 = -45; end
		29763: begin l_1 = +32;
				 l_2 = +46; end
		31249: begin l_1 = +32;
				 l_2 = -46; end
		19612: begin l_1 = -32;
				 l_2 = +46; end
		21098: begin l_1 = -32;
				 l_2 = -46; end
		29020: begin l_1 = +32;
				 l_2 = +47; end
		31992: begin l_1 = +32;
				 l_2 = -47; end
		18869: begin l_1 = -32;
				 l_2 = +47; end
		21841: begin l_1 = -32;
				 l_2 = -47; end
		27534: begin l_1 = +32;
				 l_2 = +48; end
		33478: begin l_1 = +32;
				 l_2 = -48; end
		17383: begin l_1 = -32;
				 l_2 = +48; end
		23327: begin l_1 = -32;
				 l_2 = -48; end
		24562: begin l_1 = +32;
				 l_2 = +49; end
		36450: begin l_1 = +32;
				 l_2 = -49; end
		14411: begin l_1 = -32;
				 l_2 = +49; end
		26299: begin l_1 = -32;
				 l_2 = -49; end
		18618: begin l_1 = +32;
				 l_2 = +50; end
		42394: begin l_1 = +32;
				 l_2 = -50; end
		8467: begin l_1 = -32;
				 l_2 = +50; end
		32243: begin l_1 = -32;
				 l_2 = -50; end
		6730: begin l_1 = +32;
				 l_2 = +51; end
		3421: begin l_1 = +32;
				 l_2 = -51; end
		47440: begin l_1 = -32;
				 l_2 = +51; end
		44131: begin l_1 = -32;
				 l_2 = -51; end
		33815: begin l_1 = +32;
				 l_2 = +52; end
		27197: begin l_1 = +32;
				 l_2 = -52; end
		23664: begin l_1 = -32;
				 l_2 = +52; end
		17046: begin l_1 = -32;
				 l_2 = -52; end
		37124: begin l_1 = +32;
				 l_2 = +53; end
		23888: begin l_1 = +32;
				 l_2 = -53; end
		26973: begin l_1 = -32;
				 l_2 = +53; end
		13737: begin l_1 = -32;
				 l_2 = -53; end
		43742: begin l_1 = +32;
				 l_2 = +54; end
		17270: begin l_1 = +32;
				 l_2 = -54; end
		33591: begin l_1 = -32;
				 l_2 = +54; end
		7119: begin l_1 = -32;
				 l_2 = -54; end
		6117: begin l_1 = +32;
				 l_2 = +55; end
		4034: begin l_1 = +32;
				 l_2 = -55; end
		46827: begin l_1 = -32;
				 l_2 = +55; end
		44744: begin l_1 = -32;
				 l_2 = -55; end
		32589: begin l_1 = +32;
				 l_2 = +56; end
		28423: begin l_1 = +32;
				 l_2 = -56; end
		22438: begin l_1 = -32;
				 l_2 = +56; end
		18272: begin l_1 = -32;
				 l_2 = -56; end
		34672: begin l_1 = +32;
				 l_2 = +57; end
		26340: begin l_1 = +32;
				 l_2 = -57; end
		24521: begin l_1 = -32;
				 l_2 = +57; end
		16189: begin l_1 = -32;
				 l_2 = -57; end
		38838: begin l_1 = +32;
				 l_2 = +58; end
		22174: begin l_1 = +32;
				 l_2 = -58; end
		28687: begin l_1 = -32;
				 l_2 = +58; end
		12023: begin l_1 = -32;
				 l_2 = -58; end
		47170: begin l_1 = +32;
				 l_2 = +59; end
		13842: begin l_1 = +32;
				 l_2 = -59; end
		37019: begin l_1 = -32;
				 l_2 = +59; end
		3691: begin l_1 = -32;
				 l_2 = -59; end
		12973: begin l_1 = +32;
				 l_2 = +60; end
		48039: begin l_1 = +32;
				 l_2 = -60; end
		2822: begin l_1 = -32;
				 l_2 = +60; end
		37888: begin l_1 = -32;
				 l_2 = -60; end
		46301: begin l_1 = +32;
				 l_2 = +61; end
		14711: begin l_1 = +32;
				 l_2 = -61; end
		36150: begin l_1 = -32;
				 l_2 = +61; end
		4560: begin l_1 = -32;
				 l_2 = -61; end
		11235: begin l_1 = +32;
				 l_2 = +62; end
		49777: begin l_1 = +32;
				 l_2 = -62; end
		1084: begin l_1 = -32;
				 l_2 = +62; end
		39626: begin l_1 = -32;
				 l_2 = -62; end
		42825: begin l_1 = +32;
				 l_2 = +63; end
		18187: begin l_1 = +32;
				 l_2 = -63; end
		32674: begin l_1 = -32;
				 l_2 = +63; end
		8036: begin l_1 = -32;
				 l_2 = -63; end
		4283: begin l_1 = +32;
				 l_2 = +64; end
		5868: begin l_1 = +32;
				 l_2 = -64; end
		44993: begin l_1 = -32;
				 l_2 = +64; end
		46578: begin l_1 = -32;
				 l_2 = -64; end
		28921: begin l_1 = +32;
				 l_2 = +65; end
		32091: begin l_1 = +32;
				 l_2 = -65; end
		18770: begin l_1 = -32;
				 l_2 = +65; end
		21940: begin l_1 = -32;
				 l_2 = -65; end
		27336: begin l_1 = +32;
				 l_2 = +66; end
		33676: begin l_1 = +32;
				 l_2 = -66; end
		17185: begin l_1 = -32;
				 l_2 = +66; end
		23525: begin l_1 = -32;
				 l_2 = -66; end
		24166: begin l_1 = +32;
				 l_2 = +67; end
		36846: begin l_1 = +32;
				 l_2 = -67; end
		14015: begin l_1 = -32;
				 l_2 = +67; end
		26695: begin l_1 = -32;
				 l_2 = -67; end
		17826: begin l_1 = +32;
				 l_2 = +68; end
		43186: begin l_1 = +32;
				 l_2 = -68; end
		7675: begin l_1 = -32;
				 l_2 = +68; end
		33035: begin l_1 = -32;
				 l_2 = -68; end
		30453: begin l_1 = -33;
				 l_2 = +35; end
		20408: begin l_1 = -33;
				 l_2 = -34; end
		50755: begin l_1 = +33;
				 l_2 = +35; end
		106: begin l_1 = -33;
				 l_2 = -35; end
		40498: begin l_1 = +33;
				 l_2 = +36; end
		30665: begin l_1 = +33;
				 l_2 = -36; end
		20196: begin l_1 = -33;
				 l_2 = +36; end
		10363: begin l_1 = -33;
				 l_2 = -36; end
		19984: begin l_1 = +33;
				 l_2 = +37; end
		318: begin l_1 = +33;
				 l_2 = -37; end
		50543: begin l_1 = -33;
				 l_2 = +37; end
		30877: begin l_1 = -33;
				 l_2 = -37; end
		29817: begin l_1 = +33;
				 l_2 = +38; end
		41346: begin l_1 = +33;
				 l_2 = -38; end
		9515: begin l_1 = -33;
				 l_2 = +38; end
		21044: begin l_1 = -33;
				 l_2 = -38; end
		49483: begin l_1 = +33;
				 l_2 = +39; end
		21680: begin l_1 = +33;
				 l_2 = -39; end
		29181: begin l_1 = -33;
				 l_2 = +39; end
		1378: begin l_1 = -33;
				 l_2 = -39; end
		37954: begin l_1 = +33;
				 l_2 = +40; end
		33209: begin l_1 = +33;
				 l_2 = -40; end
		17652: begin l_1 = -33;
				 l_2 = +40; end
		12907: begin l_1 = -33;
				 l_2 = -40; end
		14896: begin l_1 = +33;
				 l_2 = +41; end
		5406: begin l_1 = +33;
				 l_2 = -41; end
		45455: begin l_1 = -33;
				 l_2 = +41; end
		35965: begin l_1 = -33;
				 l_2 = -41; end
		19641: begin l_1 = +33;
				 l_2 = +42; end
		661: begin l_1 = +33;
				 l_2 = -42; end
		50200: begin l_1 = -33;
				 l_2 = +42; end
		31220: begin l_1 = -33;
				 l_2 = -42; end
		29131: begin l_1 = +33;
				 l_2 = +43; end
		42032: begin l_1 = +33;
				 l_2 = -43; end
		8829: begin l_1 = -33;
				 l_2 = +43; end
		21730: begin l_1 = -33;
				 l_2 = -43; end
		48111: begin l_1 = +33;
				 l_2 = +44; end
		23052: begin l_1 = +33;
				 l_2 = -44; end
		27809: begin l_1 = -33;
				 l_2 = +44; end
		2750: begin l_1 = -33;
				 l_2 = -44; end
		35210: begin l_1 = +33;
				 l_2 = +45; end
		35953: begin l_1 = +33;
				 l_2 = -45; end
		14908: begin l_1 = -33;
				 l_2 = +45; end
		15651: begin l_1 = -33;
				 l_2 = -45; end
		9408: begin l_1 = +33;
				 l_2 = +46; end
		10894: begin l_1 = +33;
				 l_2 = -46; end
		39967: begin l_1 = -33;
				 l_2 = +46; end
		41453: begin l_1 = -33;
				 l_2 = -46; end
		8665: begin l_1 = +33;
				 l_2 = +47; end
		11637: begin l_1 = +33;
				 l_2 = -47; end
		39224: begin l_1 = -33;
				 l_2 = +47; end
		42196: begin l_1 = -33;
				 l_2 = -47; end
		7179: begin l_1 = +33;
				 l_2 = +48; end
		13123: begin l_1 = +33;
				 l_2 = -48; end
		37738: begin l_1 = -33;
				 l_2 = +48; end
		43682: begin l_1 = -33;
				 l_2 = -48; end
		4207: begin l_1 = +33;
				 l_2 = +49; end
		16095: begin l_1 = +33;
				 l_2 = -49; end
		34766: begin l_1 = -33;
				 l_2 = +49; end
		46654: begin l_1 = -33;
				 l_2 = -49; end
		49124: begin l_1 = +33;
				 l_2 = +50; end
		22039: begin l_1 = +33;
				 l_2 = -50; end
		28822: begin l_1 = -33;
				 l_2 = +50; end
		1737: begin l_1 = -33;
				 l_2 = -50; end
		37236: begin l_1 = +33;
				 l_2 = +51; end
		33927: begin l_1 = +33;
				 l_2 = -51; end
		16934: begin l_1 = -33;
				 l_2 = +51; end
		13625: begin l_1 = -33;
				 l_2 = -51; end
		13460: begin l_1 = +33;
				 l_2 = +52; end
		6842: begin l_1 = +33;
				 l_2 = -52; end
		44019: begin l_1 = -33;
				 l_2 = +52; end
		37401: begin l_1 = -33;
				 l_2 = -52; end
		16769: begin l_1 = +33;
				 l_2 = +53; end
		3533: begin l_1 = +33;
				 l_2 = -53; end
		47328: begin l_1 = -33;
				 l_2 = +53; end
		34092: begin l_1 = -33;
				 l_2 = -53; end
		23387: begin l_1 = +33;
				 l_2 = +54; end
		47776: begin l_1 = +33;
				 l_2 = -54; end
		3085: begin l_1 = -33;
				 l_2 = +54; end
		27474: begin l_1 = -33;
				 l_2 = -54; end
		36623: begin l_1 = +33;
				 l_2 = +55; end
		34540: begin l_1 = +33;
				 l_2 = -55; end
		16321: begin l_1 = -33;
				 l_2 = +55; end
		14238: begin l_1 = -33;
				 l_2 = -55; end
		12234: begin l_1 = +33;
				 l_2 = +56; end
		8068: begin l_1 = +33;
				 l_2 = -56; end
		42793: begin l_1 = -33;
				 l_2 = +56; end
		38627: begin l_1 = -33;
				 l_2 = -56; end
		14317: begin l_1 = +33;
				 l_2 = +57; end
		5985: begin l_1 = +33;
				 l_2 = -57; end
		44876: begin l_1 = -33;
				 l_2 = +57; end
		36544: begin l_1 = -33;
				 l_2 = -57; end
		18483: begin l_1 = +33;
				 l_2 = +58; end
		1819: begin l_1 = +33;
				 l_2 = -58; end
		49042: begin l_1 = -33;
				 l_2 = +58; end
		32378: begin l_1 = -33;
				 l_2 = -58; end
		26815: begin l_1 = +33;
				 l_2 = +59; end
		44348: begin l_1 = +33;
				 l_2 = -59; end
		6513: begin l_1 = -33;
				 l_2 = +59; end
		24046: begin l_1 = -33;
				 l_2 = -59; end
		43479: begin l_1 = +33;
				 l_2 = +60; end
		27684: begin l_1 = +33;
				 l_2 = -60; end
		23177: begin l_1 = -33;
				 l_2 = +60; end
		7382: begin l_1 = -33;
				 l_2 = -60; end
		25946: begin l_1 = +33;
				 l_2 = +61; end
		45217: begin l_1 = +33;
				 l_2 = -61; end
		5644: begin l_1 = -33;
				 l_2 = +61; end
		24915: begin l_1 = -33;
				 l_2 = -61; end
		41741: begin l_1 = +33;
				 l_2 = +62; end
		29422: begin l_1 = +33;
				 l_2 = -62; end
		21439: begin l_1 = -33;
				 l_2 = +62; end
		9120: begin l_1 = -33;
				 l_2 = -62; end
		22470: begin l_1 = +33;
				 l_2 = +63; end
		48693: begin l_1 = +33;
				 l_2 = -63; end
		2168: begin l_1 = -33;
				 l_2 = +63; end
		28391: begin l_1 = -33;
				 l_2 = -63; end
		34789: begin l_1 = +33;
				 l_2 = +64; end
		36374: begin l_1 = +33;
				 l_2 = -64; end
		14487: begin l_1 = -33;
				 l_2 = +64; end
		16072: begin l_1 = -33;
				 l_2 = -64; end
		8566: begin l_1 = +33;
				 l_2 = +65; end
		11736: begin l_1 = +33;
				 l_2 = -65; end
		39125: begin l_1 = -33;
				 l_2 = +65; end
		42295: begin l_1 = -33;
				 l_2 = -65; end
		6981: begin l_1 = +33;
				 l_2 = +66; end
		13321: begin l_1 = +33;
				 l_2 = -66; end
		37540: begin l_1 = -33;
				 l_2 = +66; end
		43880: begin l_1 = -33;
				 l_2 = -66; end
		3811: begin l_1 = +33;
				 l_2 = +67; end
		16491: begin l_1 = +33;
				 l_2 = -67; end
		34370: begin l_1 = -33;
				 l_2 = +67; end
		47050: begin l_1 = -33;
				 l_2 = -67; end
		48332: begin l_1 = +33;
				 l_2 = +68; end
		22831: begin l_1 = +33;
				 l_2 = -68; end
		28030: begin l_1 = -33;
				 l_2 = +68; end
		2529: begin l_1 = -33;
				 l_2 = -68; end
		10045: begin l_1 = -34;
				 l_2 = +36; end
		40816: begin l_1 = -34;
				 l_2 = -35; end
		50649: begin l_1 = +34;
				 l_2 = +36; end
		212: begin l_1 = -34;
				 l_2 = -36; end
		30135: begin l_1 = +34;
				 l_2 = +37; end
		10469: begin l_1 = +34;
				 l_2 = -37; end
		40392: begin l_1 = -34;
				 l_2 = +37; end
		20726: begin l_1 = -34;
				 l_2 = -37; end
		39968: begin l_1 = +34;
				 l_2 = +38; end
		636: begin l_1 = +34;
				 l_2 = -38; end
		50225: begin l_1 = -34;
				 l_2 = +38; end
		10893: begin l_1 = -34;
				 l_2 = -38; end
		8773: begin l_1 = +34;
				 l_2 = +39; end
		31831: begin l_1 = +34;
				 l_2 = -39; end
		19030: begin l_1 = -34;
				 l_2 = +39; end
		42088: begin l_1 = -34;
				 l_2 = -39; end
		48105: begin l_1 = +34;
				 l_2 = +40; end
		43360: begin l_1 = +34;
				 l_2 = -40; end
		7501: begin l_1 = -34;
				 l_2 = +40; end
		2756: begin l_1 = -34;
				 l_2 = -40; end
		25047: begin l_1 = +34;
				 l_2 = +41; end
		15557: begin l_1 = +34;
				 l_2 = -41; end
		35304: begin l_1 = -34;
				 l_2 = +41; end
		25814: begin l_1 = -34;
				 l_2 = -41; end
		29792: begin l_1 = +34;
				 l_2 = +42; end
		10812: begin l_1 = +34;
				 l_2 = -42; end
		40049: begin l_1 = -34;
				 l_2 = +42; end
		21069: begin l_1 = -34;
				 l_2 = -42; end
		39282: begin l_1 = +34;
				 l_2 = +43; end
		1322: begin l_1 = +34;
				 l_2 = -43; end
		49539: begin l_1 = -34;
				 l_2 = +43; end
		11579: begin l_1 = -34;
				 l_2 = -43; end
		7401: begin l_1 = +34;
				 l_2 = +44; end
		33203: begin l_1 = +34;
				 l_2 = -44; end
		17658: begin l_1 = -34;
				 l_2 = +44; end
		43460: begin l_1 = -34;
				 l_2 = -44; end
		45361: begin l_1 = +34;
				 l_2 = +45; end
		46104: begin l_1 = +34;
				 l_2 = -45; end
		4757: begin l_1 = -34;
				 l_2 = +45; end
		5500: begin l_1 = -34;
				 l_2 = -45; end
		19559: begin l_1 = +34;
				 l_2 = +46; end
		21045: begin l_1 = +34;
				 l_2 = -46; end
		29816: begin l_1 = -34;
				 l_2 = +46; end
		31302: begin l_1 = -34;
				 l_2 = -46; end
		18816: begin l_1 = +34;
				 l_2 = +47; end
		21788: begin l_1 = +34;
				 l_2 = -47; end
		29073: begin l_1 = -34;
				 l_2 = +47; end
		32045: begin l_1 = -34;
				 l_2 = -47; end
		17330: begin l_1 = +34;
				 l_2 = +48; end
		23274: begin l_1 = +34;
				 l_2 = -48; end
		27587: begin l_1 = -34;
				 l_2 = +48; end
		33531: begin l_1 = -34;
				 l_2 = -48; end
		14358: begin l_1 = +34;
				 l_2 = +49; end
		26246: begin l_1 = +34;
				 l_2 = -49; end
		24615: begin l_1 = -34;
				 l_2 = +49; end
		36503: begin l_1 = -34;
				 l_2 = -49; end
		8414: begin l_1 = +34;
				 l_2 = +50; end
		32190: begin l_1 = +34;
				 l_2 = -50; end
		18671: begin l_1 = -34;
				 l_2 = +50; end
		42447: begin l_1 = -34;
				 l_2 = -50; end
		47387: begin l_1 = +34;
				 l_2 = +51; end
		44078: begin l_1 = +34;
				 l_2 = -51; end
		6783: begin l_1 = -34;
				 l_2 = +51; end
		3474: begin l_1 = -34;
				 l_2 = -51; end
		23611: begin l_1 = +34;
				 l_2 = +52; end
		16993: begin l_1 = +34;
				 l_2 = -52; end
		33868: begin l_1 = -34;
				 l_2 = +52; end
		27250: begin l_1 = -34;
				 l_2 = -52; end
		26920: begin l_1 = +34;
				 l_2 = +53; end
		13684: begin l_1 = +34;
				 l_2 = -53; end
		37177: begin l_1 = -34;
				 l_2 = +53; end
		23941: begin l_1 = -34;
				 l_2 = -53; end
		33538: begin l_1 = +34;
				 l_2 = +54; end
		7066: begin l_1 = +34;
				 l_2 = -54; end
		43795: begin l_1 = -34;
				 l_2 = +54; end
		17323: begin l_1 = -34;
				 l_2 = -54; end
		46774: begin l_1 = +34;
				 l_2 = +55; end
		44691: begin l_1 = +34;
				 l_2 = -55; end
		6170: begin l_1 = -34;
				 l_2 = +55; end
		4087: begin l_1 = -34;
				 l_2 = -55; end
		22385: begin l_1 = +34;
				 l_2 = +56; end
		18219: begin l_1 = +34;
				 l_2 = -56; end
		32642: begin l_1 = -34;
				 l_2 = +56; end
		28476: begin l_1 = -34;
				 l_2 = -56; end
		24468: begin l_1 = +34;
				 l_2 = +57; end
		16136: begin l_1 = +34;
				 l_2 = -57; end
		34725: begin l_1 = -34;
				 l_2 = +57; end
		26393: begin l_1 = -34;
				 l_2 = -57; end
		28634: begin l_1 = +34;
				 l_2 = +58; end
		11970: begin l_1 = +34;
				 l_2 = -58; end
		38891: begin l_1 = -34;
				 l_2 = +58; end
		22227: begin l_1 = -34;
				 l_2 = -58; end
		36966: begin l_1 = +34;
				 l_2 = +59; end
		3638: begin l_1 = +34;
				 l_2 = -59; end
		47223: begin l_1 = -34;
				 l_2 = +59; end
		13895: begin l_1 = -34;
				 l_2 = -59; end
		2769: begin l_1 = +34;
				 l_2 = +60; end
		37835: begin l_1 = +34;
				 l_2 = -60; end
		13026: begin l_1 = -34;
				 l_2 = +60; end
		48092: begin l_1 = -34;
				 l_2 = -60; end
		36097: begin l_1 = +34;
				 l_2 = +61; end
		4507: begin l_1 = +34;
				 l_2 = -61; end
		46354: begin l_1 = -34;
				 l_2 = +61; end
		14764: begin l_1 = -34;
				 l_2 = -61; end
		1031: begin l_1 = +34;
				 l_2 = +62; end
		39573: begin l_1 = +34;
				 l_2 = -62; end
		11288: begin l_1 = -34;
				 l_2 = +62; end
		49830: begin l_1 = -34;
				 l_2 = -62; end
		32621: begin l_1 = +34;
				 l_2 = +63; end
		7983: begin l_1 = +34;
				 l_2 = -63; end
		42878: begin l_1 = -34;
				 l_2 = +63; end
		18240: begin l_1 = -34;
				 l_2 = -63; end
		44940: begin l_1 = +34;
				 l_2 = +64; end
		46525: begin l_1 = +34;
				 l_2 = -64; end
		4336: begin l_1 = -34;
				 l_2 = +64; end
		5921: begin l_1 = -34;
				 l_2 = -64; end
		18717: begin l_1 = +34;
				 l_2 = +65; end
		21887: begin l_1 = +34;
				 l_2 = -65; end
		28974: begin l_1 = -34;
				 l_2 = +65; end
		32144: begin l_1 = -34;
				 l_2 = -65; end
		17132: begin l_1 = +34;
				 l_2 = +66; end
		23472: begin l_1 = +34;
				 l_2 = -66; end
		27389: begin l_1 = -34;
				 l_2 = +66; end
		33729: begin l_1 = -34;
				 l_2 = -66; end
		13962: begin l_1 = +34;
				 l_2 = +67; end
		26642: begin l_1 = +34;
				 l_2 = -67; end
		24219: begin l_1 = -34;
				 l_2 = +67; end
		36899: begin l_1 = -34;
				 l_2 = -67; end
		7622: begin l_1 = +34;
				 l_2 = +68; end
		32982: begin l_1 = +34;
				 l_2 = -68; end
		17879: begin l_1 = -34;
				 l_2 = +68; end
		43239: begin l_1 = -34;
				 l_2 = -68; end
		20090: begin l_1 = -35;
				 l_2 = +37; end
		30771: begin l_1 = -35;
				 l_2 = -36; end
		50437: begin l_1 = +35;
				 l_2 = +37; end
		424: begin l_1 = -35;
				 l_2 = -37; end
		9409: begin l_1 = +35;
				 l_2 = +38; end
		20938: begin l_1 = +35;
				 l_2 = -38; end
		29923: begin l_1 = -35;
				 l_2 = +38; end
		41452: begin l_1 = -35;
				 l_2 = -38; end
		29075: begin l_1 = +35;
				 l_2 = +39; end
		1272: begin l_1 = +35;
				 l_2 = -39; end
		49589: begin l_1 = -35;
				 l_2 = +39; end
		21786: begin l_1 = -35;
				 l_2 = -39; end
		17546: begin l_1 = +35;
				 l_2 = +40; end
		12801: begin l_1 = +35;
				 l_2 = -40; end
		38060: begin l_1 = -35;
				 l_2 = +40; end
		33315: begin l_1 = -35;
				 l_2 = -40; end
		45349: begin l_1 = +35;
				 l_2 = +41; end
		35859: begin l_1 = +35;
				 l_2 = -41; end
		15002: begin l_1 = -35;
				 l_2 = +41; end
		5512: begin l_1 = -35;
				 l_2 = -41; end
		50094: begin l_1 = +35;
				 l_2 = +42; end
		31114: begin l_1 = +35;
				 l_2 = -42; end
		19747: begin l_1 = -35;
				 l_2 = +42; end
		767: begin l_1 = -35;
				 l_2 = -42; end
		8723: begin l_1 = +35;
				 l_2 = +43; end
		21624: begin l_1 = +35;
				 l_2 = -43; end
		29237: begin l_1 = -35;
				 l_2 = +43; end
		42138: begin l_1 = -35;
				 l_2 = -43; end
		27703: begin l_1 = +35;
				 l_2 = +44; end
		2644: begin l_1 = +35;
				 l_2 = -44; end
		48217: begin l_1 = -35;
				 l_2 = +44; end
		23158: begin l_1 = -35;
				 l_2 = -44; end
		14802: begin l_1 = +35;
				 l_2 = +45; end
		15545: begin l_1 = +35;
				 l_2 = -45; end
		35316: begin l_1 = -35;
				 l_2 = +45; end
		36059: begin l_1 = -35;
				 l_2 = -45; end
		39861: begin l_1 = +35;
				 l_2 = +46; end
		41347: begin l_1 = +35;
				 l_2 = -46; end
		9514: begin l_1 = -35;
				 l_2 = +46; end
		11000: begin l_1 = -35;
				 l_2 = -46; end
		39118: begin l_1 = +35;
				 l_2 = +47; end
		42090: begin l_1 = +35;
				 l_2 = -47; end
		8771: begin l_1 = -35;
				 l_2 = +47; end
		11743: begin l_1 = -35;
				 l_2 = -47; end
		37632: begin l_1 = +35;
				 l_2 = +48; end
		43576: begin l_1 = +35;
				 l_2 = -48; end
		7285: begin l_1 = -35;
				 l_2 = +48; end
		13229: begin l_1 = -35;
				 l_2 = -48; end
		34660: begin l_1 = +35;
				 l_2 = +49; end
		46548: begin l_1 = +35;
				 l_2 = -49; end
		4313: begin l_1 = -35;
				 l_2 = +49; end
		16201: begin l_1 = -35;
				 l_2 = -49; end
		28716: begin l_1 = +35;
				 l_2 = +50; end
		1631: begin l_1 = +35;
				 l_2 = -50; end
		49230: begin l_1 = -35;
				 l_2 = +50; end
		22145: begin l_1 = -35;
				 l_2 = -50; end
		16828: begin l_1 = +35;
				 l_2 = +51; end
		13519: begin l_1 = +35;
				 l_2 = -51; end
		37342: begin l_1 = -35;
				 l_2 = +51; end
		34033: begin l_1 = -35;
				 l_2 = -51; end
		43913: begin l_1 = +35;
				 l_2 = +52; end
		37295: begin l_1 = +35;
				 l_2 = -52; end
		13566: begin l_1 = -35;
				 l_2 = +52; end
		6948: begin l_1 = -35;
				 l_2 = -52; end
		47222: begin l_1 = +35;
				 l_2 = +53; end
		33986: begin l_1 = +35;
				 l_2 = -53; end
		16875: begin l_1 = -35;
				 l_2 = +53; end
		3639: begin l_1 = -35;
				 l_2 = -53; end
		2979: begin l_1 = +35;
				 l_2 = +54; end
		27368: begin l_1 = +35;
				 l_2 = -54; end
		23493: begin l_1 = -35;
				 l_2 = +54; end
		47882: begin l_1 = -35;
				 l_2 = -54; end
		16215: begin l_1 = +35;
				 l_2 = +55; end
		14132: begin l_1 = +35;
				 l_2 = -55; end
		36729: begin l_1 = -35;
				 l_2 = +55; end
		34646: begin l_1 = -35;
				 l_2 = -55; end
		42687: begin l_1 = +35;
				 l_2 = +56; end
		38521: begin l_1 = +35;
				 l_2 = -56; end
		12340: begin l_1 = -35;
				 l_2 = +56; end
		8174: begin l_1 = -35;
				 l_2 = -56; end
		44770: begin l_1 = +35;
				 l_2 = +57; end
		36438: begin l_1 = +35;
				 l_2 = -57; end
		14423: begin l_1 = -35;
				 l_2 = +57; end
		6091: begin l_1 = -35;
				 l_2 = -57; end
		48936: begin l_1 = +35;
				 l_2 = +58; end
		32272: begin l_1 = +35;
				 l_2 = -58; end
		18589: begin l_1 = -35;
				 l_2 = +58; end
		1925: begin l_1 = -35;
				 l_2 = -58; end
		6407: begin l_1 = +35;
				 l_2 = +59; end
		23940: begin l_1 = +35;
				 l_2 = -59; end
		26921: begin l_1 = -35;
				 l_2 = +59; end
		44454: begin l_1 = -35;
				 l_2 = -59; end
		23071: begin l_1 = +35;
				 l_2 = +60; end
		7276: begin l_1 = +35;
				 l_2 = -60; end
		43585: begin l_1 = -35;
				 l_2 = +60; end
		27790: begin l_1 = -35;
				 l_2 = -60; end
		5538: begin l_1 = +35;
				 l_2 = +61; end
		24809: begin l_1 = +35;
				 l_2 = -61; end
		26052: begin l_1 = -35;
				 l_2 = +61; end
		45323: begin l_1 = -35;
				 l_2 = -61; end
		21333: begin l_1 = +35;
				 l_2 = +62; end
		9014: begin l_1 = +35;
				 l_2 = -62; end
		41847: begin l_1 = -35;
				 l_2 = +62; end
		29528: begin l_1 = -35;
				 l_2 = -62; end
		2062: begin l_1 = +35;
				 l_2 = +63; end
		28285: begin l_1 = +35;
				 l_2 = -63; end
		22576: begin l_1 = -35;
				 l_2 = +63; end
		48799: begin l_1 = -35;
				 l_2 = -63; end
		14381: begin l_1 = +35;
				 l_2 = +64; end
		15966: begin l_1 = +35;
				 l_2 = -64; end
		34895: begin l_1 = -35;
				 l_2 = +64; end
		36480: begin l_1 = -35;
				 l_2 = -64; end
		39019: begin l_1 = +35;
				 l_2 = +65; end
		42189: begin l_1 = +35;
				 l_2 = -65; end
		8672: begin l_1 = -35;
				 l_2 = +65; end
		11842: begin l_1 = -35;
				 l_2 = -65; end
		37434: begin l_1 = +35;
				 l_2 = +66; end
		43774: begin l_1 = +35;
				 l_2 = -66; end
		7087: begin l_1 = -35;
				 l_2 = +66; end
		13427: begin l_1 = -35;
				 l_2 = -66; end
		34264: begin l_1 = +35;
				 l_2 = +67; end
		46944: begin l_1 = +35;
				 l_2 = -67; end
		3917: begin l_1 = -35;
				 l_2 = +67; end
		16597: begin l_1 = -35;
				 l_2 = -67; end
		27924: begin l_1 = +35;
				 l_2 = +68; end
		2423: begin l_1 = +35;
				 l_2 = -68; end
		48438: begin l_1 = -35;
				 l_2 = +68; end
		22937: begin l_1 = -35;
				 l_2 = -68; end
		40180: begin l_1 = -36;
				 l_2 = +38; end
		10681: begin l_1 = -36;
				 l_2 = -37; end
		50013: begin l_1 = +36;
				 l_2 = +38; end
		848: begin l_1 = -36;
				 l_2 = -38; end
		18818: begin l_1 = +36;
				 l_2 = +39; end
		41876: begin l_1 = +36;
				 l_2 = -39; end
		8985: begin l_1 = -36;
				 l_2 = +39; end
		32043: begin l_1 = -36;
				 l_2 = -39; end
		7289: begin l_1 = +36;
				 l_2 = +40; end
		2544: begin l_1 = +36;
				 l_2 = -40; end
		48317: begin l_1 = -36;
				 l_2 = +40; end
		43572: begin l_1 = -36;
				 l_2 = -40; end
		35092: begin l_1 = +36;
				 l_2 = +41; end
		25602: begin l_1 = +36;
				 l_2 = -41; end
		25259: begin l_1 = -36;
				 l_2 = +41; end
		15769: begin l_1 = -36;
				 l_2 = -41; end
		39837: begin l_1 = +36;
				 l_2 = +42; end
		20857: begin l_1 = +36;
				 l_2 = -42; end
		30004: begin l_1 = -36;
				 l_2 = +42; end
		11024: begin l_1 = -36;
				 l_2 = -42; end
		49327: begin l_1 = +36;
				 l_2 = +43; end
		11367: begin l_1 = +36;
				 l_2 = -43; end
		39494: begin l_1 = -36;
				 l_2 = +43; end
		1534: begin l_1 = -36;
				 l_2 = -43; end
		17446: begin l_1 = +36;
				 l_2 = +44; end
		43248: begin l_1 = +36;
				 l_2 = -44; end
		7613: begin l_1 = -36;
				 l_2 = +44; end
		33415: begin l_1 = -36;
				 l_2 = -44; end
		4545: begin l_1 = +36;
				 l_2 = +45; end
		5288: begin l_1 = +36;
				 l_2 = -45; end
		45573: begin l_1 = -36;
				 l_2 = +45; end
		46316: begin l_1 = -36;
				 l_2 = -45; end
		29604: begin l_1 = +36;
				 l_2 = +46; end
		31090: begin l_1 = +36;
				 l_2 = -46; end
		19771: begin l_1 = -36;
				 l_2 = +46; end
		21257: begin l_1 = -36;
				 l_2 = -46; end
		28861: begin l_1 = +36;
				 l_2 = +47; end
		31833: begin l_1 = +36;
				 l_2 = -47; end
		19028: begin l_1 = -36;
				 l_2 = +47; end
		22000: begin l_1 = -36;
				 l_2 = -47; end
		27375: begin l_1 = +36;
				 l_2 = +48; end
		33319: begin l_1 = +36;
				 l_2 = -48; end
		17542: begin l_1 = -36;
				 l_2 = +48; end
		23486: begin l_1 = -36;
				 l_2 = -48; end
		24403: begin l_1 = +36;
				 l_2 = +49; end
		36291: begin l_1 = +36;
				 l_2 = -49; end
		14570: begin l_1 = -36;
				 l_2 = +49; end
		26458: begin l_1 = -36;
				 l_2 = -49; end
		18459: begin l_1 = +36;
				 l_2 = +50; end
		42235: begin l_1 = +36;
				 l_2 = -50; end
		8626: begin l_1 = -36;
				 l_2 = +50; end
		32402: begin l_1 = -36;
				 l_2 = -50; end
		6571: begin l_1 = +36;
				 l_2 = +51; end
		3262: begin l_1 = +36;
				 l_2 = -51; end
		47599: begin l_1 = -36;
				 l_2 = +51; end
		44290: begin l_1 = -36;
				 l_2 = -51; end
		33656: begin l_1 = +36;
				 l_2 = +52; end
		27038: begin l_1 = +36;
				 l_2 = -52; end
		23823: begin l_1 = -36;
				 l_2 = +52; end
		17205: begin l_1 = -36;
				 l_2 = -52; end
		36965: begin l_1 = +36;
				 l_2 = +53; end
		23729: begin l_1 = +36;
				 l_2 = -53; end
		27132: begin l_1 = -36;
				 l_2 = +53; end
		13896: begin l_1 = -36;
				 l_2 = -53; end
		43583: begin l_1 = +36;
				 l_2 = +54; end
		17111: begin l_1 = +36;
				 l_2 = -54; end
		33750: begin l_1 = -36;
				 l_2 = +54; end
		7278: begin l_1 = -36;
				 l_2 = -54; end
		5958: begin l_1 = +36;
				 l_2 = +55; end
		3875: begin l_1 = +36;
				 l_2 = -55; end
		46986: begin l_1 = -36;
				 l_2 = +55; end
		44903: begin l_1 = -36;
				 l_2 = -55; end
		32430: begin l_1 = +36;
				 l_2 = +56; end
		28264: begin l_1 = +36;
				 l_2 = -56; end
		22597: begin l_1 = -36;
				 l_2 = +56; end
		18431: begin l_1 = -36;
				 l_2 = -56; end
		34513: begin l_1 = +36;
				 l_2 = +57; end
		26181: begin l_1 = +36;
				 l_2 = -57; end
		24680: begin l_1 = -36;
				 l_2 = +57; end
		16348: begin l_1 = -36;
				 l_2 = -57; end
		38679: begin l_1 = +36;
				 l_2 = +58; end
		22015: begin l_1 = +36;
				 l_2 = -58; end
		28846: begin l_1 = -36;
				 l_2 = +58; end
		12182: begin l_1 = -36;
				 l_2 = -58; end
		47011: begin l_1 = +36;
				 l_2 = +59; end
		13683: begin l_1 = +36;
				 l_2 = -59; end
		37178: begin l_1 = -36;
				 l_2 = +59; end
		3850: begin l_1 = -36;
				 l_2 = -59; end
		12814: begin l_1 = +36;
				 l_2 = +60; end
		47880: begin l_1 = +36;
				 l_2 = -60; end
		2981: begin l_1 = -36;
				 l_2 = +60; end
		38047: begin l_1 = -36;
				 l_2 = -60; end
		46142: begin l_1 = +36;
				 l_2 = +61; end
		14552: begin l_1 = +36;
				 l_2 = -61; end
		36309: begin l_1 = -36;
				 l_2 = +61; end
		4719: begin l_1 = -36;
				 l_2 = -61; end
		11076: begin l_1 = +36;
				 l_2 = +62; end
		49618: begin l_1 = +36;
				 l_2 = -62; end
		1243: begin l_1 = -36;
				 l_2 = +62; end
		39785: begin l_1 = -36;
				 l_2 = -62; end
		42666: begin l_1 = +36;
				 l_2 = +63; end
		18028: begin l_1 = +36;
				 l_2 = -63; end
		32833: begin l_1 = -36;
				 l_2 = +63; end
		8195: begin l_1 = -36;
				 l_2 = -63; end
		4124: begin l_1 = +36;
				 l_2 = +64; end
		5709: begin l_1 = +36;
				 l_2 = -64; end
		45152: begin l_1 = -36;
				 l_2 = +64; end
		46737: begin l_1 = -36;
				 l_2 = -64; end
		28762: begin l_1 = +36;
				 l_2 = +65; end
		31932: begin l_1 = +36;
				 l_2 = -65; end
		18929: begin l_1 = -36;
				 l_2 = +65; end
		22099: begin l_1 = -36;
				 l_2 = -65; end
		27177: begin l_1 = +36;
				 l_2 = +66; end
		33517: begin l_1 = +36;
				 l_2 = -66; end
		17344: begin l_1 = -36;
				 l_2 = +66; end
		23684: begin l_1 = -36;
				 l_2 = -66; end
		24007: begin l_1 = +36;
				 l_2 = +67; end
		36687: begin l_1 = +36;
				 l_2 = -67; end
		14174: begin l_1 = -36;
				 l_2 = +67; end
		26854: begin l_1 = -36;
				 l_2 = -67; end
		17667: begin l_1 = +36;
				 l_2 = +68; end
		43027: begin l_1 = +36;
				 l_2 = -68; end
		7834: begin l_1 = -36;
				 l_2 = +68; end
		33194: begin l_1 = -36;
				 l_2 = -68; end
		29499: begin l_1 = -37;
				 l_2 = +39; end
		21362: begin l_1 = -37;
				 l_2 = -38; end
		49165: begin l_1 = +37;
				 l_2 = +39; end
		1696: begin l_1 = -37;
				 l_2 = -39; end
		37636: begin l_1 = +37;
				 l_2 = +40; end
		32891: begin l_1 = +37;
				 l_2 = -40; end
		17970: begin l_1 = -37;
				 l_2 = +40; end
		13225: begin l_1 = -37;
				 l_2 = -40; end
		14578: begin l_1 = +37;
				 l_2 = +41; end
		5088: begin l_1 = +37;
				 l_2 = -41; end
		45773: begin l_1 = -37;
				 l_2 = +41; end
		36283: begin l_1 = -37;
				 l_2 = -41; end
		19323: begin l_1 = +37;
				 l_2 = +42; end
		343: begin l_1 = +37;
				 l_2 = -42; end
		50518: begin l_1 = -37;
				 l_2 = +42; end
		31538: begin l_1 = -37;
				 l_2 = -42; end
		28813: begin l_1 = +37;
				 l_2 = +43; end
		41714: begin l_1 = +37;
				 l_2 = -43; end
		9147: begin l_1 = -37;
				 l_2 = +43; end
		22048: begin l_1 = -37;
				 l_2 = -43; end
		47793: begin l_1 = +37;
				 l_2 = +44; end
		22734: begin l_1 = +37;
				 l_2 = -44; end
		28127: begin l_1 = -37;
				 l_2 = +44; end
		3068: begin l_1 = -37;
				 l_2 = -44; end
		34892: begin l_1 = +37;
				 l_2 = +45; end
		35635: begin l_1 = +37;
				 l_2 = -45; end
		15226: begin l_1 = -37;
				 l_2 = +45; end
		15969: begin l_1 = -37;
				 l_2 = -45; end
		9090: begin l_1 = +37;
				 l_2 = +46; end
		10576: begin l_1 = +37;
				 l_2 = -46; end
		40285: begin l_1 = -37;
				 l_2 = +46; end
		41771: begin l_1 = -37;
				 l_2 = -46; end
		8347: begin l_1 = +37;
				 l_2 = +47; end
		11319: begin l_1 = +37;
				 l_2 = -47; end
		39542: begin l_1 = -37;
				 l_2 = +47; end
		42514: begin l_1 = -37;
				 l_2 = -47; end
		6861: begin l_1 = +37;
				 l_2 = +48; end
		12805: begin l_1 = +37;
				 l_2 = -48; end
		38056: begin l_1 = -37;
				 l_2 = +48; end
		44000: begin l_1 = -37;
				 l_2 = -48; end
		3889: begin l_1 = +37;
				 l_2 = +49; end
		15777: begin l_1 = +37;
				 l_2 = -49; end
		35084: begin l_1 = -37;
				 l_2 = +49; end
		46972: begin l_1 = -37;
				 l_2 = -49; end
		48806: begin l_1 = +37;
				 l_2 = +50; end
		21721: begin l_1 = +37;
				 l_2 = -50; end
		29140: begin l_1 = -37;
				 l_2 = +50; end
		2055: begin l_1 = -37;
				 l_2 = -50; end
		36918: begin l_1 = +37;
				 l_2 = +51; end
		33609: begin l_1 = +37;
				 l_2 = -51; end
		17252: begin l_1 = -37;
				 l_2 = +51; end
		13943: begin l_1 = -37;
				 l_2 = -51; end
		13142: begin l_1 = +37;
				 l_2 = +52; end
		6524: begin l_1 = +37;
				 l_2 = -52; end
		44337: begin l_1 = -37;
				 l_2 = +52; end
		37719: begin l_1 = -37;
				 l_2 = -52; end
		16451: begin l_1 = +37;
				 l_2 = +53; end
		3215: begin l_1 = +37;
				 l_2 = -53; end
		47646: begin l_1 = -37;
				 l_2 = +53; end
		34410: begin l_1 = -37;
				 l_2 = -53; end
		23069: begin l_1 = +37;
				 l_2 = +54; end
		47458: begin l_1 = +37;
				 l_2 = -54; end
		3403: begin l_1 = -37;
				 l_2 = +54; end
		27792: begin l_1 = -37;
				 l_2 = -54; end
		36305: begin l_1 = +37;
				 l_2 = +55; end
		34222: begin l_1 = +37;
				 l_2 = -55; end
		16639: begin l_1 = -37;
				 l_2 = +55; end
		14556: begin l_1 = -37;
				 l_2 = -55; end
		11916: begin l_1 = +37;
				 l_2 = +56; end
		7750: begin l_1 = +37;
				 l_2 = -56; end
		43111: begin l_1 = -37;
				 l_2 = +56; end
		38945: begin l_1 = -37;
				 l_2 = -56; end
		13999: begin l_1 = +37;
				 l_2 = +57; end
		5667: begin l_1 = +37;
				 l_2 = -57; end
		45194: begin l_1 = -37;
				 l_2 = +57; end
		36862: begin l_1 = -37;
				 l_2 = -57; end
		18165: begin l_1 = +37;
				 l_2 = +58; end
		1501: begin l_1 = +37;
				 l_2 = -58; end
		49360: begin l_1 = -37;
				 l_2 = +58; end
		32696: begin l_1 = -37;
				 l_2 = -58; end
		26497: begin l_1 = +37;
				 l_2 = +59; end
		44030: begin l_1 = +37;
				 l_2 = -59; end
		6831: begin l_1 = -37;
				 l_2 = +59; end
		24364: begin l_1 = -37;
				 l_2 = -59; end
		43161: begin l_1 = +37;
				 l_2 = +60; end
		27366: begin l_1 = +37;
				 l_2 = -60; end
		23495: begin l_1 = -37;
				 l_2 = +60; end
		7700: begin l_1 = -37;
				 l_2 = -60; end
		25628: begin l_1 = +37;
				 l_2 = +61; end
		44899: begin l_1 = +37;
				 l_2 = -61; end
		5962: begin l_1 = -37;
				 l_2 = +61; end
		25233: begin l_1 = -37;
				 l_2 = -61; end
		41423: begin l_1 = +37;
				 l_2 = +62; end
		29104: begin l_1 = +37;
				 l_2 = -62; end
		21757: begin l_1 = -37;
				 l_2 = +62; end
		9438: begin l_1 = -37;
				 l_2 = -62; end
		22152: begin l_1 = +37;
				 l_2 = +63; end
		48375: begin l_1 = +37;
				 l_2 = -63; end
		2486: begin l_1 = -37;
				 l_2 = +63; end
		28709: begin l_1 = -37;
				 l_2 = -63; end
		34471: begin l_1 = +37;
				 l_2 = +64; end
		36056: begin l_1 = +37;
				 l_2 = -64; end
		14805: begin l_1 = -37;
				 l_2 = +64; end
		16390: begin l_1 = -37;
				 l_2 = -64; end
		8248: begin l_1 = +37;
				 l_2 = +65; end
		11418: begin l_1 = +37;
				 l_2 = -65; end
		39443: begin l_1 = -37;
				 l_2 = +65; end
		42613: begin l_1 = -37;
				 l_2 = -65; end
		6663: begin l_1 = +37;
				 l_2 = +66; end
		13003: begin l_1 = +37;
				 l_2 = -66; end
		37858: begin l_1 = -37;
				 l_2 = +66; end
		44198: begin l_1 = -37;
				 l_2 = -66; end
		3493: begin l_1 = +37;
				 l_2 = +67; end
		16173: begin l_1 = +37;
				 l_2 = -67; end
		34688: begin l_1 = -37;
				 l_2 = +67; end
		47368: begin l_1 = -37;
				 l_2 = -67; end
		48014: begin l_1 = +37;
				 l_2 = +68; end
		22513: begin l_1 = +37;
				 l_2 = -68; end
		28348: begin l_1 = -37;
				 l_2 = +68; end
		2847: begin l_1 = -37;
				 l_2 = -68; end
		8137: begin l_1 = -38;
				 l_2 = +40; end
		42724: begin l_1 = -38;
				 l_2 = -39; end
		47469: begin l_1 = +38;
				 l_2 = +40; end
		3392: begin l_1 = -38;
				 l_2 = -40; end
		24411: begin l_1 = +38;
				 l_2 = +41; end
		14921: begin l_1 = +38;
				 l_2 = -41; end
		35940: begin l_1 = -38;
				 l_2 = +41; end
		26450: begin l_1 = -38;
				 l_2 = -41; end
		29156: begin l_1 = +38;
				 l_2 = +42; end
		10176: begin l_1 = +38;
				 l_2 = -42; end
		40685: begin l_1 = -38;
				 l_2 = +42; end
		21705: begin l_1 = -38;
				 l_2 = -42; end
		38646: begin l_1 = +38;
				 l_2 = +43; end
		686: begin l_1 = +38;
				 l_2 = -43; end
		50175: begin l_1 = -38;
				 l_2 = +43; end
		12215: begin l_1 = -38;
				 l_2 = -43; end
		6765: begin l_1 = +38;
				 l_2 = +44; end
		32567: begin l_1 = +38;
				 l_2 = -44; end
		18294: begin l_1 = -38;
				 l_2 = +44; end
		44096: begin l_1 = -38;
				 l_2 = -44; end
		44725: begin l_1 = +38;
				 l_2 = +45; end
		45468: begin l_1 = +38;
				 l_2 = -45; end
		5393: begin l_1 = -38;
				 l_2 = +45; end
		6136: begin l_1 = -38;
				 l_2 = -45; end
		18923: begin l_1 = +38;
				 l_2 = +46; end
		20409: begin l_1 = +38;
				 l_2 = -46; end
		30452: begin l_1 = -38;
				 l_2 = +46; end
		31938: begin l_1 = -38;
				 l_2 = -46; end
		18180: begin l_1 = +38;
				 l_2 = +47; end
		21152: begin l_1 = +38;
				 l_2 = -47; end
		29709: begin l_1 = -38;
				 l_2 = +47; end
		32681: begin l_1 = -38;
				 l_2 = -47; end
		16694: begin l_1 = +38;
				 l_2 = +48; end
		22638: begin l_1 = +38;
				 l_2 = -48; end
		28223: begin l_1 = -38;
				 l_2 = +48; end
		34167: begin l_1 = -38;
				 l_2 = -48; end
		13722: begin l_1 = +38;
				 l_2 = +49; end
		25610: begin l_1 = +38;
				 l_2 = -49; end
		25251: begin l_1 = -38;
				 l_2 = +49; end
		37139: begin l_1 = -38;
				 l_2 = -49; end
		7778: begin l_1 = +38;
				 l_2 = +50; end
		31554: begin l_1 = +38;
				 l_2 = -50; end
		19307: begin l_1 = -38;
				 l_2 = +50; end
		43083: begin l_1 = -38;
				 l_2 = -50; end
		46751: begin l_1 = +38;
				 l_2 = +51; end
		43442: begin l_1 = +38;
				 l_2 = -51; end
		7419: begin l_1 = -38;
				 l_2 = +51; end
		4110: begin l_1 = -38;
				 l_2 = -51; end
		22975: begin l_1 = +38;
				 l_2 = +52; end
		16357: begin l_1 = +38;
				 l_2 = -52; end
		34504: begin l_1 = -38;
				 l_2 = +52; end
		27886: begin l_1 = -38;
				 l_2 = -52; end
		26284: begin l_1 = +38;
				 l_2 = +53; end
		13048: begin l_1 = +38;
				 l_2 = -53; end
		37813: begin l_1 = -38;
				 l_2 = +53; end
		24577: begin l_1 = -38;
				 l_2 = -53; end
		32902: begin l_1 = +38;
				 l_2 = +54; end
		6430: begin l_1 = +38;
				 l_2 = -54; end
		44431: begin l_1 = -38;
				 l_2 = +54; end
		17959: begin l_1 = -38;
				 l_2 = -54; end
		46138: begin l_1 = +38;
				 l_2 = +55; end
		44055: begin l_1 = +38;
				 l_2 = -55; end
		6806: begin l_1 = -38;
				 l_2 = +55; end
		4723: begin l_1 = -38;
				 l_2 = -55; end
		21749: begin l_1 = +38;
				 l_2 = +56; end
		17583: begin l_1 = +38;
				 l_2 = -56; end
		33278: begin l_1 = -38;
				 l_2 = +56; end
		29112: begin l_1 = -38;
				 l_2 = -56; end
		23832: begin l_1 = +38;
				 l_2 = +57; end
		15500: begin l_1 = +38;
				 l_2 = -57; end
		35361: begin l_1 = -38;
				 l_2 = +57; end
		27029: begin l_1 = -38;
				 l_2 = -57; end
		27998: begin l_1 = +38;
				 l_2 = +58; end
		11334: begin l_1 = +38;
				 l_2 = -58; end
		39527: begin l_1 = -38;
				 l_2 = +58; end
		22863: begin l_1 = -38;
				 l_2 = -58; end
		36330: begin l_1 = +38;
				 l_2 = +59; end
		3002: begin l_1 = +38;
				 l_2 = -59; end
		47859: begin l_1 = -38;
				 l_2 = +59; end
		14531: begin l_1 = -38;
				 l_2 = -59; end
		2133: begin l_1 = +38;
				 l_2 = +60; end
		37199: begin l_1 = +38;
				 l_2 = -60; end
		13662: begin l_1 = -38;
				 l_2 = +60; end
		48728: begin l_1 = -38;
				 l_2 = -60; end
		35461: begin l_1 = +38;
				 l_2 = +61; end
		3871: begin l_1 = +38;
				 l_2 = -61; end
		46990: begin l_1 = -38;
				 l_2 = +61; end
		15400: begin l_1 = -38;
				 l_2 = -61; end
		395: begin l_1 = +38;
				 l_2 = +62; end
		38937: begin l_1 = +38;
				 l_2 = -62; end
		11924: begin l_1 = -38;
				 l_2 = +62; end
		50466: begin l_1 = -38;
				 l_2 = -62; end
		31985: begin l_1 = +38;
				 l_2 = +63; end
		7347: begin l_1 = +38;
				 l_2 = -63; end
		43514: begin l_1 = -38;
				 l_2 = +63; end
		18876: begin l_1 = -38;
				 l_2 = -63; end
		44304: begin l_1 = +38;
				 l_2 = +64; end
		45889: begin l_1 = +38;
				 l_2 = -64; end
		4972: begin l_1 = -38;
				 l_2 = +64; end
		6557: begin l_1 = -38;
				 l_2 = -64; end
		18081: begin l_1 = +38;
				 l_2 = +65; end
		21251: begin l_1 = +38;
				 l_2 = -65; end
		29610: begin l_1 = -38;
				 l_2 = +65; end
		32780: begin l_1 = -38;
				 l_2 = -65; end
		16496: begin l_1 = +38;
				 l_2 = +66; end
		22836: begin l_1 = +38;
				 l_2 = -66; end
		28025: begin l_1 = -38;
				 l_2 = +66; end
		34365: begin l_1 = -38;
				 l_2 = -66; end
		13326: begin l_1 = +38;
				 l_2 = +67; end
		26006: begin l_1 = +38;
				 l_2 = -67; end
		24855: begin l_1 = -38;
				 l_2 = +67; end
		37535: begin l_1 = -38;
				 l_2 = -67; end
		6986: begin l_1 = +38;
				 l_2 = +68; end
		32346: begin l_1 = +38;
				 l_2 = -68; end
		18515: begin l_1 = -38;
				 l_2 = +68; end
		43875: begin l_1 = -38;
				 l_2 = -68; end
		16274: begin l_1 = -39;
				 l_2 = +41; end
		34587: begin l_1 = -39;
				 l_2 = -40; end
		44077: begin l_1 = +39;
				 l_2 = +41; end
		6784: begin l_1 = -39;
				 l_2 = -41; end
		48822: begin l_1 = +39;
				 l_2 = +42; end
		29842: begin l_1 = +39;
				 l_2 = -42; end
		21019: begin l_1 = -39;
				 l_2 = +42; end
		2039: begin l_1 = -39;
				 l_2 = -42; end
		7451: begin l_1 = +39;
				 l_2 = +43; end
		20352: begin l_1 = +39;
				 l_2 = -43; end
		30509: begin l_1 = -39;
				 l_2 = +43; end
		43410: begin l_1 = -39;
				 l_2 = -43; end
		26431: begin l_1 = +39;
				 l_2 = +44; end
		1372: begin l_1 = +39;
				 l_2 = -44; end
		49489: begin l_1 = -39;
				 l_2 = +44; end
		24430: begin l_1 = -39;
				 l_2 = -44; end
		13530: begin l_1 = +39;
				 l_2 = +45; end
		14273: begin l_1 = +39;
				 l_2 = -45; end
		36588: begin l_1 = -39;
				 l_2 = +45; end
		37331: begin l_1 = -39;
				 l_2 = -45; end
		38589: begin l_1 = +39;
				 l_2 = +46; end
		40075: begin l_1 = +39;
				 l_2 = -46; end
		10786: begin l_1 = -39;
				 l_2 = +46; end
		12272: begin l_1 = -39;
				 l_2 = -46; end
		37846: begin l_1 = +39;
				 l_2 = +47; end
		40818: begin l_1 = +39;
				 l_2 = -47; end
		10043: begin l_1 = -39;
				 l_2 = +47; end
		13015: begin l_1 = -39;
				 l_2 = -47; end
		36360: begin l_1 = +39;
				 l_2 = +48; end
		42304: begin l_1 = +39;
				 l_2 = -48; end
		8557: begin l_1 = -39;
				 l_2 = +48; end
		14501: begin l_1 = -39;
				 l_2 = -48; end
		33388: begin l_1 = +39;
				 l_2 = +49; end
		45276: begin l_1 = +39;
				 l_2 = -49; end
		5585: begin l_1 = -39;
				 l_2 = +49; end
		17473: begin l_1 = -39;
				 l_2 = -49; end
		27444: begin l_1 = +39;
				 l_2 = +50; end
		359: begin l_1 = +39;
				 l_2 = -50; end
		50502: begin l_1 = -39;
				 l_2 = +50; end
		23417: begin l_1 = -39;
				 l_2 = -50; end
		15556: begin l_1 = +39;
				 l_2 = +51; end
		12247: begin l_1 = +39;
				 l_2 = -51; end
		38614: begin l_1 = -39;
				 l_2 = +51; end
		35305: begin l_1 = -39;
				 l_2 = -51; end
		42641: begin l_1 = +39;
				 l_2 = +52; end
		36023: begin l_1 = +39;
				 l_2 = -52; end
		14838: begin l_1 = -39;
				 l_2 = +52; end
		8220: begin l_1 = -39;
				 l_2 = -52; end
		45950: begin l_1 = +39;
				 l_2 = +53; end
		32714: begin l_1 = +39;
				 l_2 = -53; end
		18147: begin l_1 = -39;
				 l_2 = +53; end
		4911: begin l_1 = -39;
				 l_2 = -53; end
		1707: begin l_1 = +39;
				 l_2 = +54; end
		26096: begin l_1 = +39;
				 l_2 = -54; end
		24765: begin l_1 = -39;
				 l_2 = +54; end
		49154: begin l_1 = -39;
				 l_2 = -54; end
		14943: begin l_1 = +39;
				 l_2 = +55; end
		12860: begin l_1 = +39;
				 l_2 = -55; end
		38001: begin l_1 = -39;
				 l_2 = +55; end
		35918: begin l_1 = -39;
				 l_2 = -55; end
		41415: begin l_1 = +39;
				 l_2 = +56; end
		37249: begin l_1 = +39;
				 l_2 = -56; end
		13612: begin l_1 = -39;
				 l_2 = +56; end
		9446: begin l_1 = -39;
				 l_2 = -56; end
		43498: begin l_1 = +39;
				 l_2 = +57; end
		35166: begin l_1 = +39;
				 l_2 = -57; end
		15695: begin l_1 = -39;
				 l_2 = +57; end
		7363: begin l_1 = -39;
				 l_2 = -57; end
		47664: begin l_1 = +39;
				 l_2 = +58; end
		31000: begin l_1 = +39;
				 l_2 = -58; end
		19861: begin l_1 = -39;
				 l_2 = +58; end
		3197: begin l_1 = -39;
				 l_2 = -58; end
		5135: begin l_1 = +39;
				 l_2 = +59; end
		22668: begin l_1 = +39;
				 l_2 = -59; end
		28193: begin l_1 = -39;
				 l_2 = +59; end
		45726: begin l_1 = -39;
				 l_2 = -59; end
		21799: begin l_1 = +39;
				 l_2 = +60; end
		6004: begin l_1 = +39;
				 l_2 = -60; end
		44857: begin l_1 = -39;
				 l_2 = +60; end
		29062: begin l_1 = -39;
				 l_2 = -60; end
		4266: begin l_1 = +39;
				 l_2 = +61; end
		23537: begin l_1 = +39;
				 l_2 = -61; end
		27324: begin l_1 = -39;
				 l_2 = +61; end
		46595: begin l_1 = -39;
				 l_2 = -61; end
		20061: begin l_1 = +39;
				 l_2 = +62; end
		7742: begin l_1 = +39;
				 l_2 = -62; end
		43119: begin l_1 = -39;
				 l_2 = +62; end
		30800: begin l_1 = -39;
				 l_2 = -62; end
		790: begin l_1 = +39;
				 l_2 = +63; end
		27013: begin l_1 = +39;
				 l_2 = -63; end
		23848: begin l_1 = -39;
				 l_2 = +63; end
		50071: begin l_1 = -39;
				 l_2 = -63; end
		13109: begin l_1 = +39;
				 l_2 = +64; end
		14694: begin l_1 = +39;
				 l_2 = -64; end
		36167: begin l_1 = -39;
				 l_2 = +64; end
		37752: begin l_1 = -39;
				 l_2 = -64; end
		37747: begin l_1 = +39;
				 l_2 = +65; end
		40917: begin l_1 = +39;
				 l_2 = -65; end
		9944: begin l_1 = -39;
				 l_2 = +65; end
		13114: begin l_1 = -39;
				 l_2 = -65; end
		36162: begin l_1 = +39;
				 l_2 = +66; end
		42502: begin l_1 = +39;
				 l_2 = -66; end
		8359: begin l_1 = -39;
				 l_2 = +66; end
		14699: begin l_1 = -39;
				 l_2 = -66; end
		32992: begin l_1 = +39;
				 l_2 = +67; end
		45672: begin l_1 = +39;
				 l_2 = -67; end
		5189: begin l_1 = -39;
				 l_2 = +67; end
		17869: begin l_1 = -39;
				 l_2 = -67; end
		26652: begin l_1 = +39;
				 l_2 = +68; end
		1151: begin l_1 = +39;
				 l_2 = -68; end
		49710: begin l_1 = -39;
				 l_2 = +68; end
		24209: begin l_1 = -39;
				 l_2 = -68; end
		32548: begin l_1 = -40;
				 l_2 = +42; end
		18313: begin l_1 = -40;
				 l_2 = -41; end
		37293: begin l_1 = +40;
				 l_2 = +42; end
		13568: begin l_1 = -40;
				 l_2 = -42; end
		46783: begin l_1 = +40;
				 l_2 = +43; end
		8823: begin l_1 = +40;
				 l_2 = -43; end
		42038: begin l_1 = -40;
				 l_2 = +43; end
		4078: begin l_1 = -40;
				 l_2 = -43; end
		14902: begin l_1 = +40;
				 l_2 = +44; end
		40704: begin l_1 = +40;
				 l_2 = -44; end
		10157: begin l_1 = -40;
				 l_2 = +44; end
		35959: begin l_1 = -40;
				 l_2 = -44; end
		2001: begin l_1 = +40;
				 l_2 = +45; end
		2744: begin l_1 = +40;
				 l_2 = -45; end
		48117: begin l_1 = -40;
				 l_2 = +45; end
		48860: begin l_1 = -40;
				 l_2 = -45; end
		27060: begin l_1 = +40;
				 l_2 = +46; end
		28546: begin l_1 = +40;
				 l_2 = -46; end
		22315: begin l_1 = -40;
				 l_2 = +46; end
		23801: begin l_1 = -40;
				 l_2 = -46; end
		26317: begin l_1 = +40;
				 l_2 = +47; end
		29289: begin l_1 = +40;
				 l_2 = -47; end
		21572: begin l_1 = -40;
				 l_2 = +47; end
		24544: begin l_1 = -40;
				 l_2 = -47; end
		24831: begin l_1 = +40;
				 l_2 = +48; end
		30775: begin l_1 = +40;
				 l_2 = -48; end
		20086: begin l_1 = -40;
				 l_2 = +48; end
		26030: begin l_1 = -40;
				 l_2 = -48; end
		21859: begin l_1 = +40;
				 l_2 = +49; end
		33747: begin l_1 = +40;
				 l_2 = -49; end
		17114: begin l_1 = -40;
				 l_2 = +49; end
		29002: begin l_1 = -40;
				 l_2 = -49; end
		15915: begin l_1 = +40;
				 l_2 = +50; end
		39691: begin l_1 = +40;
				 l_2 = -50; end
		11170: begin l_1 = -40;
				 l_2 = +50; end
		34946: begin l_1 = -40;
				 l_2 = -50; end
		4027: begin l_1 = +40;
				 l_2 = +51; end
		718: begin l_1 = +40;
				 l_2 = -51; end
		50143: begin l_1 = -40;
				 l_2 = +51; end
		46834: begin l_1 = -40;
				 l_2 = -51; end
		31112: begin l_1 = +40;
				 l_2 = +52; end
		24494: begin l_1 = +40;
				 l_2 = -52; end
		26367: begin l_1 = -40;
				 l_2 = +52; end
		19749: begin l_1 = -40;
				 l_2 = -52; end
		34421: begin l_1 = +40;
				 l_2 = +53; end
		21185: begin l_1 = +40;
				 l_2 = -53; end
		29676: begin l_1 = -40;
				 l_2 = +53; end
		16440: begin l_1 = -40;
				 l_2 = -53; end
		41039: begin l_1 = +40;
				 l_2 = +54; end
		14567: begin l_1 = +40;
				 l_2 = -54; end
		36294: begin l_1 = -40;
				 l_2 = +54; end
		9822: begin l_1 = -40;
				 l_2 = -54; end
		3414: begin l_1 = +40;
				 l_2 = +55; end
		1331: begin l_1 = +40;
				 l_2 = -55; end
		49530: begin l_1 = -40;
				 l_2 = +55; end
		47447: begin l_1 = -40;
				 l_2 = -55; end
		29886: begin l_1 = +40;
				 l_2 = +56; end
		25720: begin l_1 = +40;
				 l_2 = -56; end
		25141: begin l_1 = -40;
				 l_2 = +56; end
		20975: begin l_1 = -40;
				 l_2 = -56; end
		31969: begin l_1 = +40;
				 l_2 = +57; end
		23637: begin l_1 = +40;
				 l_2 = -57; end
		27224: begin l_1 = -40;
				 l_2 = +57; end
		18892: begin l_1 = -40;
				 l_2 = -57; end
		36135: begin l_1 = +40;
				 l_2 = +58; end
		19471: begin l_1 = +40;
				 l_2 = -58; end
		31390: begin l_1 = -40;
				 l_2 = +58; end
		14726: begin l_1 = -40;
				 l_2 = -58; end
		44467: begin l_1 = +40;
				 l_2 = +59; end
		11139: begin l_1 = +40;
				 l_2 = -59; end
		39722: begin l_1 = -40;
				 l_2 = +59; end
		6394: begin l_1 = -40;
				 l_2 = -59; end
		10270: begin l_1 = +40;
				 l_2 = +60; end
		45336: begin l_1 = +40;
				 l_2 = -60; end
		5525: begin l_1 = -40;
				 l_2 = +60; end
		40591: begin l_1 = -40;
				 l_2 = -60; end
		43598: begin l_1 = +40;
				 l_2 = +61; end
		12008: begin l_1 = +40;
				 l_2 = -61; end
		38853: begin l_1 = -40;
				 l_2 = +61; end
		7263: begin l_1 = -40;
				 l_2 = -61; end
		8532: begin l_1 = +40;
				 l_2 = +62; end
		47074: begin l_1 = +40;
				 l_2 = -62; end
		3787: begin l_1 = -40;
				 l_2 = +62; end
		42329: begin l_1 = -40;
				 l_2 = -62; end
		40122: begin l_1 = +40;
				 l_2 = +63; end
		15484: begin l_1 = +40;
				 l_2 = -63; end
		35377: begin l_1 = -40;
				 l_2 = +63; end
		10739: begin l_1 = -40;
				 l_2 = -63; end
		1580: begin l_1 = +40;
				 l_2 = +64; end
		3165: begin l_1 = +40;
				 l_2 = -64; end
		47696: begin l_1 = -40;
				 l_2 = +64; end
		49281: begin l_1 = -40;
				 l_2 = -64; end
		26218: begin l_1 = +40;
				 l_2 = +65; end
		29388: begin l_1 = +40;
				 l_2 = -65; end
		21473: begin l_1 = -40;
				 l_2 = +65; end
		24643: begin l_1 = -40;
				 l_2 = -65; end
		24633: begin l_1 = +40;
				 l_2 = +66; end
		30973: begin l_1 = +40;
				 l_2 = -66; end
		19888: begin l_1 = -40;
				 l_2 = +66; end
		26228: begin l_1 = -40;
				 l_2 = -66; end
		21463: begin l_1 = +40;
				 l_2 = +67; end
		34143: begin l_1 = +40;
				 l_2 = -67; end
		16718: begin l_1 = -40;
				 l_2 = +67; end
		29398: begin l_1 = -40;
				 l_2 = -67; end
		15123: begin l_1 = +40;
				 l_2 = +68; end
		40483: begin l_1 = +40;
				 l_2 = -68; end
		10378: begin l_1 = -40;
				 l_2 = +68; end
		35738: begin l_1 = -40;
				 l_2 = -68; end
		14235: begin l_1 = -41;
				 l_2 = +43; end
		36626: begin l_1 = -41;
				 l_2 = -42; end
		23725: begin l_1 = +41;
				 l_2 = +43; end
		27136: begin l_1 = -41;
				 l_2 = -43; end
		42705: begin l_1 = +41;
				 l_2 = +44; end
		17646: begin l_1 = +41;
				 l_2 = -44; end
		33215: begin l_1 = -41;
				 l_2 = +44; end
		8156: begin l_1 = -41;
				 l_2 = -44; end
		29804: begin l_1 = +41;
				 l_2 = +45; end
		30547: begin l_1 = +41;
				 l_2 = -45; end
		20314: begin l_1 = -41;
				 l_2 = +45; end
		21057: begin l_1 = -41;
				 l_2 = -45; end
		4002: begin l_1 = +41;
				 l_2 = +46; end
		5488: begin l_1 = +41;
				 l_2 = -46; end
		45373: begin l_1 = -41;
				 l_2 = +46; end
		46859: begin l_1 = -41;
				 l_2 = -46; end
		3259: begin l_1 = +41;
				 l_2 = +47; end
		6231: begin l_1 = +41;
				 l_2 = -47; end
		44630: begin l_1 = -41;
				 l_2 = +47; end
		47602: begin l_1 = -41;
				 l_2 = -47; end
		1773: begin l_1 = +41;
				 l_2 = +48; end
		7717: begin l_1 = +41;
				 l_2 = -48; end
		43144: begin l_1 = -41;
				 l_2 = +48; end
		49088: begin l_1 = -41;
				 l_2 = -48; end
		49662: begin l_1 = +41;
				 l_2 = +49; end
		10689: begin l_1 = +41;
				 l_2 = -49; end
		40172: begin l_1 = -41;
				 l_2 = +49; end
		1199: begin l_1 = -41;
				 l_2 = -49; end
		43718: begin l_1 = +41;
				 l_2 = +50; end
		16633: begin l_1 = +41;
				 l_2 = -50; end
		34228: begin l_1 = -41;
				 l_2 = +50; end
		7143: begin l_1 = -41;
				 l_2 = -50; end
		31830: begin l_1 = +41;
				 l_2 = +51; end
		28521: begin l_1 = +41;
				 l_2 = -51; end
		22340: begin l_1 = -41;
				 l_2 = +51; end
		19031: begin l_1 = -41;
				 l_2 = -51; end
		8054: begin l_1 = +41;
				 l_2 = +52; end
		1436: begin l_1 = +41;
				 l_2 = -52; end
		49425: begin l_1 = -41;
				 l_2 = +52; end
		42807: begin l_1 = -41;
				 l_2 = -52; end
		11363: begin l_1 = +41;
				 l_2 = +53; end
		48988: begin l_1 = +41;
				 l_2 = -53; end
		1873: begin l_1 = -41;
				 l_2 = +53; end
		39498: begin l_1 = -41;
				 l_2 = -53; end
		17981: begin l_1 = +41;
				 l_2 = +54; end
		42370: begin l_1 = +41;
				 l_2 = -54; end
		8491: begin l_1 = -41;
				 l_2 = +54; end
		32880: begin l_1 = -41;
				 l_2 = -54; end
		31217: begin l_1 = +41;
				 l_2 = +55; end
		29134: begin l_1 = +41;
				 l_2 = -55; end
		21727: begin l_1 = -41;
				 l_2 = +55; end
		19644: begin l_1 = -41;
				 l_2 = -55; end
		6828: begin l_1 = +41;
				 l_2 = +56; end
		2662: begin l_1 = +41;
				 l_2 = -56; end
		48199: begin l_1 = -41;
				 l_2 = +56; end
		44033: begin l_1 = -41;
				 l_2 = -56; end
		8911: begin l_1 = +41;
				 l_2 = +57; end
		579: begin l_1 = +41;
				 l_2 = -57; end
		50282: begin l_1 = -41;
				 l_2 = +57; end
		41950: begin l_1 = -41;
				 l_2 = -57; end
		13077: begin l_1 = +41;
				 l_2 = +58; end
		47274: begin l_1 = +41;
				 l_2 = -58; end
		3587: begin l_1 = -41;
				 l_2 = +58; end
		37784: begin l_1 = -41;
				 l_2 = -58; end
		21409: begin l_1 = +41;
				 l_2 = +59; end
		38942: begin l_1 = +41;
				 l_2 = -59; end
		11919: begin l_1 = -41;
				 l_2 = +59; end
		29452: begin l_1 = -41;
				 l_2 = -59; end
		38073: begin l_1 = +41;
				 l_2 = +60; end
		22278: begin l_1 = +41;
				 l_2 = -60; end
		28583: begin l_1 = -41;
				 l_2 = +60; end
		12788: begin l_1 = -41;
				 l_2 = -60; end
		20540: begin l_1 = +41;
				 l_2 = +61; end
		39811: begin l_1 = +41;
				 l_2 = -61; end
		11050: begin l_1 = -41;
				 l_2 = +61; end
		30321: begin l_1 = -41;
				 l_2 = -61; end
		36335: begin l_1 = +41;
				 l_2 = +62; end
		24016: begin l_1 = +41;
				 l_2 = -62; end
		26845: begin l_1 = -41;
				 l_2 = +62; end
		14526: begin l_1 = -41;
				 l_2 = -62; end
		17064: begin l_1 = +41;
				 l_2 = +63; end
		43287: begin l_1 = +41;
				 l_2 = -63; end
		7574: begin l_1 = -41;
				 l_2 = +63; end
		33797: begin l_1 = -41;
				 l_2 = -63; end
		29383: begin l_1 = +41;
				 l_2 = +64; end
		30968: begin l_1 = +41;
				 l_2 = -64; end
		19893: begin l_1 = -41;
				 l_2 = +64; end
		21478: begin l_1 = -41;
				 l_2 = -64; end
		3160: begin l_1 = +41;
				 l_2 = +65; end
		6330: begin l_1 = +41;
				 l_2 = -65; end
		44531: begin l_1 = -41;
				 l_2 = +65; end
		47701: begin l_1 = -41;
				 l_2 = -65; end
		1575: begin l_1 = +41;
				 l_2 = +66; end
		7915: begin l_1 = +41;
				 l_2 = -66; end
		42946: begin l_1 = -41;
				 l_2 = +66; end
		49286: begin l_1 = -41;
				 l_2 = -66; end
		49266: begin l_1 = +41;
				 l_2 = +67; end
		11085: begin l_1 = +41;
				 l_2 = -67; end
		39776: begin l_1 = -41;
				 l_2 = +67; end
		1595: begin l_1 = -41;
				 l_2 = -67; end
		42926: begin l_1 = +41;
				 l_2 = +68; end
		17425: begin l_1 = +41;
				 l_2 = -68; end
		33436: begin l_1 = -41;
				 l_2 = +68; end
		7935: begin l_1 = -41;
				 l_2 = -68; end
		28470: begin l_1 = -42;
				 l_2 = +44; end
		22391: begin l_1 = -42;
				 l_2 = -43; end
		47450: begin l_1 = +42;
				 l_2 = +44; end
		3411: begin l_1 = -42;
				 l_2 = -44; end
		34549: begin l_1 = +42;
				 l_2 = +45; end
		35292: begin l_1 = +42;
				 l_2 = -45; end
		15569: begin l_1 = -42;
				 l_2 = +45; end
		16312: begin l_1 = -42;
				 l_2 = -45; end
		8747: begin l_1 = +42;
				 l_2 = +46; end
		10233: begin l_1 = +42;
				 l_2 = -46; end
		40628: begin l_1 = -42;
				 l_2 = +46; end
		42114: begin l_1 = -42;
				 l_2 = -46; end
		8004: begin l_1 = +42;
				 l_2 = +47; end
		10976: begin l_1 = +42;
				 l_2 = -47; end
		39885: begin l_1 = -42;
				 l_2 = +47; end
		42857: begin l_1 = -42;
				 l_2 = -47; end
		6518: begin l_1 = +42;
				 l_2 = +48; end
		12462: begin l_1 = +42;
				 l_2 = -48; end
		38399: begin l_1 = -42;
				 l_2 = +48; end
		44343: begin l_1 = -42;
				 l_2 = -48; end
		3546: begin l_1 = +42;
				 l_2 = +49; end
		15434: begin l_1 = +42;
				 l_2 = -49; end
		35427: begin l_1 = -42;
				 l_2 = +49; end
		47315: begin l_1 = -42;
				 l_2 = -49; end
		48463: begin l_1 = +42;
				 l_2 = +50; end
		21378: begin l_1 = +42;
				 l_2 = -50; end
		29483: begin l_1 = -42;
				 l_2 = +50; end
		2398: begin l_1 = -42;
				 l_2 = -50; end
		36575: begin l_1 = +42;
				 l_2 = +51; end
		33266: begin l_1 = +42;
				 l_2 = -51; end
		17595: begin l_1 = -42;
				 l_2 = +51; end
		14286: begin l_1 = -42;
				 l_2 = -51; end
		12799: begin l_1 = +42;
				 l_2 = +52; end
		6181: begin l_1 = +42;
				 l_2 = -52; end
		44680: begin l_1 = -42;
				 l_2 = +52; end
		38062: begin l_1 = -42;
				 l_2 = -52; end
		16108: begin l_1 = +42;
				 l_2 = +53; end
		2872: begin l_1 = +42;
				 l_2 = -53; end
		47989: begin l_1 = -42;
				 l_2 = +53; end
		34753: begin l_1 = -42;
				 l_2 = -53; end
		22726: begin l_1 = +42;
				 l_2 = +54; end
		47115: begin l_1 = +42;
				 l_2 = -54; end
		3746: begin l_1 = -42;
				 l_2 = +54; end
		28135: begin l_1 = -42;
				 l_2 = -54; end
		35962: begin l_1 = +42;
				 l_2 = +55; end
		33879: begin l_1 = +42;
				 l_2 = -55; end
		16982: begin l_1 = -42;
				 l_2 = +55; end
		14899: begin l_1 = -42;
				 l_2 = -55; end
		11573: begin l_1 = +42;
				 l_2 = +56; end
		7407: begin l_1 = +42;
				 l_2 = -56; end
		43454: begin l_1 = -42;
				 l_2 = +56; end
		39288: begin l_1 = -42;
				 l_2 = -56; end
		13656: begin l_1 = +42;
				 l_2 = +57; end
		5324: begin l_1 = +42;
				 l_2 = -57; end
		45537: begin l_1 = -42;
				 l_2 = +57; end
		37205: begin l_1 = -42;
				 l_2 = -57; end
		17822: begin l_1 = +42;
				 l_2 = +58; end
		1158: begin l_1 = +42;
				 l_2 = -58; end
		49703: begin l_1 = -42;
				 l_2 = +58; end
		33039: begin l_1 = -42;
				 l_2 = -58; end
		26154: begin l_1 = +42;
				 l_2 = +59; end
		43687: begin l_1 = +42;
				 l_2 = -59; end
		7174: begin l_1 = -42;
				 l_2 = +59; end
		24707: begin l_1 = -42;
				 l_2 = -59; end
		42818: begin l_1 = +42;
				 l_2 = +60; end
		27023: begin l_1 = +42;
				 l_2 = -60; end
		23838: begin l_1 = -42;
				 l_2 = +60; end
		8043: begin l_1 = -42;
				 l_2 = -60; end
		25285: begin l_1 = +42;
				 l_2 = +61; end
		44556: begin l_1 = +42;
				 l_2 = -61; end
		6305: begin l_1 = -42;
				 l_2 = +61; end
		25576: begin l_1 = -42;
				 l_2 = -61; end
		41080: begin l_1 = +42;
				 l_2 = +62; end
		28761: begin l_1 = +42;
				 l_2 = -62; end
		22100: begin l_1 = -42;
				 l_2 = +62; end
		9781: begin l_1 = -42;
				 l_2 = -62; end
		21809: begin l_1 = +42;
				 l_2 = +63; end
		48032: begin l_1 = +42;
				 l_2 = -63; end
		2829: begin l_1 = -42;
				 l_2 = +63; end
		29052: begin l_1 = -42;
				 l_2 = -63; end
		34128: begin l_1 = +42;
				 l_2 = +64; end
		35713: begin l_1 = +42;
				 l_2 = -64; end
		15148: begin l_1 = -42;
				 l_2 = +64; end
		16733: begin l_1 = -42;
				 l_2 = -64; end
		7905: begin l_1 = +42;
				 l_2 = +65; end
		11075: begin l_1 = +42;
				 l_2 = -65; end
		39786: begin l_1 = -42;
				 l_2 = +65; end
		42956: begin l_1 = -42;
				 l_2 = -65; end
		6320: begin l_1 = +42;
				 l_2 = +66; end
		12660: begin l_1 = +42;
				 l_2 = -66; end
		38201: begin l_1 = -42;
				 l_2 = +66; end
		44541: begin l_1 = -42;
				 l_2 = -66; end
		3150: begin l_1 = +42;
				 l_2 = +67; end
		15830: begin l_1 = +42;
				 l_2 = -67; end
		35031: begin l_1 = -42;
				 l_2 = +67; end
		47711: begin l_1 = -42;
				 l_2 = -67; end
		47671: begin l_1 = +42;
				 l_2 = +68; end
		22170: begin l_1 = +42;
				 l_2 = -68; end
		28691: begin l_1 = -42;
				 l_2 = +68; end
		3190: begin l_1 = -42;
				 l_2 = -68; end
		6079: begin l_1 = -43;
				 l_2 = +45; end
		44782: begin l_1 = -43;
				 l_2 = -44; end
		44039: begin l_1 = +43;
				 l_2 = +45; end
		6822: begin l_1 = -43;
				 l_2 = -45; end
		18237: begin l_1 = +43;
				 l_2 = +46; end
		19723: begin l_1 = +43;
				 l_2 = -46; end
		31138: begin l_1 = -43;
				 l_2 = +46; end
		32624: begin l_1 = -43;
				 l_2 = -46; end
		17494: begin l_1 = +43;
				 l_2 = +47; end
		20466: begin l_1 = +43;
				 l_2 = -47; end
		30395: begin l_1 = -43;
				 l_2 = +47; end
		33367: begin l_1 = -43;
				 l_2 = -47; end
		16008: begin l_1 = +43;
				 l_2 = +48; end
		21952: begin l_1 = +43;
				 l_2 = -48; end
		28909: begin l_1 = -43;
				 l_2 = +48; end
		34853: begin l_1 = -43;
				 l_2 = -48; end
		13036: begin l_1 = +43;
				 l_2 = +49; end
		24924: begin l_1 = +43;
				 l_2 = -49; end
		25937: begin l_1 = -43;
				 l_2 = +49; end
		37825: begin l_1 = -43;
				 l_2 = -49; end
		7092: begin l_1 = +43;
				 l_2 = +50; end
		30868: begin l_1 = +43;
				 l_2 = -50; end
		19993: begin l_1 = -43;
				 l_2 = +50; end
		43769: begin l_1 = -43;
				 l_2 = -50; end
		46065: begin l_1 = +43;
				 l_2 = +51; end
		42756: begin l_1 = +43;
				 l_2 = -51; end
		8105: begin l_1 = -43;
				 l_2 = +51; end
		4796: begin l_1 = -43;
				 l_2 = -51; end
		22289: begin l_1 = +43;
				 l_2 = +52; end
		15671: begin l_1 = +43;
				 l_2 = -52; end
		35190: begin l_1 = -43;
				 l_2 = +52; end
		28572: begin l_1 = -43;
				 l_2 = -52; end
		25598: begin l_1 = +43;
				 l_2 = +53; end
		12362: begin l_1 = +43;
				 l_2 = -53; end
		38499: begin l_1 = -43;
				 l_2 = +53; end
		25263: begin l_1 = -43;
				 l_2 = -53; end
		32216: begin l_1 = +43;
				 l_2 = +54; end
		5744: begin l_1 = +43;
				 l_2 = -54; end
		45117: begin l_1 = -43;
				 l_2 = +54; end
		18645: begin l_1 = -43;
				 l_2 = -54; end
		45452: begin l_1 = +43;
				 l_2 = +55; end
		43369: begin l_1 = +43;
				 l_2 = -55; end
		7492: begin l_1 = -43;
				 l_2 = +55; end
		5409: begin l_1 = -43;
				 l_2 = -55; end
		21063: begin l_1 = +43;
				 l_2 = +56; end
		16897: begin l_1 = +43;
				 l_2 = -56; end
		33964: begin l_1 = -43;
				 l_2 = +56; end
		29798: begin l_1 = -43;
				 l_2 = -56; end
		23146: begin l_1 = +43;
				 l_2 = +57; end
		14814: begin l_1 = +43;
				 l_2 = -57; end
		36047: begin l_1 = -43;
				 l_2 = +57; end
		27715: begin l_1 = -43;
				 l_2 = -57; end
		27312: begin l_1 = +43;
				 l_2 = +58; end
		10648: begin l_1 = +43;
				 l_2 = -58; end
		40213: begin l_1 = -43;
				 l_2 = +58; end
		23549: begin l_1 = -43;
				 l_2 = -58; end
		35644: begin l_1 = +43;
				 l_2 = +59; end
		2316: begin l_1 = +43;
				 l_2 = -59; end
		48545: begin l_1 = -43;
				 l_2 = +59; end
		15217: begin l_1 = -43;
				 l_2 = -59; end
		1447: begin l_1 = +43;
				 l_2 = +60; end
		36513: begin l_1 = +43;
				 l_2 = -60; end
		14348: begin l_1 = -43;
				 l_2 = +60; end
		49414: begin l_1 = -43;
				 l_2 = -60; end
		34775: begin l_1 = +43;
				 l_2 = +61; end
		3185: begin l_1 = +43;
				 l_2 = -61; end
		47676: begin l_1 = -43;
				 l_2 = +61; end
		16086: begin l_1 = -43;
				 l_2 = -61; end
		50570: begin l_1 = +43;
				 l_2 = +62; end
		38251: begin l_1 = +43;
				 l_2 = -62; end
		12610: begin l_1 = -43;
				 l_2 = +62; end
		291: begin l_1 = -43;
				 l_2 = -62; end
		31299: begin l_1 = +43;
				 l_2 = +63; end
		6661: begin l_1 = +43;
				 l_2 = -63; end
		44200: begin l_1 = -43;
				 l_2 = +63; end
		19562: begin l_1 = -43;
				 l_2 = -63; end
		43618: begin l_1 = +43;
				 l_2 = +64; end
		45203: begin l_1 = +43;
				 l_2 = -64; end
		5658: begin l_1 = -43;
				 l_2 = +64; end
		7243: begin l_1 = -43;
				 l_2 = -64; end
		17395: begin l_1 = +43;
				 l_2 = +65; end
		20565: begin l_1 = +43;
				 l_2 = -65; end
		30296: begin l_1 = -43;
				 l_2 = +65; end
		33466: begin l_1 = -43;
				 l_2 = -65; end
		15810: begin l_1 = +43;
				 l_2 = +66; end
		22150: begin l_1 = +43;
				 l_2 = -66; end
		28711: begin l_1 = -43;
				 l_2 = +66; end
		35051: begin l_1 = -43;
				 l_2 = -66; end
		12640: begin l_1 = +43;
				 l_2 = +67; end
		25320: begin l_1 = +43;
				 l_2 = -67; end
		25541: begin l_1 = -43;
				 l_2 = +67; end
		38221: begin l_1 = -43;
				 l_2 = -67; end
		6300: begin l_1 = +43;
				 l_2 = +68; end
		31660: begin l_1 = +43;
				 l_2 = -68; end
		19201: begin l_1 = -43;
				 l_2 = +68; end
		44561: begin l_1 = -43;
				 l_2 = -68; end
		12158: begin l_1 = -44;
				 l_2 = +46; end
		38703: begin l_1 = -44;
				 l_2 = -45; end
		37217: begin l_1 = +44;
				 l_2 = +46; end
		13644: begin l_1 = -44;
				 l_2 = -46; end
		36474: begin l_1 = +44;
				 l_2 = +47; end
		39446: begin l_1 = +44;
				 l_2 = -47; end
		11415: begin l_1 = -44;
				 l_2 = +47; end
		14387: begin l_1 = -44;
				 l_2 = -47; end
		34988: begin l_1 = +44;
				 l_2 = +48; end
		40932: begin l_1 = +44;
				 l_2 = -48; end
		9929: begin l_1 = -44;
				 l_2 = +48; end
		15873: begin l_1 = -44;
				 l_2 = -48; end
		32016: begin l_1 = +44;
				 l_2 = +49; end
		43904: begin l_1 = +44;
				 l_2 = -49; end
		6957: begin l_1 = -44;
				 l_2 = +49; end
		18845: begin l_1 = -44;
				 l_2 = -49; end
		26072: begin l_1 = +44;
				 l_2 = +50; end
		49848: begin l_1 = +44;
				 l_2 = -50; end
		1013: begin l_1 = -44;
				 l_2 = +50; end
		24789: begin l_1 = -44;
				 l_2 = -50; end
		14184: begin l_1 = +44;
				 l_2 = +51; end
		10875: begin l_1 = +44;
				 l_2 = -51; end
		39986: begin l_1 = -44;
				 l_2 = +51; end
		36677: begin l_1 = -44;
				 l_2 = -51; end
		41269: begin l_1 = +44;
				 l_2 = +52; end
		34651: begin l_1 = +44;
				 l_2 = -52; end
		16210: begin l_1 = -44;
				 l_2 = +52; end
		9592: begin l_1 = -44;
				 l_2 = -52; end
		44578: begin l_1 = +44;
				 l_2 = +53; end
		31342: begin l_1 = +44;
				 l_2 = -53; end
		19519: begin l_1 = -44;
				 l_2 = +53; end
		6283: begin l_1 = -44;
				 l_2 = -53; end
		335: begin l_1 = +44;
				 l_2 = +54; end
		24724: begin l_1 = +44;
				 l_2 = -54; end
		26137: begin l_1 = -44;
				 l_2 = +54; end
		50526: begin l_1 = -44;
				 l_2 = -54; end
		13571: begin l_1 = +44;
				 l_2 = +55; end
		11488: begin l_1 = +44;
				 l_2 = -55; end
		39373: begin l_1 = -44;
				 l_2 = +55; end
		37290: begin l_1 = -44;
				 l_2 = -55; end
		40043: begin l_1 = +44;
				 l_2 = +56; end
		35877: begin l_1 = +44;
				 l_2 = -56; end
		14984: begin l_1 = -44;
				 l_2 = +56; end
		10818: begin l_1 = -44;
				 l_2 = -56; end
		42126: begin l_1 = +44;
				 l_2 = +57; end
		33794: begin l_1 = +44;
				 l_2 = -57; end
		17067: begin l_1 = -44;
				 l_2 = +57; end
		8735: begin l_1 = -44;
				 l_2 = -57; end
		46292: begin l_1 = +44;
				 l_2 = +58; end
		29628: begin l_1 = +44;
				 l_2 = -58; end
		21233: begin l_1 = -44;
				 l_2 = +58; end
		4569: begin l_1 = -44;
				 l_2 = -58; end
		3763: begin l_1 = +44;
				 l_2 = +59; end
		21296: begin l_1 = +44;
				 l_2 = -59; end
		29565: begin l_1 = -44;
				 l_2 = +59; end
		47098: begin l_1 = -44;
				 l_2 = -59; end
		20427: begin l_1 = +44;
				 l_2 = +60; end
		4632: begin l_1 = +44;
				 l_2 = -60; end
		46229: begin l_1 = -44;
				 l_2 = +60; end
		30434: begin l_1 = -44;
				 l_2 = -60; end
		2894: begin l_1 = +44;
				 l_2 = +61; end
		22165: begin l_1 = +44;
				 l_2 = -61; end
		28696: begin l_1 = -44;
				 l_2 = +61; end
		47967: begin l_1 = -44;
				 l_2 = -61; end
		18689: begin l_1 = +44;
				 l_2 = +62; end
		6370: begin l_1 = +44;
				 l_2 = -62; end
		44491: begin l_1 = -44;
				 l_2 = +62; end
		32172: begin l_1 = -44;
				 l_2 = -62; end
		50279: begin l_1 = +44;
				 l_2 = +63; end
		25641: begin l_1 = +44;
				 l_2 = -63; end
		25220: begin l_1 = -44;
				 l_2 = +63; end
		582: begin l_1 = -44;
				 l_2 = -63; end
		11737: begin l_1 = +44;
				 l_2 = +64; end
		13322: begin l_1 = +44;
				 l_2 = -64; end
		37539: begin l_1 = -44;
				 l_2 = +64; end
		39124: begin l_1 = -44;
				 l_2 = -64; end
		36375: begin l_1 = +44;
				 l_2 = +65; end
		39545: begin l_1 = +44;
				 l_2 = -65; end
		11316: begin l_1 = -44;
				 l_2 = +65; end
		14486: begin l_1 = -44;
				 l_2 = -65; end
		34790: begin l_1 = +44;
				 l_2 = +66; end
		41130: begin l_1 = +44;
				 l_2 = -66; end
		9731: begin l_1 = -44;
				 l_2 = +66; end
		16071: begin l_1 = -44;
				 l_2 = -66; end
		31620: begin l_1 = +44;
				 l_2 = +67; end
		44300: begin l_1 = +44;
				 l_2 = -67; end
		6561: begin l_1 = -44;
				 l_2 = +67; end
		19241: begin l_1 = -44;
				 l_2 = -67; end
		25280: begin l_1 = +44;
				 l_2 = +68; end
		50640: begin l_1 = +44;
				 l_2 = -68; end
		221: begin l_1 = -44;
				 l_2 = +68; end
		25581: begin l_1 = -44;
				 l_2 = -68; end
		24316: begin l_1 = -45;
				 l_2 = +47; end
		26545: begin l_1 = -45;
				 l_2 = -46; end
		23573: begin l_1 = +45;
				 l_2 = +47; end
		27288: begin l_1 = -45;
				 l_2 = -47; end
		22087: begin l_1 = +45;
				 l_2 = +48; end
		28031: begin l_1 = +45;
				 l_2 = -48; end
		22830: begin l_1 = -45;
				 l_2 = +48; end
		28774: begin l_1 = -45;
				 l_2 = -48; end
		19115: begin l_1 = +45;
				 l_2 = +49; end
		31003: begin l_1 = +45;
				 l_2 = -49; end
		19858: begin l_1 = -45;
				 l_2 = +49; end
		31746: begin l_1 = -45;
				 l_2 = -49; end
		13171: begin l_1 = +45;
				 l_2 = +50; end
		36947: begin l_1 = +45;
				 l_2 = -50; end
		13914: begin l_1 = -45;
				 l_2 = +50; end
		37690: begin l_1 = -45;
				 l_2 = -50; end
		1283: begin l_1 = +45;
				 l_2 = +51; end
		48835: begin l_1 = +45;
				 l_2 = -51; end
		2026: begin l_1 = -45;
				 l_2 = +51; end
		49578: begin l_1 = -45;
				 l_2 = -51; end
		28368: begin l_1 = +45;
				 l_2 = +52; end
		21750: begin l_1 = +45;
				 l_2 = -52; end
		29111: begin l_1 = -45;
				 l_2 = +52; end
		22493: begin l_1 = -45;
				 l_2 = -52; end
		31677: begin l_1 = +45;
				 l_2 = +53; end
		18441: begin l_1 = +45;
				 l_2 = -53; end
		32420: begin l_1 = -45;
				 l_2 = +53; end
		19184: begin l_1 = -45;
				 l_2 = -53; end
		38295: begin l_1 = +45;
				 l_2 = +54; end
		11823: begin l_1 = +45;
				 l_2 = -54; end
		39038: begin l_1 = -45;
				 l_2 = +54; end
		12566: begin l_1 = -45;
				 l_2 = -54; end
		670: begin l_1 = +45;
				 l_2 = +55; end
		49448: begin l_1 = +45;
				 l_2 = -55; end
		1413: begin l_1 = -45;
				 l_2 = +55; end
		50191: begin l_1 = -45;
				 l_2 = -55; end
		27142: begin l_1 = +45;
				 l_2 = +56; end
		22976: begin l_1 = +45;
				 l_2 = -56; end
		27885: begin l_1 = -45;
				 l_2 = +56; end
		23719: begin l_1 = -45;
				 l_2 = -56; end
		29225: begin l_1 = +45;
				 l_2 = +57; end
		20893: begin l_1 = +45;
				 l_2 = -57; end
		29968: begin l_1 = -45;
				 l_2 = +57; end
		21636: begin l_1 = -45;
				 l_2 = -57; end
		33391: begin l_1 = +45;
				 l_2 = +58; end
		16727: begin l_1 = +45;
				 l_2 = -58; end
		34134: begin l_1 = -45;
				 l_2 = +58; end
		17470: begin l_1 = -45;
				 l_2 = -58; end
		41723: begin l_1 = +45;
				 l_2 = +59; end
		8395: begin l_1 = +45;
				 l_2 = -59; end
		42466: begin l_1 = -45;
				 l_2 = +59; end
		9138: begin l_1 = -45;
				 l_2 = -59; end
		7526: begin l_1 = +45;
				 l_2 = +60; end
		42592: begin l_1 = +45;
				 l_2 = -60; end
		8269: begin l_1 = -45;
				 l_2 = +60; end
		43335: begin l_1 = -45;
				 l_2 = -60; end
		40854: begin l_1 = +45;
				 l_2 = +61; end
		9264: begin l_1 = +45;
				 l_2 = -61; end
		41597: begin l_1 = -45;
				 l_2 = +61; end
		10007: begin l_1 = -45;
				 l_2 = -61; end
		5788: begin l_1 = +45;
				 l_2 = +62; end
		44330: begin l_1 = +45;
				 l_2 = -62; end
		6531: begin l_1 = -45;
				 l_2 = +62; end
		45073: begin l_1 = -45;
				 l_2 = -62; end
		37378: begin l_1 = +45;
				 l_2 = +63; end
		12740: begin l_1 = +45;
				 l_2 = -63; end
		38121: begin l_1 = -45;
				 l_2 = +63; end
		13483: begin l_1 = -45;
				 l_2 = -63; end
		49697: begin l_1 = +45;
				 l_2 = +64; end
		421: begin l_1 = +45;
				 l_2 = -64; end
		50440: begin l_1 = -45;
				 l_2 = +64; end
		1164: begin l_1 = -45;
				 l_2 = -64; end
		23474: begin l_1 = +45;
				 l_2 = +65; end
		26644: begin l_1 = +45;
				 l_2 = -65; end
		24217: begin l_1 = -45;
				 l_2 = +65; end
		27387: begin l_1 = -45;
				 l_2 = -65; end
		21889: begin l_1 = +45;
				 l_2 = +66; end
		28229: begin l_1 = +45;
				 l_2 = -66; end
		22632: begin l_1 = -45;
				 l_2 = +66; end
		28972: begin l_1 = -45;
				 l_2 = -66; end
		18719: begin l_1 = +45;
				 l_2 = +67; end
		31399: begin l_1 = +45;
				 l_2 = -67; end
		19462: begin l_1 = -45;
				 l_2 = +67; end
		32142: begin l_1 = -45;
				 l_2 = -67; end
		12379: begin l_1 = +45;
				 l_2 = +68; end
		37739: begin l_1 = +45;
				 l_2 = -68; end
		13122: begin l_1 = -45;
				 l_2 = +68; end
		38482: begin l_1 = -45;
				 l_2 = -68; end
		48632: begin l_1 = -46;
				 l_2 = +48; end
		2229: begin l_1 = -46;
				 l_2 = -47; end
		47146: begin l_1 = +46;
				 l_2 = +48; end
		3715: begin l_1 = -46;
				 l_2 = -48; end
		44174: begin l_1 = +46;
				 l_2 = +49; end
		5201: begin l_1 = +46;
				 l_2 = -49; end
		45660: begin l_1 = -46;
				 l_2 = +49; end
		6687: begin l_1 = -46;
				 l_2 = -49; end
		38230: begin l_1 = +46;
				 l_2 = +50; end
		11145: begin l_1 = +46;
				 l_2 = -50; end
		39716: begin l_1 = -46;
				 l_2 = +50; end
		12631: begin l_1 = -46;
				 l_2 = -50; end
		26342: begin l_1 = +46;
				 l_2 = +51; end
		23033: begin l_1 = +46;
				 l_2 = -51; end
		27828: begin l_1 = -46;
				 l_2 = +51; end
		24519: begin l_1 = -46;
				 l_2 = -51; end
		2566: begin l_1 = +46;
				 l_2 = +52; end
		46809: begin l_1 = +46;
				 l_2 = -52; end
		4052: begin l_1 = -46;
				 l_2 = +52; end
		48295: begin l_1 = -46;
				 l_2 = -52; end
		5875: begin l_1 = +46;
				 l_2 = +53; end
		43500: begin l_1 = +46;
				 l_2 = -53; end
		7361: begin l_1 = -46;
				 l_2 = +53; end
		44986: begin l_1 = -46;
				 l_2 = -53; end
		12493: begin l_1 = +46;
				 l_2 = +54; end
		36882: begin l_1 = +46;
				 l_2 = -54; end
		13979: begin l_1 = -46;
				 l_2 = +54; end
		38368: begin l_1 = -46;
				 l_2 = -54; end
		25729: begin l_1 = +46;
				 l_2 = +55; end
		23646: begin l_1 = +46;
				 l_2 = -55; end
		27215: begin l_1 = -46;
				 l_2 = +55; end
		25132: begin l_1 = -46;
				 l_2 = -55; end
		1340: begin l_1 = +46;
				 l_2 = +56; end
		48035: begin l_1 = +46;
				 l_2 = -56; end
		2826: begin l_1 = -46;
				 l_2 = +56; end
		49521: begin l_1 = -46;
				 l_2 = -56; end
		3423: begin l_1 = +46;
				 l_2 = +57; end
		45952: begin l_1 = +46;
				 l_2 = -57; end
		4909: begin l_1 = -46;
				 l_2 = +57; end
		47438: begin l_1 = -46;
				 l_2 = -57; end
		7589: begin l_1 = +46;
				 l_2 = +58; end
		41786: begin l_1 = +46;
				 l_2 = -58; end
		9075: begin l_1 = -46;
				 l_2 = +58; end
		43272: begin l_1 = -46;
				 l_2 = -58; end
		15921: begin l_1 = +46;
				 l_2 = +59; end
		33454: begin l_1 = +46;
				 l_2 = -59; end
		17407: begin l_1 = -46;
				 l_2 = +59; end
		34940: begin l_1 = -46;
				 l_2 = -59; end
		32585: begin l_1 = +46;
				 l_2 = +60; end
		16790: begin l_1 = +46;
				 l_2 = -60; end
		34071: begin l_1 = -46;
				 l_2 = +60; end
		18276: begin l_1 = -46;
				 l_2 = -60; end
		15052: begin l_1 = +46;
				 l_2 = +61; end
		34323: begin l_1 = +46;
				 l_2 = -61; end
		16538: begin l_1 = -46;
				 l_2 = +61; end
		35809: begin l_1 = -46;
				 l_2 = -61; end
		30847: begin l_1 = +46;
				 l_2 = +62; end
		18528: begin l_1 = +46;
				 l_2 = -62; end
		32333: begin l_1 = -46;
				 l_2 = +62; end
		20014: begin l_1 = -46;
				 l_2 = -62; end
		11576: begin l_1 = +46;
				 l_2 = +63; end
		37799: begin l_1 = +46;
				 l_2 = -63; end
		13062: begin l_1 = -46;
				 l_2 = +63; end
		39285: begin l_1 = -46;
				 l_2 = -63; end
		23895: begin l_1 = +46;
				 l_2 = +64; end
		25480: begin l_1 = +46;
				 l_2 = -64; end
		25381: begin l_1 = -46;
				 l_2 = +64; end
		26966: begin l_1 = -46;
				 l_2 = -64; end
		48533: begin l_1 = +46;
				 l_2 = +65; end
		842: begin l_1 = +46;
				 l_2 = -65; end
		50019: begin l_1 = -46;
				 l_2 = +65; end
		2328: begin l_1 = -46;
				 l_2 = -65; end
		46948: begin l_1 = +46;
				 l_2 = +66; end
		2427: begin l_1 = +46;
				 l_2 = -66; end
		48434: begin l_1 = -46;
				 l_2 = +66; end
		3913: begin l_1 = -46;
				 l_2 = -66; end
		43778: begin l_1 = +46;
				 l_2 = +67; end
		5597: begin l_1 = +46;
				 l_2 = -67; end
		45264: begin l_1 = -46;
				 l_2 = +67; end
		7083: begin l_1 = -46;
				 l_2 = -67; end
		37438: begin l_1 = +46;
				 l_2 = +68; end
		11937: begin l_1 = +46;
				 l_2 = -68; end
		38924: begin l_1 = -46;
				 l_2 = +68; end
		13423: begin l_1 = -46;
				 l_2 = -68; end
		46403: begin l_1 = -47;
				 l_2 = +49; end
		4458: begin l_1 = -47;
				 l_2 = -48; end
		43431: begin l_1 = +47;
				 l_2 = +49; end
		7430: begin l_1 = -47;
				 l_2 = -49; end
		37487: begin l_1 = +47;
				 l_2 = +50; end
		10402: begin l_1 = +47;
				 l_2 = -50; end
		40459: begin l_1 = -47;
				 l_2 = +50; end
		13374: begin l_1 = -47;
				 l_2 = -50; end
		25599: begin l_1 = +47;
				 l_2 = +51; end
		22290: begin l_1 = +47;
				 l_2 = -51; end
		28571: begin l_1 = -47;
				 l_2 = +51; end
		25262: begin l_1 = -47;
				 l_2 = -51; end
		1823: begin l_1 = +47;
				 l_2 = +52; end
		46066: begin l_1 = +47;
				 l_2 = -52; end
		4795: begin l_1 = -47;
				 l_2 = +52; end
		49038: begin l_1 = -47;
				 l_2 = -52; end
		5132: begin l_1 = +47;
				 l_2 = +53; end
		42757: begin l_1 = +47;
				 l_2 = -53; end
		8104: begin l_1 = -47;
				 l_2 = +53; end
		45729: begin l_1 = -47;
				 l_2 = -53; end
		11750: begin l_1 = +47;
				 l_2 = +54; end
		36139: begin l_1 = +47;
				 l_2 = -54; end
		14722: begin l_1 = -47;
				 l_2 = +54; end
		39111: begin l_1 = -47;
				 l_2 = -54; end
		24986: begin l_1 = +47;
				 l_2 = +55; end
		22903: begin l_1 = +47;
				 l_2 = -55; end
		27958: begin l_1 = -47;
				 l_2 = +55; end
		25875: begin l_1 = -47;
				 l_2 = -55; end
		597: begin l_1 = +47;
				 l_2 = +56; end
		47292: begin l_1 = +47;
				 l_2 = -56; end
		3569: begin l_1 = -47;
				 l_2 = +56; end
		50264: begin l_1 = -47;
				 l_2 = -56; end
		2680: begin l_1 = +47;
				 l_2 = +57; end
		45209: begin l_1 = +47;
				 l_2 = -57; end
		5652: begin l_1 = -47;
				 l_2 = +57; end
		48181: begin l_1 = -47;
				 l_2 = -57; end
		6846: begin l_1 = +47;
				 l_2 = +58; end
		41043: begin l_1 = +47;
				 l_2 = -58; end
		9818: begin l_1 = -47;
				 l_2 = +58; end
		44015: begin l_1 = -47;
				 l_2 = -58; end
		15178: begin l_1 = +47;
				 l_2 = +59; end
		32711: begin l_1 = +47;
				 l_2 = -59; end
		18150: begin l_1 = -47;
				 l_2 = +59; end
		35683: begin l_1 = -47;
				 l_2 = -59; end
		31842: begin l_1 = +47;
				 l_2 = +60; end
		16047: begin l_1 = +47;
				 l_2 = -60; end
		34814: begin l_1 = -47;
				 l_2 = +60; end
		19019: begin l_1 = -47;
				 l_2 = -60; end
		14309: begin l_1 = +47;
				 l_2 = +61; end
		33580: begin l_1 = +47;
				 l_2 = -61; end
		17281: begin l_1 = -47;
				 l_2 = +61; end
		36552: begin l_1 = -47;
				 l_2 = -61; end
		30104: begin l_1 = +47;
				 l_2 = +62; end
		17785: begin l_1 = +47;
				 l_2 = -62; end
		33076: begin l_1 = -47;
				 l_2 = +62; end
		20757: begin l_1 = -47;
				 l_2 = -62; end
		10833: begin l_1 = +47;
				 l_2 = +63; end
		37056: begin l_1 = +47;
				 l_2 = -63; end
		13805: begin l_1 = -47;
				 l_2 = +63; end
		40028: begin l_1 = -47;
				 l_2 = -63; end
		23152: begin l_1 = +47;
				 l_2 = +64; end
		24737: begin l_1 = +47;
				 l_2 = -64; end
		26124: begin l_1 = -47;
				 l_2 = +64; end
		27709: begin l_1 = -47;
				 l_2 = -64; end
		47790: begin l_1 = +47;
				 l_2 = +65; end
		99: begin l_1 = +47;
				 l_2 = -65; end
		50762: begin l_1 = -47;
				 l_2 = +65; end
		3071: begin l_1 = -47;
				 l_2 = -65; end
		46205: begin l_1 = +47;
				 l_2 = +66; end
		1684: begin l_1 = +47;
				 l_2 = -66; end
		49177: begin l_1 = -47;
				 l_2 = +66; end
		4656: begin l_1 = -47;
				 l_2 = -66; end
		43035: begin l_1 = +47;
				 l_2 = +67; end
		4854: begin l_1 = +47;
				 l_2 = -67; end
		46007: begin l_1 = -47;
				 l_2 = +67; end
		7826: begin l_1 = -47;
				 l_2 = -67; end
		36695: begin l_1 = +47;
				 l_2 = +68; end
		11194: begin l_1 = +47;
				 l_2 = -68; end
		39667: begin l_1 = -47;
				 l_2 = +68; end
		14166: begin l_1 = -47;
				 l_2 = -68; end
		41945: begin l_1 = -48;
				 l_2 = +50; end
		8916: begin l_1 = -48;
				 l_2 = -49; end
		36001: begin l_1 = +48;
				 l_2 = +50; end
		14860: begin l_1 = -48;
				 l_2 = -50; end
		24113: begin l_1 = +48;
				 l_2 = +51; end
		20804: begin l_1 = +48;
				 l_2 = -51; end
		30057: begin l_1 = -48;
				 l_2 = +51; end
		26748: begin l_1 = -48;
				 l_2 = -51; end
		337: begin l_1 = +48;
				 l_2 = +52; end
		44580: begin l_1 = +48;
				 l_2 = -52; end
		6281: begin l_1 = -48;
				 l_2 = +52; end
		50524: begin l_1 = -48;
				 l_2 = -52; end
		3646: begin l_1 = +48;
				 l_2 = +53; end
		41271: begin l_1 = +48;
				 l_2 = -53; end
		9590: begin l_1 = -48;
				 l_2 = +53; end
		47215: begin l_1 = -48;
				 l_2 = -53; end
		10264: begin l_1 = +48;
				 l_2 = +54; end
		34653: begin l_1 = +48;
				 l_2 = -54; end
		16208: begin l_1 = -48;
				 l_2 = +54; end
		40597: begin l_1 = -48;
				 l_2 = -54; end
		23500: begin l_1 = +48;
				 l_2 = +55; end
		21417: begin l_1 = +48;
				 l_2 = -55; end
		29444: begin l_1 = -48;
				 l_2 = +55; end
		27361: begin l_1 = -48;
				 l_2 = -55; end
		49972: begin l_1 = +48;
				 l_2 = +56; end
		45806: begin l_1 = +48;
				 l_2 = -56; end
		5055: begin l_1 = -48;
				 l_2 = +56; end
		889: begin l_1 = -48;
				 l_2 = -56; end
		1194: begin l_1 = +48;
				 l_2 = +57; end
		43723: begin l_1 = +48;
				 l_2 = -57; end
		7138: begin l_1 = -48;
				 l_2 = +57; end
		49667: begin l_1 = -48;
				 l_2 = -57; end
		5360: begin l_1 = +48;
				 l_2 = +58; end
		39557: begin l_1 = +48;
				 l_2 = -58; end
		11304: begin l_1 = -48;
				 l_2 = +58; end
		45501: begin l_1 = -48;
				 l_2 = -58; end
		13692: begin l_1 = +48;
				 l_2 = +59; end
		31225: begin l_1 = +48;
				 l_2 = -59; end
		19636: begin l_1 = -48;
				 l_2 = +59; end
		37169: begin l_1 = -48;
				 l_2 = -59; end
		30356: begin l_1 = +48;
				 l_2 = +60; end
		14561: begin l_1 = +48;
				 l_2 = -60; end
		36300: begin l_1 = -48;
				 l_2 = +60; end
		20505: begin l_1 = -48;
				 l_2 = -60; end
		12823: begin l_1 = +48;
				 l_2 = +61; end
		32094: begin l_1 = +48;
				 l_2 = -61; end
		18767: begin l_1 = -48;
				 l_2 = +61; end
		38038: begin l_1 = -48;
				 l_2 = -61; end
		28618: begin l_1 = +48;
				 l_2 = +62; end
		16299: begin l_1 = +48;
				 l_2 = -62; end
		34562: begin l_1 = -48;
				 l_2 = +62; end
		22243: begin l_1 = -48;
				 l_2 = -62; end
		9347: begin l_1 = +48;
				 l_2 = +63; end
		35570: begin l_1 = +48;
				 l_2 = -63; end
		15291: begin l_1 = -48;
				 l_2 = +63; end
		41514: begin l_1 = -48;
				 l_2 = -63; end
		21666: begin l_1 = +48;
				 l_2 = +64; end
		23251: begin l_1 = +48;
				 l_2 = -64; end
		27610: begin l_1 = -48;
				 l_2 = +64; end
		29195: begin l_1 = -48;
				 l_2 = -64; end
		46304: begin l_1 = +48;
				 l_2 = +65; end
		49474: begin l_1 = +48;
				 l_2 = -65; end
		1387: begin l_1 = -48;
				 l_2 = +65; end
		4557: begin l_1 = -48;
				 l_2 = -65; end
		44719: begin l_1 = +48;
				 l_2 = +66; end
		198: begin l_1 = +48;
				 l_2 = -66; end
		50663: begin l_1 = -48;
				 l_2 = +66; end
		6142: begin l_1 = -48;
				 l_2 = -66; end
		41549: begin l_1 = +48;
				 l_2 = +67; end
		3368: begin l_1 = +48;
				 l_2 = -67; end
		47493: begin l_1 = -48;
				 l_2 = +67; end
		9312: begin l_1 = -48;
				 l_2 = -67; end
		35209: begin l_1 = +48;
				 l_2 = +68; end
		9708: begin l_1 = +48;
				 l_2 = -68; end
		41153: begin l_1 = -48;
				 l_2 = +68; end
		15652: begin l_1 = -48;
				 l_2 = -68; end
		33029: begin l_1 = -49;
				 l_2 = +51; end
		17832: begin l_1 = -49;
				 l_2 = -50; end
		21141: begin l_1 = +49;
				 l_2 = +51; end
		29720: begin l_1 = -49;
				 l_2 = -51; end
		48226: begin l_1 = +49;
				 l_2 = +52; end
		41608: begin l_1 = +49;
				 l_2 = -52; end
		9253: begin l_1 = -49;
				 l_2 = +52; end
		2635: begin l_1 = -49;
				 l_2 = -52; end
		674: begin l_1 = +49;
				 l_2 = +53; end
		38299: begin l_1 = +49;
				 l_2 = -53; end
		12562: begin l_1 = -49;
				 l_2 = +53; end
		50187: begin l_1 = -49;
				 l_2 = -53; end
		7292: begin l_1 = +49;
				 l_2 = +54; end
		31681: begin l_1 = +49;
				 l_2 = -54; end
		19180: begin l_1 = -49;
				 l_2 = +54; end
		43569: begin l_1 = -49;
				 l_2 = -54; end
		20528: begin l_1 = +49;
				 l_2 = +55; end
		18445: begin l_1 = +49;
				 l_2 = -55; end
		32416: begin l_1 = -49;
				 l_2 = +55; end
		30333: begin l_1 = -49;
				 l_2 = -55; end
		47000: begin l_1 = +49;
				 l_2 = +56; end
		42834: begin l_1 = +49;
				 l_2 = -56; end
		8027: begin l_1 = -49;
				 l_2 = +56; end
		3861: begin l_1 = -49;
				 l_2 = -56; end
		49083: begin l_1 = +49;
				 l_2 = +57; end
		40751: begin l_1 = +49;
				 l_2 = -57; end
		10110: begin l_1 = -49;
				 l_2 = +57; end
		1778: begin l_1 = -49;
				 l_2 = -57; end
		2388: begin l_1 = +49;
				 l_2 = +58; end
		36585: begin l_1 = +49;
				 l_2 = -58; end
		14276: begin l_1 = -49;
				 l_2 = +58; end
		48473: begin l_1 = -49;
				 l_2 = -58; end
		10720: begin l_1 = +49;
				 l_2 = +59; end
		28253: begin l_1 = +49;
				 l_2 = -59; end
		22608: begin l_1 = -49;
				 l_2 = +59; end
		40141: begin l_1 = -49;
				 l_2 = -59; end
		27384: begin l_1 = +49;
				 l_2 = +60; end
		11589: begin l_1 = +49;
				 l_2 = -60; end
		39272: begin l_1 = -49;
				 l_2 = +60; end
		23477: begin l_1 = -49;
				 l_2 = -60; end
		9851: begin l_1 = +49;
				 l_2 = +61; end
		29122: begin l_1 = +49;
				 l_2 = -61; end
		21739: begin l_1 = -49;
				 l_2 = +61; end
		41010: begin l_1 = -49;
				 l_2 = -61; end
		25646: begin l_1 = +49;
				 l_2 = +62; end
		13327: begin l_1 = +49;
				 l_2 = -62; end
		37534: begin l_1 = -49;
				 l_2 = +62; end
		25215: begin l_1 = -49;
				 l_2 = -62; end
		6375: begin l_1 = +49;
				 l_2 = +63; end
		32598: begin l_1 = +49;
				 l_2 = -63; end
		18263: begin l_1 = -49;
				 l_2 = +63; end
		44486: begin l_1 = -49;
				 l_2 = -63; end
		18694: begin l_1 = +49;
				 l_2 = +64; end
		20279: begin l_1 = +49;
				 l_2 = -64; end
		30582: begin l_1 = -49;
				 l_2 = +64; end
		32167: begin l_1 = -49;
				 l_2 = -64; end
		43332: begin l_1 = +49;
				 l_2 = +65; end
		46502: begin l_1 = +49;
				 l_2 = -65; end
		4359: begin l_1 = -49;
				 l_2 = +65; end
		7529: begin l_1 = -49;
				 l_2 = -65; end
		41747: begin l_1 = +49;
				 l_2 = +66; end
		48087: begin l_1 = +49;
				 l_2 = -66; end
		2774: begin l_1 = -49;
				 l_2 = +66; end
		9114: begin l_1 = -49;
				 l_2 = -66; end
		38577: begin l_1 = +49;
				 l_2 = +67; end
		396: begin l_1 = +49;
				 l_2 = -67; end
		50465: begin l_1 = -49;
				 l_2 = +67; end
		12284: begin l_1 = -49;
				 l_2 = -67; end
		32237: begin l_1 = +49;
				 l_2 = +68; end
		6736: begin l_1 = +49;
				 l_2 = -68; end
		44125: begin l_1 = -49;
				 l_2 = +68; end
		18624: begin l_1 = -49;
				 l_2 = -68; end
		15197: begin l_1 = -50;
				 l_2 = +52; end
		35664: begin l_1 = -50;
				 l_2 = -51; end
		42282: begin l_1 = +50;
				 l_2 = +52; end
		8579: begin l_1 = -50;
				 l_2 = -52; end
		45591: begin l_1 = +50;
				 l_2 = +53; end
		32355: begin l_1 = +50;
				 l_2 = -53; end
		18506: begin l_1 = -50;
				 l_2 = +53; end
		5270: begin l_1 = -50;
				 l_2 = -53; end
		1348: begin l_1 = +50;
				 l_2 = +54; end
		25737: begin l_1 = +50;
				 l_2 = -54; end
		25124: begin l_1 = -50;
				 l_2 = +54; end
		49513: begin l_1 = -50;
				 l_2 = -54; end
		14584: begin l_1 = +50;
				 l_2 = +55; end
		12501: begin l_1 = +50;
				 l_2 = -55; end
		38360: begin l_1 = -50;
				 l_2 = +55; end
		36277: begin l_1 = -50;
				 l_2 = -55; end
		41056: begin l_1 = +50;
				 l_2 = +56; end
		36890: begin l_1 = +50;
				 l_2 = -56; end
		13971: begin l_1 = -50;
				 l_2 = +56; end
		9805: begin l_1 = -50;
				 l_2 = -56; end
		43139: begin l_1 = +50;
				 l_2 = +57; end
		34807: begin l_1 = +50;
				 l_2 = -57; end
		16054: begin l_1 = -50;
				 l_2 = +57; end
		7722: begin l_1 = -50;
				 l_2 = -57; end
		47305: begin l_1 = +50;
				 l_2 = +58; end
		30641: begin l_1 = +50;
				 l_2 = -58; end
		20220: begin l_1 = -50;
				 l_2 = +58; end
		3556: begin l_1 = -50;
				 l_2 = -58; end
		4776: begin l_1 = +50;
				 l_2 = +59; end
		22309: begin l_1 = +50;
				 l_2 = -59; end
		28552: begin l_1 = -50;
				 l_2 = +59; end
		46085: begin l_1 = -50;
				 l_2 = -59; end
		21440: begin l_1 = +50;
				 l_2 = +60; end
		5645: begin l_1 = +50;
				 l_2 = -60; end
		45216: begin l_1 = -50;
				 l_2 = +60; end
		29421: begin l_1 = -50;
				 l_2 = -60; end
		3907: begin l_1 = +50;
				 l_2 = +61; end
		23178: begin l_1 = +50;
				 l_2 = -61; end
		27683: begin l_1 = -50;
				 l_2 = +61; end
		46954: begin l_1 = -50;
				 l_2 = -61; end
		19702: begin l_1 = +50;
				 l_2 = +62; end
		7383: begin l_1 = +50;
				 l_2 = -62; end
		43478: begin l_1 = -50;
				 l_2 = +62; end
		31159: begin l_1 = -50;
				 l_2 = -62; end
		431: begin l_1 = +50;
				 l_2 = +63; end
		26654: begin l_1 = +50;
				 l_2 = -63; end
		24207: begin l_1 = -50;
				 l_2 = +63; end
		50430: begin l_1 = -50;
				 l_2 = -63; end
		12750: begin l_1 = +50;
				 l_2 = +64; end
		14335: begin l_1 = +50;
				 l_2 = -64; end
		36526: begin l_1 = -50;
				 l_2 = +64; end
		38111: begin l_1 = -50;
				 l_2 = -64; end
		37388: begin l_1 = +50;
				 l_2 = +65; end
		40558: begin l_1 = +50;
				 l_2 = -65; end
		10303: begin l_1 = -50;
				 l_2 = +65; end
		13473: begin l_1 = -50;
				 l_2 = -65; end
		35803: begin l_1 = +50;
				 l_2 = +66; end
		42143: begin l_1 = +50;
				 l_2 = -66; end
		8718: begin l_1 = -50;
				 l_2 = +66; end
		15058: begin l_1 = -50;
				 l_2 = -66; end
		32633: begin l_1 = +50;
				 l_2 = +67; end
		45313: begin l_1 = +50;
				 l_2 = -67; end
		5548: begin l_1 = -50;
				 l_2 = +67; end
		18228: begin l_1 = -50;
				 l_2 = -67; end
		26293: begin l_1 = +50;
				 l_2 = +68; end
		792: begin l_1 = +50;
				 l_2 = -68; end
		50069: begin l_1 = -50;
				 l_2 = +68; end
		24568: begin l_1 = -50;
				 l_2 = -68; end
		30394: begin l_1 = -51;
				 l_2 = +53; end
		20467: begin l_1 = -51;
				 l_2 = -52; end
		33703: begin l_1 = +51;
				 l_2 = +53; end
		17158: begin l_1 = -51;
				 l_2 = -53; end
		40321: begin l_1 = +51;
				 l_2 = +54; end
		13849: begin l_1 = +51;
				 l_2 = -54; end
		37012: begin l_1 = -51;
				 l_2 = +54; end
		10540: begin l_1 = -51;
				 l_2 = -54; end
		2696: begin l_1 = +51;
				 l_2 = +55; end
		613: begin l_1 = +51;
				 l_2 = -55; end
		50248: begin l_1 = -51;
				 l_2 = +55; end
		48165: begin l_1 = -51;
				 l_2 = -55; end
		29168: begin l_1 = +51;
				 l_2 = +56; end
		25002: begin l_1 = +51;
				 l_2 = -56; end
		25859: begin l_1 = -51;
				 l_2 = +56; end
		21693: begin l_1 = -51;
				 l_2 = -56; end
		31251: begin l_1 = +51;
				 l_2 = +57; end
		22919: begin l_1 = +51;
				 l_2 = -57; end
		27942: begin l_1 = -51;
				 l_2 = +57; end
		19610: begin l_1 = -51;
				 l_2 = -57; end
		35417: begin l_1 = +51;
				 l_2 = +58; end
		18753: begin l_1 = +51;
				 l_2 = -58; end
		32108: begin l_1 = -51;
				 l_2 = +58; end
		15444: begin l_1 = -51;
				 l_2 = -58; end
		43749: begin l_1 = +51;
				 l_2 = +59; end
		10421: begin l_1 = +51;
				 l_2 = -59; end
		40440: begin l_1 = -51;
				 l_2 = +59; end
		7112: begin l_1 = -51;
				 l_2 = -59; end
		9552: begin l_1 = +51;
				 l_2 = +60; end
		44618: begin l_1 = +51;
				 l_2 = -60; end
		6243: begin l_1 = -51;
				 l_2 = +60; end
		41309: begin l_1 = -51;
				 l_2 = -60; end
		42880: begin l_1 = +51;
				 l_2 = +61; end
		11290: begin l_1 = +51;
				 l_2 = -61; end
		39571: begin l_1 = -51;
				 l_2 = +61; end
		7981: begin l_1 = -51;
				 l_2 = -61; end
		7814: begin l_1 = +51;
				 l_2 = +62; end
		46356: begin l_1 = +51;
				 l_2 = -62; end
		4505: begin l_1 = -51;
				 l_2 = +62; end
		43047: begin l_1 = -51;
				 l_2 = -62; end
		39404: begin l_1 = +51;
				 l_2 = +63; end
		14766: begin l_1 = +51;
				 l_2 = -63; end
		36095: begin l_1 = -51;
				 l_2 = +63; end
		11457: begin l_1 = -51;
				 l_2 = -63; end
		862: begin l_1 = +51;
				 l_2 = +64; end
		2447: begin l_1 = +51;
				 l_2 = -64; end
		48414: begin l_1 = -51;
				 l_2 = +64; end
		49999: begin l_1 = -51;
				 l_2 = -64; end
		25500: begin l_1 = +51;
				 l_2 = +65; end
		28670: begin l_1 = +51;
				 l_2 = -65; end
		22191: begin l_1 = -51;
				 l_2 = +65; end
		25361: begin l_1 = -51;
				 l_2 = -65; end
		23915: begin l_1 = +51;
				 l_2 = +66; end
		30255: begin l_1 = +51;
				 l_2 = -66; end
		20606: begin l_1 = -51;
				 l_2 = +66; end
		26946: begin l_1 = -51;
				 l_2 = -66; end
		20745: begin l_1 = +51;
				 l_2 = +67; end
		33425: begin l_1 = +51;
				 l_2 = -67; end
		17436: begin l_1 = -51;
				 l_2 = +67; end
		30116: begin l_1 = -51;
				 l_2 = -67; end
		14405: begin l_1 = +51;
				 l_2 = +68; end
		39765: begin l_1 = +51;
				 l_2 = -68; end
		11096: begin l_1 = -51;
				 l_2 = +68; end
		36456: begin l_1 = -51;
				 l_2 = -68; end
		9927: begin l_1 = -52;
				 l_2 = +54; end
		40934: begin l_1 = -52;
				 l_2 = -53; end
		16545: begin l_1 = +52;
				 l_2 = +54; end
		34316: begin l_1 = -52;
				 l_2 = -54; end
		29781: begin l_1 = +52;
				 l_2 = +55; end
		27698: begin l_1 = +52;
				 l_2 = -55; end
		23163: begin l_1 = -52;
				 l_2 = +55; end
		21080: begin l_1 = -52;
				 l_2 = -55; end
		5392: begin l_1 = +52;
				 l_2 = +56; end
		1226: begin l_1 = +52;
				 l_2 = -56; end
		49635: begin l_1 = -52;
				 l_2 = +56; end
		45469: begin l_1 = -52;
				 l_2 = -56; end
		7475: begin l_1 = +52;
				 l_2 = +57; end
		50004: begin l_1 = +52;
				 l_2 = -57; end
		857: begin l_1 = -52;
				 l_2 = +57; end
		43386: begin l_1 = -52;
				 l_2 = -57; end
		11641: begin l_1 = +52;
				 l_2 = +58; end
		45838: begin l_1 = +52;
				 l_2 = -58; end
		5023: begin l_1 = -52;
				 l_2 = +58; end
		39220: begin l_1 = -52;
				 l_2 = -58; end
		19973: begin l_1 = +52;
				 l_2 = +59; end
		37506: begin l_1 = +52;
				 l_2 = -59; end
		13355: begin l_1 = -52;
				 l_2 = +59; end
		30888: begin l_1 = -52;
				 l_2 = -59; end
		36637: begin l_1 = +52;
				 l_2 = +60; end
		20842: begin l_1 = +52;
				 l_2 = -60; end
		30019: begin l_1 = -52;
				 l_2 = +60; end
		14224: begin l_1 = -52;
				 l_2 = -60; end
		19104: begin l_1 = +52;
				 l_2 = +61; end
		38375: begin l_1 = +52;
				 l_2 = -61; end
		12486: begin l_1 = -52;
				 l_2 = +61; end
		31757: begin l_1 = -52;
				 l_2 = -61; end
		34899: begin l_1 = +52;
				 l_2 = +62; end
		22580: begin l_1 = +52;
				 l_2 = -62; end
		28281: begin l_1 = -52;
				 l_2 = +62; end
		15962: begin l_1 = -52;
				 l_2 = -62; end
		15628: begin l_1 = +52;
				 l_2 = +63; end
		41851: begin l_1 = +52;
				 l_2 = -63; end
		9010: begin l_1 = -52;
				 l_2 = +63; end
		35233: begin l_1 = -52;
				 l_2 = -63; end
		27947: begin l_1 = +52;
				 l_2 = +64; end
		29532: begin l_1 = +52;
				 l_2 = -64; end
		21329: begin l_1 = -52;
				 l_2 = +64; end
		22914: begin l_1 = -52;
				 l_2 = -64; end
		1724: begin l_1 = +52;
				 l_2 = +65; end
		4894: begin l_1 = +52;
				 l_2 = -65; end
		45967: begin l_1 = -52;
				 l_2 = +65; end
		49137: begin l_1 = -52;
				 l_2 = -65; end
		139: begin l_1 = +52;
				 l_2 = +66; end
		6479: begin l_1 = +52;
				 l_2 = -66; end
		44382: begin l_1 = -52;
				 l_2 = +66; end
		50722: begin l_1 = -52;
				 l_2 = -66; end
		47830: begin l_1 = +52;
				 l_2 = +67; end
		9649: begin l_1 = +52;
				 l_2 = -67; end
		41212: begin l_1 = -52;
				 l_2 = +67; end
		3031: begin l_1 = -52;
				 l_2 = -67; end
		41490: begin l_1 = +52;
				 l_2 = +68; end
		15989: begin l_1 = +52;
				 l_2 = -68; end
		34872: begin l_1 = -52;
				 l_2 = +68; end
		9371: begin l_1 = -52;
				 l_2 = -68; end
		19854: begin l_1 = -53;
				 l_2 = +55; end
		31007: begin l_1 = -53;
				 l_2 = -54; end
		33090: begin l_1 = +53;
				 l_2 = +55; end
		17771: begin l_1 = -53;
				 l_2 = -55; end
		8701: begin l_1 = +53;
				 l_2 = +56; end
		4535: begin l_1 = +53;
				 l_2 = -56; end
		46326: begin l_1 = -53;
				 l_2 = +56; end
		42160: begin l_1 = -53;
				 l_2 = -56; end
		10784: begin l_1 = +53;
				 l_2 = +57; end
		2452: begin l_1 = +53;
				 l_2 = -57; end
		48409: begin l_1 = -53;
				 l_2 = +57; end
		40077: begin l_1 = -53;
				 l_2 = -57; end
		14950: begin l_1 = +53;
				 l_2 = +58; end
		49147: begin l_1 = +53;
				 l_2 = -58; end
		1714: begin l_1 = -53;
				 l_2 = +58; end
		35911: begin l_1 = -53;
				 l_2 = -58; end
		23282: begin l_1 = +53;
				 l_2 = +59; end
		40815: begin l_1 = +53;
				 l_2 = -59; end
		10046: begin l_1 = -53;
				 l_2 = +59; end
		27579: begin l_1 = -53;
				 l_2 = -59; end
		39946: begin l_1 = +53;
				 l_2 = +60; end
		24151: begin l_1 = +53;
				 l_2 = -60; end
		26710: begin l_1 = -53;
				 l_2 = +60; end
		10915: begin l_1 = -53;
				 l_2 = -60; end
		22413: begin l_1 = +53;
				 l_2 = +61; end
		41684: begin l_1 = +53;
				 l_2 = -61; end
		9177: begin l_1 = -53;
				 l_2 = +61; end
		28448: begin l_1 = -53;
				 l_2 = -61; end
		38208: begin l_1 = +53;
				 l_2 = +62; end
		25889: begin l_1 = +53;
				 l_2 = -62; end
		24972: begin l_1 = -53;
				 l_2 = +62; end
		12653: begin l_1 = -53;
				 l_2 = -62; end
		18937: begin l_1 = +53;
				 l_2 = +63; end
		45160: begin l_1 = +53;
				 l_2 = -63; end
		5701: begin l_1 = -53;
				 l_2 = +63; end
		31924: begin l_1 = -53;
				 l_2 = -63; end
		31256: begin l_1 = +53;
				 l_2 = +64; end
		32841: begin l_1 = +53;
				 l_2 = -64; end
		18020: begin l_1 = -53;
				 l_2 = +64; end
		19605: begin l_1 = -53;
				 l_2 = -64; end
		5033: begin l_1 = +53;
				 l_2 = +65; end
		8203: begin l_1 = +53;
				 l_2 = -65; end
		42658: begin l_1 = -53;
				 l_2 = +65; end
		45828: begin l_1 = -53;
				 l_2 = -65; end
		3448: begin l_1 = +53;
				 l_2 = +66; end
		9788: begin l_1 = +53;
				 l_2 = -66; end
		41073: begin l_1 = -53;
				 l_2 = +66; end
		47413: begin l_1 = -53;
				 l_2 = -66; end
		278: begin l_1 = +53;
				 l_2 = +67; end
		12958: begin l_1 = +53;
				 l_2 = -67; end
		37903: begin l_1 = -53;
				 l_2 = +67; end
		50583: begin l_1 = -53;
				 l_2 = -67; end
		44799: begin l_1 = +53;
				 l_2 = +68; end
		19298: begin l_1 = +53;
				 l_2 = -68; end
		31563: begin l_1 = -53;
				 l_2 = +68; end
		6062: begin l_1 = -53;
				 l_2 = -68; end
		39708: begin l_1 = -54;
				 l_2 = +56; end
		11153: begin l_1 = -54;
				 l_2 = -55; end
		15319: begin l_1 = +54;
				 l_2 = +56; end
		35542: begin l_1 = -54;
				 l_2 = -56; end
		17402: begin l_1 = +54;
				 l_2 = +57; end
		9070: begin l_1 = +54;
				 l_2 = -57; end
		41791: begin l_1 = -54;
				 l_2 = +57; end
		33459: begin l_1 = -54;
				 l_2 = -57; end
		21568: begin l_1 = +54;
				 l_2 = +58; end
		4904: begin l_1 = +54;
				 l_2 = -58; end
		45957: begin l_1 = -54;
				 l_2 = +58; end
		29293: begin l_1 = -54;
				 l_2 = -58; end
		29900: begin l_1 = +54;
				 l_2 = +59; end
		47433: begin l_1 = +54;
				 l_2 = -59; end
		3428: begin l_1 = -54;
				 l_2 = +59; end
		20961: begin l_1 = -54;
				 l_2 = -59; end
		46564: begin l_1 = +54;
				 l_2 = +60; end
		30769: begin l_1 = +54;
				 l_2 = -60; end
		20092: begin l_1 = -54;
				 l_2 = +60; end
		4297: begin l_1 = -54;
				 l_2 = -60; end
		29031: begin l_1 = +54;
				 l_2 = +61; end
		48302: begin l_1 = +54;
				 l_2 = -61; end
		2559: begin l_1 = -54;
				 l_2 = +61; end
		21830: begin l_1 = -54;
				 l_2 = -61; end
		44826: begin l_1 = +54;
				 l_2 = +62; end
		32507: begin l_1 = +54;
				 l_2 = -62; end
		18354: begin l_1 = -54;
				 l_2 = +62; end
		6035: begin l_1 = -54;
				 l_2 = -62; end
		25555: begin l_1 = +54;
				 l_2 = +63; end
		917: begin l_1 = +54;
				 l_2 = -63; end
		49944: begin l_1 = -54;
				 l_2 = +63; end
		25306: begin l_1 = -54;
				 l_2 = -63; end
		37874: begin l_1 = +54;
				 l_2 = +64; end
		39459: begin l_1 = +54;
				 l_2 = -64; end
		11402: begin l_1 = -54;
				 l_2 = +64; end
		12987: begin l_1 = -54;
				 l_2 = -64; end
		11651: begin l_1 = +54;
				 l_2 = +65; end
		14821: begin l_1 = +54;
				 l_2 = -65; end
		36040: begin l_1 = -54;
				 l_2 = +65; end
		39210: begin l_1 = -54;
				 l_2 = -65; end
		10066: begin l_1 = +54;
				 l_2 = +66; end
		16406: begin l_1 = +54;
				 l_2 = -66; end
		34455: begin l_1 = -54;
				 l_2 = +66; end
		40795: begin l_1 = -54;
				 l_2 = -66; end
		6896: begin l_1 = +54;
				 l_2 = +67; end
		19576: begin l_1 = +54;
				 l_2 = -67; end
		31285: begin l_1 = -54;
				 l_2 = +67; end
		43965: begin l_1 = -54;
				 l_2 = -67; end
		556: begin l_1 = +54;
				 l_2 = +68; end
		25916: begin l_1 = +54;
				 l_2 = -68; end
		24945: begin l_1 = -54;
				 l_2 = +68; end
		50305: begin l_1 = -54;
				 l_2 = -68; end
		28555: begin l_1 = -55;
				 l_2 = +57; end
		22306: begin l_1 = -55;
				 l_2 = -56; end
		30638: begin l_1 = +55;
				 l_2 = +57; end
		20223: begin l_1 = -55;
				 l_2 = -57; end
		34804: begin l_1 = +55;
				 l_2 = +58; end
		18140: begin l_1 = +55;
				 l_2 = -58; end
		32721: begin l_1 = -55;
				 l_2 = +58; end
		16057: begin l_1 = -55;
				 l_2 = -58; end
		43136: begin l_1 = +55;
				 l_2 = +59; end
		9808: begin l_1 = +55;
				 l_2 = -59; end
		41053: begin l_1 = -55;
				 l_2 = +59; end
		7725: begin l_1 = -55;
				 l_2 = -59; end
		8939: begin l_1 = +55;
				 l_2 = +60; end
		44005: begin l_1 = +55;
				 l_2 = -60; end
		6856: begin l_1 = -55;
				 l_2 = +60; end
		41922: begin l_1 = -55;
				 l_2 = -60; end
		42267: begin l_1 = +55;
				 l_2 = +61; end
		10677: begin l_1 = +55;
				 l_2 = -61; end
		40184: begin l_1 = -55;
				 l_2 = +61; end
		8594: begin l_1 = -55;
				 l_2 = -61; end
		7201: begin l_1 = +55;
				 l_2 = +62; end
		45743: begin l_1 = +55;
				 l_2 = -62; end
		5118: begin l_1 = -55;
				 l_2 = +62; end
		43660: begin l_1 = -55;
				 l_2 = -62; end
		38791: begin l_1 = +55;
				 l_2 = +63; end
		14153: begin l_1 = +55;
				 l_2 = -63; end
		36708: begin l_1 = -55;
				 l_2 = +63; end
		12070: begin l_1 = -55;
				 l_2 = -63; end
		249: begin l_1 = +55;
				 l_2 = +64; end
		1834: begin l_1 = +55;
				 l_2 = -64; end
		49027: begin l_1 = -55;
				 l_2 = +64; end
		50612: begin l_1 = -55;
				 l_2 = -64; end
		24887: begin l_1 = +55;
				 l_2 = +65; end
		28057: begin l_1 = +55;
				 l_2 = -65; end
		22804: begin l_1 = -55;
				 l_2 = +65; end
		25974: begin l_1 = -55;
				 l_2 = -65; end
		23302: begin l_1 = +55;
				 l_2 = +66; end
		29642: begin l_1 = +55;
				 l_2 = -66; end
		21219: begin l_1 = -55;
				 l_2 = +66; end
		27559: begin l_1 = -55;
				 l_2 = -66; end
		20132: begin l_1 = +55;
				 l_2 = +67; end
		32812: begin l_1 = +55;
				 l_2 = -67; end
		18049: begin l_1 = -55;
				 l_2 = +67; end
		30729: begin l_1 = -55;
				 l_2 = -67; end
		13792: begin l_1 = +55;
				 l_2 = +68; end
		39152: begin l_1 = +55;
				 l_2 = -68; end
		11709: begin l_1 = -55;
				 l_2 = +68; end
		37069: begin l_1 = -55;
				 l_2 = -68; end
		6249: begin l_1 = -56;
				 l_2 = +58; end
		44612: begin l_1 = -56;
				 l_2 = -57; end
		10415: begin l_1 = +56;
				 l_2 = +58; end
		40446: begin l_1 = -56;
				 l_2 = -58; end
		18747: begin l_1 = +56;
				 l_2 = +59; end
		36280: begin l_1 = +56;
				 l_2 = -59; end
		14581: begin l_1 = -56;
				 l_2 = +59; end
		32114: begin l_1 = -56;
				 l_2 = -59; end
		35411: begin l_1 = +56;
				 l_2 = +60; end
		19616: begin l_1 = +56;
				 l_2 = -60; end
		31245: begin l_1 = -56;
				 l_2 = +60; end
		15450: begin l_1 = -56;
				 l_2 = -60; end
		17878: begin l_1 = +56;
				 l_2 = +61; end
		37149: begin l_1 = +56;
				 l_2 = -61; end
		13712: begin l_1 = -56;
				 l_2 = +61; end
		32983: begin l_1 = -56;
				 l_2 = -61; end
		33673: begin l_1 = +56;
				 l_2 = +62; end
		21354: begin l_1 = +56;
				 l_2 = -62; end
		29507: begin l_1 = -56;
				 l_2 = +62; end
		17188: begin l_1 = -56;
				 l_2 = -62; end
		14402: begin l_1 = +56;
				 l_2 = +63; end
		40625: begin l_1 = +56;
				 l_2 = -63; end
		10236: begin l_1 = -56;
				 l_2 = +63; end
		36459: begin l_1 = -56;
				 l_2 = -63; end
		26721: begin l_1 = +56;
				 l_2 = +64; end
		28306: begin l_1 = +56;
				 l_2 = -64; end
		22555: begin l_1 = -56;
				 l_2 = +64; end
		24140: begin l_1 = -56;
				 l_2 = -64; end
		498: begin l_1 = +56;
				 l_2 = +65; end
		3668: begin l_1 = +56;
				 l_2 = -65; end
		47193: begin l_1 = -56;
				 l_2 = +65; end
		50363: begin l_1 = -56;
				 l_2 = -65; end
		49774: begin l_1 = +56;
				 l_2 = +66; end
		5253: begin l_1 = +56;
				 l_2 = -66; end
		45608: begin l_1 = -56;
				 l_2 = +66; end
		1087: begin l_1 = -56;
				 l_2 = -66; end
		46604: begin l_1 = +56;
				 l_2 = +67; end
		8423: begin l_1 = +56;
				 l_2 = -67; end
		42438: begin l_1 = -56;
				 l_2 = +67; end
		4257: begin l_1 = -56;
				 l_2 = -67; end
		40264: begin l_1 = +56;
				 l_2 = +68; end
		14763: begin l_1 = +56;
				 l_2 = -68; end
		36098: begin l_1 = -56;
				 l_2 = +68; end
		10597: begin l_1 = -56;
				 l_2 = -68; end
		12498: begin l_1 = -57;
				 l_2 = +59; end
		38363: begin l_1 = -57;
				 l_2 = -58; end
		20830: begin l_1 = +57;
				 l_2 = +59; end
		30031: begin l_1 = -57;
				 l_2 = -59; end
		37494: begin l_1 = +57;
				 l_2 = +60; end
		21699: begin l_1 = +57;
				 l_2 = -60; end
		29162: begin l_1 = -57;
				 l_2 = +60; end
		13367: begin l_1 = -57;
				 l_2 = -60; end
		19961: begin l_1 = +57;
				 l_2 = +61; end
		39232: begin l_1 = +57;
				 l_2 = -61; end
		11629: begin l_1 = -57;
				 l_2 = +61; end
		30900: begin l_1 = -57;
				 l_2 = -61; end
		35756: begin l_1 = +57;
				 l_2 = +62; end
		23437: begin l_1 = +57;
				 l_2 = -62; end
		27424: begin l_1 = -57;
				 l_2 = +62; end
		15105: begin l_1 = -57;
				 l_2 = -62; end
		16485: begin l_1 = +57;
				 l_2 = +63; end
		42708: begin l_1 = +57;
				 l_2 = -63; end
		8153: begin l_1 = -57;
				 l_2 = +63; end
		34376: begin l_1 = -57;
				 l_2 = -63; end
		28804: begin l_1 = +57;
				 l_2 = +64; end
		30389: begin l_1 = +57;
				 l_2 = -64; end
		20472: begin l_1 = -57;
				 l_2 = +64; end
		22057: begin l_1 = -57;
				 l_2 = -64; end
		2581: begin l_1 = +57;
				 l_2 = +65; end
		5751: begin l_1 = +57;
				 l_2 = -65; end
		45110: begin l_1 = -57;
				 l_2 = +65; end
		48280: begin l_1 = -57;
				 l_2 = -65; end
		996: begin l_1 = +57;
				 l_2 = +66; end
		7336: begin l_1 = +57;
				 l_2 = -66; end
		43525: begin l_1 = -57;
				 l_2 = +66; end
		49865: begin l_1 = -57;
				 l_2 = -66; end
		48687: begin l_1 = +57;
				 l_2 = +67; end
		10506: begin l_1 = +57;
				 l_2 = -67; end
		40355: begin l_1 = -57;
				 l_2 = +67; end
		2174: begin l_1 = -57;
				 l_2 = -67; end
		42347: begin l_1 = +57;
				 l_2 = +68; end
		16846: begin l_1 = +57;
				 l_2 = -68; end
		34015: begin l_1 = -57;
				 l_2 = +68; end
		8514: begin l_1 = -57;
				 l_2 = -68; end
		24996: begin l_1 = -58;
				 l_2 = +60; end
		25865: begin l_1 = -58;
				 l_2 = -59; end
		41660: begin l_1 = +58;
				 l_2 = +60; end
		9201: begin l_1 = -58;
				 l_2 = -60; end
		24127: begin l_1 = +58;
				 l_2 = +61; end
		43398: begin l_1 = +58;
				 l_2 = -61; end
		7463: begin l_1 = -58;
				 l_2 = +61; end
		26734: begin l_1 = -58;
				 l_2 = -61; end
		39922: begin l_1 = +58;
				 l_2 = +62; end
		27603: begin l_1 = +58;
				 l_2 = -62; end
		23258: begin l_1 = -58;
				 l_2 = +62; end
		10939: begin l_1 = -58;
				 l_2 = -62; end
		20651: begin l_1 = +58;
				 l_2 = +63; end
		46874: begin l_1 = +58;
				 l_2 = -63; end
		3987: begin l_1 = -58;
				 l_2 = +63; end
		30210: begin l_1 = -58;
				 l_2 = -63; end
		32970: begin l_1 = +58;
				 l_2 = +64; end
		34555: begin l_1 = +58;
				 l_2 = -64; end
		16306: begin l_1 = -58;
				 l_2 = +64; end
		17891: begin l_1 = -58;
				 l_2 = -64; end
		6747: begin l_1 = +58;
				 l_2 = +65; end
		9917: begin l_1 = +58;
				 l_2 = -65; end
		40944: begin l_1 = -58;
				 l_2 = +65; end
		44114: begin l_1 = -58;
				 l_2 = -65; end
		5162: begin l_1 = +58;
				 l_2 = +66; end
		11502: begin l_1 = +58;
				 l_2 = -66; end
		39359: begin l_1 = -58;
				 l_2 = +66; end
		45699: begin l_1 = -58;
				 l_2 = -66; end
		1992: begin l_1 = +58;
				 l_2 = +67; end
		14672: begin l_1 = +58;
				 l_2 = -67; end
		36189: begin l_1 = -58;
				 l_2 = +67; end
		48869: begin l_1 = -58;
				 l_2 = -67; end
		46513: begin l_1 = +58;
				 l_2 = +68; end
		21012: begin l_1 = +58;
				 l_2 = -68; end
		29849: begin l_1 = -58;
				 l_2 = +68; end
		4348: begin l_1 = -58;
				 l_2 = -68; end
		49992: begin l_1 = -59;
				 l_2 = +61; end
		869: begin l_1 = -59;
				 l_2 = -60; end
		32459: begin l_1 = +59;
				 l_2 = +61; end
		18402: begin l_1 = -59;
				 l_2 = -61; end
		48254: begin l_1 = +59;
				 l_2 = +62; end
		35935: begin l_1 = +59;
				 l_2 = -62; end
		14926: begin l_1 = -59;
				 l_2 = +62; end
		2607: begin l_1 = -59;
				 l_2 = -62; end
		28983: begin l_1 = +59;
				 l_2 = +63; end
		4345: begin l_1 = +59;
				 l_2 = -63; end
		46516: begin l_1 = -59;
				 l_2 = +63; end
		21878: begin l_1 = -59;
				 l_2 = -63; end
		41302: begin l_1 = +59;
				 l_2 = +64; end
		42887: begin l_1 = +59;
				 l_2 = -64; end
		7974: begin l_1 = -59;
				 l_2 = +64; end
		9559: begin l_1 = -59;
				 l_2 = -64; end
		15079: begin l_1 = +59;
				 l_2 = +65; end
		18249: begin l_1 = +59;
				 l_2 = -65; end
		32612: begin l_1 = -59;
				 l_2 = +65; end
		35782: begin l_1 = -59;
				 l_2 = -65; end
		13494: begin l_1 = +59;
				 l_2 = +66; end
		19834: begin l_1 = +59;
				 l_2 = -66; end
		31027: begin l_1 = -59;
				 l_2 = +66; end
		37367: begin l_1 = -59;
				 l_2 = -66; end
		10324: begin l_1 = +59;
				 l_2 = +67; end
		23004: begin l_1 = +59;
				 l_2 = -67; end
		27857: begin l_1 = -59;
				 l_2 = +67; end
		40537: begin l_1 = -59;
				 l_2 = -67; end
		3984: begin l_1 = +59;
				 l_2 = +68; end
		29344: begin l_1 = +59;
				 l_2 = -68; end
		21517: begin l_1 = -59;
				 l_2 = +68; end
		46877: begin l_1 = -59;
				 l_2 = -68; end
		49123: begin l_1 = -60;
				 l_2 = +62; end
		1738: begin l_1 = -60;
				 l_2 = -61; end
		14057: begin l_1 = +60;
				 l_2 = +62; end
		36804: begin l_1 = -60;
				 l_2 = -62; end
		45647: begin l_1 = +60;
				 l_2 = +63; end
		21009: begin l_1 = +60;
				 l_2 = -63; end
		29852: begin l_1 = -60;
				 l_2 = +63; end
		5214: begin l_1 = -60;
				 l_2 = -63; end
		7105: begin l_1 = +60;
				 l_2 = +64; end
		8690: begin l_1 = +60;
				 l_2 = -64; end
		42171: begin l_1 = -60;
				 l_2 = +64; end
		43756: begin l_1 = -60;
				 l_2 = -64; end
		31743: begin l_1 = +60;
				 l_2 = +65; end
		34913: begin l_1 = +60;
				 l_2 = -65; end
		15948: begin l_1 = -60;
				 l_2 = +65; end
		19118: begin l_1 = -60;
				 l_2 = -65; end
		30158: begin l_1 = +60;
				 l_2 = +66; end
		36498: begin l_1 = +60;
				 l_2 = -66; end
		14363: begin l_1 = -60;
				 l_2 = +66; end
		20703: begin l_1 = -60;
				 l_2 = -66; end
		26988: begin l_1 = +60;
				 l_2 = +67; end
		39668: begin l_1 = +60;
				 l_2 = -67; end
		11193: begin l_1 = -60;
				 l_2 = +67; end
		23873: begin l_1 = -60;
				 l_2 = -67; end
		20648: begin l_1 = +60;
				 l_2 = +68; end
		46008: begin l_1 = +60;
				 l_2 = -68; end
		4853: begin l_1 = -60;
				 l_2 = +68; end
		30213: begin l_1 = -60;
				 l_2 = -68; end
		47385: begin l_1 = -61;
				 l_2 = +63; end
		3476: begin l_1 = -61;
				 l_2 = -62; end
		28114: begin l_1 = +61;
				 l_2 = +63; end
		22747: begin l_1 = -61;
				 l_2 = -63; end
		40433: begin l_1 = +61;
				 l_2 = +64; end
		42018: begin l_1 = +61;
				 l_2 = -64; end
		8843: begin l_1 = -61;
				 l_2 = +64; end
		10428: begin l_1 = -61;
				 l_2 = -64; end
		14210: begin l_1 = +61;
				 l_2 = +65; end
		17380: begin l_1 = +61;
				 l_2 = -65; end
		33481: begin l_1 = -61;
				 l_2 = +65; end
		36651: begin l_1 = -61;
				 l_2 = -65; end
		12625: begin l_1 = +61;
				 l_2 = +66; end
		18965: begin l_1 = +61;
				 l_2 = -66; end
		31896: begin l_1 = -61;
				 l_2 = +66; end
		38236: begin l_1 = -61;
				 l_2 = -66; end
		9455: begin l_1 = +61;
				 l_2 = +67; end
		22135: begin l_1 = +61;
				 l_2 = -67; end
		28726: begin l_1 = -61;
				 l_2 = +67; end
		41406: begin l_1 = -61;
				 l_2 = -67; end
		3115: begin l_1 = +61;
				 l_2 = +68; end
		28475: begin l_1 = +61;
				 l_2 = -68; end
		22386: begin l_1 = -61;
				 l_2 = +68; end
		47746: begin l_1 = -61;
				 l_2 = -68; end
		43909: begin l_1 = -62;
				 l_2 = +64; end
		6952: begin l_1 = -62;
				 l_2 = -63; end
		5367: begin l_1 = +62;
				 l_2 = +64; end
		45494: begin l_1 = -62;
				 l_2 = -64; end
		30005: begin l_1 = +62;
				 l_2 = +65; end
		33175: begin l_1 = +62;
				 l_2 = -65; end
		17686: begin l_1 = -62;
				 l_2 = +65; end
		20856: begin l_1 = -62;
				 l_2 = -65; end
		28420: begin l_1 = +62;
				 l_2 = +66; end
		34760: begin l_1 = +62;
				 l_2 = -66; end
		16101: begin l_1 = -62;
				 l_2 = +66; end
		22441: begin l_1 = -62;
				 l_2 = -66; end
		25250: begin l_1 = +62;
				 l_2 = +67; end
		37930: begin l_1 = +62;
				 l_2 = -67; end
		12931: begin l_1 = -62;
				 l_2 = +67; end
		25611: begin l_1 = -62;
				 l_2 = -67; end
		18910: begin l_1 = +62;
				 l_2 = +68; end
		44270: begin l_1 = +62;
				 l_2 = -68; end
		6591: begin l_1 = -62;
				 l_2 = +68; end
		31951: begin l_1 = -62;
				 l_2 = -68; end
		36957: begin l_1 = -63;
				 l_2 = +65; end
		13904: begin l_1 = -63;
				 l_2 = -64; end
		10734: begin l_1 = +63;
				 l_2 = +65; end
		40127: begin l_1 = -63;
				 l_2 = -65; end
		9149: begin l_1 = +63;
				 l_2 = +66; end
		15489: begin l_1 = +63;
				 l_2 = -66; end
		35372: begin l_1 = -63;
				 l_2 = +66; end
		41712: begin l_1 = -63;
				 l_2 = -66; end
		5979: begin l_1 = +63;
				 l_2 = +67; end
		18659: begin l_1 = +63;
				 l_2 = -67; end
		32202: begin l_1 = -63;
				 l_2 = +67; end
		44882: begin l_1 = -63;
				 l_2 = -67; end
		50500: begin l_1 = +63;
				 l_2 = +68; end
		24999: begin l_1 = +63;
				 l_2 = -68; end
		25862: begin l_1 = -63;
				 l_2 = +68; end
		361: begin l_1 = -63;
				 l_2 = -68; end
		23053: begin l_1 = -64;
				 l_2 = +66; end
		27808: begin l_1 = -64;
				 l_2 = -65; end
		21468: begin l_1 = +64;
				 l_2 = +66; end
		29393: begin l_1 = -64;
				 l_2 = -66; end
		18298: begin l_1 = +64;
				 l_2 = +67; end
		30978: begin l_1 = +64;
				 l_2 = -67; end
		19883: begin l_1 = -64;
				 l_2 = +67; end
		32563: begin l_1 = -64;
				 l_2 = -67; end
		11958: begin l_1 = +64;
				 l_2 = +68; end
		37318: begin l_1 = +64;
				 l_2 = -68; end
		13543: begin l_1 = -64;
				 l_2 = +68; end
		38903: begin l_1 = -64;
				 l_2 = -68; end
		46106: begin l_1 = -65;
				 l_2 = +67; end
		4755: begin l_1 = -65;
				 l_2 = -66; end
		42936: begin l_1 = +65;
				 l_2 = +67; end
		7925: begin l_1 = -65;
				 l_2 = -67; end
		36596: begin l_1 = +65;
				 l_2 = +68; end
		11095: begin l_1 = +65;
				 l_2 = -68; end
		39766: begin l_1 = -65;
				 l_2 = +68; end
		14265: begin l_1 = -65;
				 l_2 = -68; end
		41351: begin l_1 = -66;
				 l_2 = +68; end
		9510: begin l_1 = -66;
				 l_2 = -67; end
		35011: begin l_1 = +66;
				 l_2 = +68; end
		15850: begin l_1 = -66;
				 l_2 = -68; end
		31841: begin l_1 = +67;
				 l_2 = +68; end
		19020: begin l_1 = -67;
				 l_2 = -68; end
		default: begin l_1 = 0;
					   l_2 = 0; end
	endcase
end

endmodule

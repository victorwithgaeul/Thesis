// Product (AN) Code DEC_LUT_Decoder
// DEC_LUT_Decoder28bits.v
// Received codeword W = AN + E, E is double AWE (E = e1 + e2), +2^i or -2^i.
module DEC_LUT_Decoder28bits(W, N);
input 	[42:0]	W;
output	[27:0]	N;
parameter A = 17619;

wire 	[27:0]	Q;
wire 	[14:0]	R;
assign Q = W / A;
assign R = W - (A * Q);

reg	signed	[43:0]	Delta;
always@(*) begin
	case(R)
		1: Delta = 44'sb00000000000000000000000000000000000000000001;
		17618: Delta = 44'sb11111111111111111111111111111111111111111111;
		2: Delta = 44'sb00000000000000000000000000000000000000000010;
		17617: Delta = 44'sb11111111111111111111111111111111111111111110;
		4: Delta = 44'sb00000000000000000000000000000000000000000100;
		17615: Delta = 44'sb11111111111111111111111111111111111111111100;
		8: Delta = 44'sb00000000000000000000000000000000000000001000;
		17611: Delta = 44'sb11111111111111111111111111111111111111111000;
		16: Delta = 44'sb00000000000000000000000000000000000000010000;
		17603: Delta = 44'sb11111111111111111111111111111111111111110000;
		32: Delta = 44'sb00000000000000000000000000000000000000100000;
		17587: Delta = 44'sb11111111111111111111111111111111111111100000;
		64: Delta = 44'sb00000000000000000000000000000000000001000000;
		17555: Delta = 44'sb11111111111111111111111111111111111111000000;
		128: Delta = 44'sb00000000000000000000000000000000000010000000;
		17491: Delta = 44'sb11111111111111111111111111111111111110000000;
		256: Delta = 44'sb00000000000000000000000000000000000100000000;
		17363: Delta = 44'sb11111111111111111111111111111111111100000000;
		512: Delta = 44'sb00000000000000000000000000000000001000000000;
		17107: Delta = 44'sb11111111111111111111111111111111111000000000;
		1024: Delta = 44'sb00000000000000000000000000000000010000000000;
		16595: Delta = 44'sb11111111111111111111111111111111110000000000;
		2048: Delta = 44'sb00000000000000000000000000000000100000000000;
		15571: Delta = 44'sb11111111111111111111111111111111100000000000;
		4096: Delta = 44'sb00000000000000000000000000000001000000000000;
		13523: Delta = 44'sb11111111111111111111111111111111000000000000;
		8192: Delta = 44'sb00000000000000000000000000000010000000000000;
		9427: Delta = 44'sb11111111111111111111111111111110000000000000;
		16384: Delta = 44'sb00000000000000000000000000000100000000000000;
		1235: Delta = 44'sb11111111111111111111111111111100000000000000;
		15149: Delta = 44'sb00000000000000000000000000001000000000000000;
		2470: Delta = 44'sb11111111111111111111111111111000000000000000;
		12679: Delta = 44'sb00000000000000000000000000010000000000000000;
		4940: Delta = 44'sb11111111111111111111111111110000000000000000;
		7739: Delta = 44'sb00000000000000000000000000100000000000000000;
		9880: Delta = 44'sb11111111111111111111111111100000000000000000;
		15478: Delta = 44'sb00000000000000000000000001000000000000000000;
		2141: Delta = 44'sb11111111111111111111111111000000000000000000;
		13337: Delta = 44'sb00000000000000000000000010000000000000000000;
		4282: Delta = 44'sb11111111111111111111111110000000000000000000;
		9055: Delta = 44'sb00000000000000000000000100000000000000000000;
		8564: Delta = 44'sb11111111111111111111111100000000000000000000;
		491: Delta = 44'sb00000000000000000000001000000000000000000000;
		17128: Delta = 44'sb11111111111111111111111000000000000000000000;
		982: Delta = 44'sb00000000000000000000010000000000000000000000;
		16637: Delta = 44'sb11111111111111111111110000000000000000000000;
		1964: Delta = 44'sb00000000000000000000100000000000000000000000;
		15655: Delta = 44'sb11111111111111111111100000000000000000000000;
		3928: Delta = 44'sb00000000000000000001000000000000000000000000;
		13691: Delta = 44'sb11111111111111111111000000000000000000000000;
		7856: Delta = 44'sb00000000000000000010000000000000000000000000;
		9763: Delta = 44'sb11111111111111111110000000000000000000000000;
		15712: Delta = 44'sb00000000000000000100000000000000000000000000;
		1907: Delta = 44'sb11111111111111111100000000000000000000000000;
		13805: Delta = 44'sb00000000000000001000000000000000000000000000;
		3814: Delta = 44'sb11111111111111111000000000000000000000000000;
		9991: Delta = 44'sb00000000000000010000000000000000000000000000;
		7628: Delta = 44'sb11111111111111110000000000000000000000000000;
		2363: Delta = 44'sb00000000000000100000000000000000000000000000;
		15256: Delta = 44'sb11111111111111100000000000000000000000000000;
		4726: Delta = 44'sb00000000000001000000000000000000000000000000;
		12893: Delta = 44'sb11111111111111000000000000000000000000000000;
		9452: Delta = 44'sb00000000000010000000000000000000000000000000;
		8167: Delta = 44'sb11111111111110000000000000000000000000000000;
		1285: Delta = 44'sb00000000000100000000000000000000000000000000;
		16334: Delta = 44'sb11111111111100000000000000000000000000000000;
		2570: Delta = 44'sb00000000001000000000000000000000000000000000;
		15049: Delta = 44'sb11111111111000000000000000000000000000000000;
		5140: Delta = 44'sb00000000010000000000000000000000000000000000;
		12479: Delta = 44'sb11111111110000000000000000000000000000000000;
		10280: Delta = 44'sb00000000100000000000000000000000000000000000;
		7339: Delta = 44'sb11111111100000000000000000000000000000000000;
		2941: Delta = 44'sb00000001000000000000000000000000000000000000;
		14678: Delta = 44'sb11111111000000000000000000000000000000000000;
		5882: Delta = 44'sb00000010000000000000000000000000000000000000;
		11737: Delta = 44'sb11111110000000000000000000000000000000000000;
		11764: Delta = 44'sb00000100000000000000000000000000000000000000;
		5855: Delta = 44'sb11111100000000000000000000000000000000000000;
		5909: Delta = 44'sb00001000000000000000000000000000000000000000;
		11710: Delta = 44'sb11111000000000000000000000000000000000000000;
		11818: Delta = 44'sb00010000000000000000000000000000000000000000;
		5801: Delta = 44'sb11110000000000000000000000000000000000000000;
		6017: Delta = 44'sb00100000000000000000000000000000000000000000;
		11602: Delta = 44'sb11100000000000000000000000000000000000000000;
		12034: Delta = 44'sb01000000000000000000000000000000000000000000;
		5585: Delta = 44'sb11000000000000000000000000000000000000000000;
		3: Delta = 44'sb00000000000000000000000000000000000000000011;
		17616: Delta = 44'sb11111111111111111111111111111111111111111101;
		5: Delta = 44'sb00000000000000000000000000000000000000000101;
		17614: Delta = 44'sb11111111111111111111111111111111111111111011;
		9: Delta = 44'sb00000000000000000000000000000000000000001001;
		17612: Delta = 44'sb11111111111111111111111111111111111111111001;
		7: Delta = 44'sb00000000000000000000000000000000000000000111;
		17610: Delta = 44'sb11111111111111111111111111111111111111110111;
		17: Delta = 44'sb00000000000000000000000000000000000000010001;
		17604: Delta = 44'sb11111111111111111111111111111111111111110001;
		15: Delta = 44'sb00000000000000000000000000000000000000001111;
		17602: Delta = 44'sb11111111111111111111111111111111111111101111;
		33: Delta = 44'sb00000000000000000000000000000000000000100001;
		17588: Delta = 44'sb11111111111111111111111111111111111111100001;
		31: Delta = 44'sb00000000000000000000000000000000000000011111;
		17586: Delta = 44'sb11111111111111111111111111111111111111011111;
		65: Delta = 44'sb00000000000000000000000000000000000001000001;
		17556: Delta = 44'sb11111111111111111111111111111111111111000001;
		63: Delta = 44'sb00000000000000000000000000000000000000111111;
		17554: Delta = 44'sb11111111111111111111111111111111111110111111;
		129: Delta = 44'sb00000000000000000000000000000000000010000001;
		17492: Delta = 44'sb11111111111111111111111111111111111110000001;
		127: Delta = 44'sb00000000000000000000000000000000000001111111;
		17490: Delta = 44'sb11111111111111111111111111111111111101111111;
		257: Delta = 44'sb00000000000000000000000000000000000100000001;
		17364: Delta = 44'sb11111111111111111111111111111111111100000001;
		255: Delta = 44'sb00000000000000000000000000000000000011111111;
		17362: Delta = 44'sb11111111111111111111111111111111111011111111;
		513: Delta = 44'sb00000000000000000000000000000000001000000001;
		17108: Delta = 44'sb11111111111111111111111111111111111000000001;
		511: Delta = 44'sb00000000000000000000000000000000000111111111;
		17106: Delta = 44'sb11111111111111111111111111111111110111111111;
		1025: Delta = 44'sb00000000000000000000000000000000010000000001;
		16596: Delta = 44'sb11111111111111111111111111111111110000000001;
		1023: Delta = 44'sb00000000000000000000000000000000001111111111;
		16594: Delta = 44'sb11111111111111111111111111111111101111111111;
		2049: Delta = 44'sb00000000000000000000000000000000100000000001;
		15572: Delta = 44'sb11111111111111111111111111111111100000000001;
		2047: Delta = 44'sb00000000000000000000000000000000011111111111;
		15570: Delta = 44'sb11111111111111111111111111111111011111111111;
		4097: Delta = 44'sb00000000000000000000000000000001000000000001;
		13524: Delta = 44'sb11111111111111111111111111111111000000000001;
		4095: Delta = 44'sb00000000000000000000000000000000111111111111;
		13522: Delta = 44'sb11111111111111111111111111111110111111111111;
		8193: Delta = 44'sb00000000000000000000000000000010000000000001;
		9428: Delta = 44'sb11111111111111111111111111111110000000000001;
		8191: Delta = 44'sb00000000000000000000000000000001111111111111;
		9426: Delta = 44'sb11111111111111111111111111111101111111111111;
		16385: Delta = 44'sb00000000000000000000000000000100000000000001;
		1236: Delta = 44'sb11111111111111111111111111111100000000000001;
		16383: Delta = 44'sb00000000000000000000000000000011111111111111;
		1234: Delta = 44'sb11111111111111111111111111111011111111111111;
		15150: Delta = 44'sb00000000000000000000000000001000000000000001;
		2471: Delta = 44'sb11111111111111111111111111111000000000000001;
		15148: Delta = 44'sb00000000000000000000000000000111111111111111;
		2469: Delta = 44'sb11111111111111111111111111110111111111111111;
		12680: Delta = 44'sb00000000000000000000000000010000000000000001;
		4941: Delta = 44'sb11111111111111111111111111110000000000000001;
		12678: Delta = 44'sb00000000000000000000000000001111111111111111;
		4939: Delta = 44'sb11111111111111111111111111101111111111111111;
		7740: Delta = 44'sb00000000000000000000000000100000000000000001;
		9881: Delta = 44'sb11111111111111111111111111100000000000000001;
		7738: Delta = 44'sb00000000000000000000000000011111111111111111;
		9879: Delta = 44'sb11111111111111111111111111011111111111111111;
		15479: Delta = 44'sb00000000000000000000000001000000000000000001;
		2142: Delta = 44'sb11111111111111111111111111000000000000000001;
		15477: Delta = 44'sb00000000000000000000000000111111111111111111;
		2140: Delta = 44'sb11111111111111111111111110111111111111111111;
		13338: Delta = 44'sb00000000000000000000000010000000000000000001;
		4283: Delta = 44'sb11111111111111111111111110000000000000000001;
		13336: Delta = 44'sb00000000000000000000000001111111111111111111;
		4281: Delta = 44'sb11111111111111111111111101111111111111111111;
		9056: Delta = 44'sb00000000000000000000000100000000000000000001;
		8565: Delta = 44'sb11111111111111111111111100000000000000000001;
		9054: Delta = 44'sb00000000000000000000000011111111111111111111;
		8563: Delta = 44'sb11111111111111111111111011111111111111111111;
		492: Delta = 44'sb00000000000000000000001000000000000000000001;
		17129: Delta = 44'sb11111111111111111111111000000000000000000001;
		490: Delta = 44'sb00000000000000000000000111111111111111111111;
		17127: Delta = 44'sb11111111111111111111110111111111111111111111;
		983: Delta = 44'sb00000000000000000000010000000000000000000001;
		16638: Delta = 44'sb11111111111111111111110000000000000000000001;
		981: Delta = 44'sb00000000000000000000001111111111111111111111;
		16636: Delta = 44'sb11111111111111111111101111111111111111111111;
		1965: Delta = 44'sb00000000000000000000100000000000000000000001;
		15656: Delta = 44'sb11111111111111111111100000000000000000000001;
		1963: Delta = 44'sb00000000000000000000011111111111111111111111;
		15654: Delta = 44'sb11111111111111111111011111111111111111111111;
		3929: Delta = 44'sb00000000000000000001000000000000000000000001;
		13692: Delta = 44'sb11111111111111111111000000000000000000000001;
		3927: Delta = 44'sb00000000000000000000111111111111111111111111;
		13690: Delta = 44'sb11111111111111111110111111111111111111111111;
		7857: Delta = 44'sb00000000000000000010000000000000000000000001;
		9764: Delta = 44'sb11111111111111111110000000000000000000000001;
		7855: Delta = 44'sb00000000000000000001111111111111111111111111;
		9762: Delta = 44'sb11111111111111111101111111111111111111111111;
		15713: Delta = 44'sb00000000000000000100000000000000000000000001;
		1908: Delta = 44'sb11111111111111111100000000000000000000000001;
		15711: Delta = 44'sb00000000000000000011111111111111111111111111;
		1906: Delta = 44'sb11111111111111111011111111111111111111111111;
		13806: Delta = 44'sb00000000000000001000000000000000000000000001;
		3815: Delta = 44'sb11111111111111111000000000000000000000000001;
		13804: Delta = 44'sb00000000000000000111111111111111111111111111;
		3813: Delta = 44'sb11111111111111110111111111111111111111111111;
		9992: Delta = 44'sb00000000000000010000000000000000000000000001;
		7629: Delta = 44'sb11111111111111110000000000000000000000000001;
		9990: Delta = 44'sb00000000000000001111111111111111111111111111;
		7627: Delta = 44'sb11111111111111101111111111111111111111111111;
		2364: Delta = 44'sb00000000000000100000000000000000000000000001;
		15257: Delta = 44'sb11111111111111100000000000000000000000000001;
		2362: Delta = 44'sb00000000000000011111111111111111111111111111;
		15255: Delta = 44'sb11111111111111011111111111111111111111111111;
		4727: Delta = 44'sb00000000000001000000000000000000000000000001;
		12894: Delta = 44'sb11111111111111000000000000000000000000000001;
		4725: Delta = 44'sb00000000000000111111111111111111111111111111;
		12892: Delta = 44'sb11111111111110111111111111111111111111111111;
		9453: Delta = 44'sb00000000000010000000000000000000000000000001;
		8168: Delta = 44'sb11111111111110000000000000000000000000000001;
		9451: Delta = 44'sb00000000000001111111111111111111111111111111;
		8166: Delta = 44'sb11111111111101111111111111111111111111111111;
		1286: Delta = 44'sb00000000000100000000000000000000000000000001;
		16335: Delta = 44'sb11111111111100000000000000000000000000000001;
		1284: Delta = 44'sb00000000000011111111111111111111111111111111;
		16333: Delta = 44'sb11111111111011111111111111111111111111111111;
		2571: Delta = 44'sb00000000001000000000000000000000000000000001;
		15050: Delta = 44'sb11111111111000000000000000000000000000000001;
		2569: Delta = 44'sb00000000000111111111111111111111111111111111;
		15048: Delta = 44'sb11111111110111111111111111111111111111111111;
		5141: Delta = 44'sb00000000010000000000000000000000000000000001;
		12480: Delta = 44'sb11111111110000000000000000000000000000000001;
		5139: Delta = 44'sb00000000001111111111111111111111111111111111;
		12478: Delta = 44'sb11111111101111111111111111111111111111111111;
		10281: Delta = 44'sb00000000100000000000000000000000000000000001;
		7340: Delta = 44'sb11111111100000000000000000000000000000000001;
		10279: Delta = 44'sb00000000011111111111111111111111111111111111;
		7338: Delta = 44'sb11111111011111111111111111111111111111111111;
		2942: Delta = 44'sb00000001000000000000000000000000000000000001;
		14679: Delta = 44'sb11111111000000000000000000000000000000000001;
		2940: Delta = 44'sb00000000111111111111111111111111111111111111;
		14677: Delta = 44'sb11111110111111111111111111111111111111111111;
		5883: Delta = 44'sb00000010000000000000000000000000000000000001;
		11738: Delta = 44'sb11111110000000000000000000000000000000000001;
		5881: Delta = 44'sb00000001111111111111111111111111111111111111;
		11736: Delta = 44'sb11111101111111111111111111111111111111111111;
		11765: Delta = 44'sb00000100000000000000000000000000000000000001;
		5856: Delta = 44'sb11111100000000000000000000000000000000000001;
		11763: Delta = 44'sb00000011111111111111111111111111111111111111;
		5854: Delta = 44'sb11111011111111111111111111111111111111111111;
		5910: Delta = 44'sb00001000000000000000000000000000000000000001;
		11711: Delta = 44'sb11111000000000000000000000000000000000000001;
		5908: Delta = 44'sb00000111111111111111111111111111111111111111;
		11709: Delta = 44'sb11110111111111111111111111111111111111111111;
		11819: Delta = 44'sb00010000000000000000000000000000000000000001;
		5802: Delta = 44'sb11110000000000000000000000000000000000000001;
		11817: Delta = 44'sb00001111111111111111111111111111111111111111;
		5800: Delta = 44'sb11101111111111111111111111111111111111111111;
		6018: Delta = 44'sb00100000000000000000000000000000000000000001;
		11603: Delta = 44'sb11100000000000000000000000000000000000000001;
		6016: Delta = 44'sb00011111111111111111111111111111111111111111;
		11601: Delta = 44'sb11011111111111111111111111111111111111111111;
		12035: Delta = 44'sb01000000000000000000000000000000000000000001;
		5586: Delta = 44'sb11000000000000000000000000000000000000000001;
		12033: Delta = 44'sb00111111111111111111111111111111111111111111;
		5584: Delta = 44'sb10111111111111111111111111111111111111111111;
		6: Delta = 44'sb00000000000000000000000000000000000000000110;
		17613: Delta = 44'sb11111111111111111111111111111111111111111010;
		10: Delta = 44'sb00000000000000000000000000000000000000001010;
		17609: Delta = 44'sb11111111111111111111111111111111111111110110;
		18: Delta = 44'sb00000000000000000000000000000000000000010010;
		17605: Delta = 44'sb11111111111111111111111111111111111111110010;
		14: Delta = 44'sb00000000000000000000000000000000000000001110;
		17601: Delta = 44'sb11111111111111111111111111111111111111101110;
		34: Delta = 44'sb00000000000000000000000000000000000000100010;
		17589: Delta = 44'sb11111111111111111111111111111111111111100010;
		30: Delta = 44'sb00000000000000000000000000000000000000011110;
		17585: Delta = 44'sb11111111111111111111111111111111111111011110;
		66: Delta = 44'sb00000000000000000000000000000000000001000010;
		17557: Delta = 44'sb11111111111111111111111111111111111111000010;
		62: Delta = 44'sb00000000000000000000000000000000000000111110;
		17553: Delta = 44'sb11111111111111111111111111111111111110111110;
		130: Delta = 44'sb00000000000000000000000000000000000010000010;
		17493: Delta = 44'sb11111111111111111111111111111111111110000010;
		126: Delta = 44'sb00000000000000000000000000000000000001111110;
		17489: Delta = 44'sb11111111111111111111111111111111111101111110;
		258: Delta = 44'sb00000000000000000000000000000000000100000010;
		17365: Delta = 44'sb11111111111111111111111111111111111100000010;
		254: Delta = 44'sb00000000000000000000000000000000000011111110;
		17361: Delta = 44'sb11111111111111111111111111111111111011111110;
		514: Delta = 44'sb00000000000000000000000000000000001000000010;
		17109: Delta = 44'sb11111111111111111111111111111111111000000010;
		510: Delta = 44'sb00000000000000000000000000000000000111111110;
		17105: Delta = 44'sb11111111111111111111111111111111110111111110;
		1026: Delta = 44'sb00000000000000000000000000000000010000000010;
		16597: Delta = 44'sb11111111111111111111111111111111110000000010;
		1022: Delta = 44'sb00000000000000000000000000000000001111111110;
		16593: Delta = 44'sb11111111111111111111111111111111101111111110;
		2050: Delta = 44'sb00000000000000000000000000000000100000000010;
		15573: Delta = 44'sb11111111111111111111111111111111100000000010;
		2046: Delta = 44'sb00000000000000000000000000000000011111111110;
		15569: Delta = 44'sb11111111111111111111111111111111011111111110;
		4098: Delta = 44'sb00000000000000000000000000000001000000000010;
		13525: Delta = 44'sb11111111111111111111111111111111000000000010;
		4094: Delta = 44'sb00000000000000000000000000000000111111111110;
		13521: Delta = 44'sb11111111111111111111111111111110111111111110;
		8194: Delta = 44'sb00000000000000000000000000000010000000000010;
		9429: Delta = 44'sb11111111111111111111111111111110000000000010;
		8190: Delta = 44'sb00000000000000000000000000000001111111111110;
		9425: Delta = 44'sb11111111111111111111111111111101111111111110;
		16386: Delta = 44'sb00000000000000000000000000000100000000000010;
		1237: Delta = 44'sb11111111111111111111111111111100000000000010;
		16382: Delta = 44'sb00000000000000000000000000000011111111111110;
		1233: Delta = 44'sb11111111111111111111111111111011111111111110;
		15151: Delta = 44'sb00000000000000000000000000001000000000000010;
		2472: Delta = 44'sb11111111111111111111111111111000000000000010;
		15147: Delta = 44'sb00000000000000000000000000000111111111111110;
		2468: Delta = 44'sb11111111111111111111111111110111111111111110;
		12681: Delta = 44'sb00000000000000000000000000010000000000000010;
		4942: Delta = 44'sb11111111111111111111111111110000000000000010;
		12677: Delta = 44'sb00000000000000000000000000001111111111111110;
		4938: Delta = 44'sb11111111111111111111111111101111111111111110;
		7741: Delta = 44'sb00000000000000000000000000100000000000000010;
		9882: Delta = 44'sb11111111111111111111111111100000000000000010;
		7737: Delta = 44'sb00000000000000000000000000011111111111111110;
		9878: Delta = 44'sb11111111111111111111111111011111111111111110;
		15480: Delta = 44'sb00000000000000000000000001000000000000000010;
		2143: Delta = 44'sb11111111111111111111111111000000000000000010;
		15476: Delta = 44'sb00000000000000000000000000111111111111111110;
		2139: Delta = 44'sb11111111111111111111111110111111111111111110;
		13339: Delta = 44'sb00000000000000000000000010000000000000000010;
		4284: Delta = 44'sb11111111111111111111111110000000000000000010;
		13335: Delta = 44'sb00000000000000000000000001111111111111111110;
		4280: Delta = 44'sb11111111111111111111111101111111111111111110;
		9057: Delta = 44'sb00000000000000000000000100000000000000000010;
		8566: Delta = 44'sb11111111111111111111111100000000000000000010;
		9053: Delta = 44'sb00000000000000000000000011111111111111111110;
		8562: Delta = 44'sb11111111111111111111111011111111111111111110;
		493: Delta = 44'sb00000000000000000000001000000000000000000010;
		17130: Delta = 44'sb11111111111111111111111000000000000000000010;
		489: Delta = 44'sb00000000000000000000000111111111111111111110;
		17126: Delta = 44'sb11111111111111111111110111111111111111111110;
		984: Delta = 44'sb00000000000000000000010000000000000000000010;
		16639: Delta = 44'sb11111111111111111111110000000000000000000010;
		980: Delta = 44'sb00000000000000000000001111111111111111111110;
		16635: Delta = 44'sb11111111111111111111101111111111111111111110;
		1966: Delta = 44'sb00000000000000000000100000000000000000000010;
		15657: Delta = 44'sb11111111111111111111100000000000000000000010;
		1962: Delta = 44'sb00000000000000000000011111111111111111111110;
		15653: Delta = 44'sb11111111111111111111011111111111111111111110;
		3930: Delta = 44'sb00000000000000000001000000000000000000000010;
		13693: Delta = 44'sb11111111111111111111000000000000000000000010;
		3926: Delta = 44'sb00000000000000000000111111111111111111111110;
		13689: Delta = 44'sb11111111111111111110111111111111111111111110;
		7858: Delta = 44'sb00000000000000000010000000000000000000000010;
		9765: Delta = 44'sb11111111111111111110000000000000000000000010;
		7854: Delta = 44'sb00000000000000000001111111111111111111111110;
		9761: Delta = 44'sb11111111111111111101111111111111111111111110;
		15714: Delta = 44'sb00000000000000000100000000000000000000000010;
		1909: Delta = 44'sb11111111111111111100000000000000000000000010;
		15710: Delta = 44'sb00000000000000000011111111111111111111111110;
		1905: Delta = 44'sb11111111111111111011111111111111111111111110;
		13807: Delta = 44'sb00000000000000001000000000000000000000000010;
		3816: Delta = 44'sb11111111111111111000000000000000000000000010;
		13803: Delta = 44'sb00000000000000000111111111111111111111111110;
		3812: Delta = 44'sb11111111111111110111111111111111111111111110;
		9993: Delta = 44'sb00000000000000010000000000000000000000000010;
		7630: Delta = 44'sb11111111111111110000000000000000000000000010;
		9989: Delta = 44'sb00000000000000001111111111111111111111111110;
		7626: Delta = 44'sb11111111111111101111111111111111111111111110;
		2365: Delta = 44'sb00000000000000100000000000000000000000000010;
		15258: Delta = 44'sb11111111111111100000000000000000000000000010;
		2361: Delta = 44'sb00000000000000011111111111111111111111111110;
		15254: Delta = 44'sb11111111111111011111111111111111111111111110;
		4728: Delta = 44'sb00000000000001000000000000000000000000000010;
		12895: Delta = 44'sb11111111111111000000000000000000000000000010;
		4724: Delta = 44'sb00000000000000111111111111111111111111111110;
		12891: Delta = 44'sb11111111111110111111111111111111111111111110;
		9454: Delta = 44'sb00000000000010000000000000000000000000000010;
		8169: Delta = 44'sb11111111111110000000000000000000000000000010;
		9450: Delta = 44'sb00000000000001111111111111111111111111111110;
		8165: Delta = 44'sb11111111111101111111111111111111111111111110;
		1287: Delta = 44'sb00000000000100000000000000000000000000000010;
		16336: Delta = 44'sb11111111111100000000000000000000000000000010;
		1283: Delta = 44'sb00000000000011111111111111111111111111111110;
		16332: Delta = 44'sb11111111111011111111111111111111111111111110;
		2572: Delta = 44'sb00000000001000000000000000000000000000000010;
		15051: Delta = 44'sb11111111111000000000000000000000000000000010;
		2568: Delta = 44'sb00000000000111111111111111111111111111111110;
		15047: Delta = 44'sb11111111110111111111111111111111111111111110;
		5142: Delta = 44'sb00000000010000000000000000000000000000000010;
		12481: Delta = 44'sb11111111110000000000000000000000000000000010;
		5138: Delta = 44'sb00000000001111111111111111111111111111111110;
		12477: Delta = 44'sb11111111101111111111111111111111111111111110;
		10282: Delta = 44'sb00000000100000000000000000000000000000000010;
		7341: Delta = 44'sb11111111100000000000000000000000000000000010;
		10278: Delta = 44'sb00000000011111111111111111111111111111111110;
		7337: Delta = 44'sb11111111011111111111111111111111111111111110;
		2943: Delta = 44'sb00000001000000000000000000000000000000000010;
		14680: Delta = 44'sb11111111000000000000000000000000000000000010;
		2939: Delta = 44'sb00000000111111111111111111111111111111111110;
		14676: Delta = 44'sb11111110111111111111111111111111111111111110;
		5884: Delta = 44'sb00000010000000000000000000000000000000000010;
		11739: Delta = 44'sb11111110000000000000000000000000000000000010;
		5880: Delta = 44'sb00000001111111111111111111111111111111111110;
		11735: Delta = 44'sb11111101111111111111111111111111111111111110;
		11766: Delta = 44'sb00000100000000000000000000000000000000000010;
		5857: Delta = 44'sb11111100000000000000000000000000000000000010;
		11762: Delta = 44'sb00000011111111111111111111111111111111111110;
		5853: Delta = 44'sb11111011111111111111111111111111111111111110;
		5911: Delta = 44'sb00001000000000000000000000000000000000000010;
		11712: Delta = 44'sb11111000000000000000000000000000000000000010;
		5907: Delta = 44'sb00000111111111111111111111111111111111111110;
		11708: Delta = 44'sb11110111111111111111111111111111111111111110;
		11820: Delta = 44'sb00010000000000000000000000000000000000000010;
		5803: Delta = 44'sb11110000000000000000000000000000000000000010;
		11816: Delta = 44'sb00001111111111111111111111111111111111111110;
		5799: Delta = 44'sb11101111111111111111111111111111111111111110;
		6019: Delta = 44'sb00100000000000000000000000000000000000000010;
		11604: Delta = 44'sb11100000000000000000000000000000000000000010;
		6015: Delta = 44'sb00011111111111111111111111111111111111111110;
		11600: Delta = 44'sb11011111111111111111111111111111111111111110;
		12036: Delta = 44'sb01000000000000000000000000000000000000000010;
		5587: Delta = 44'sb11000000000000000000000000000000000000000010;
		12032: Delta = 44'sb00111111111111111111111111111111111111111110;
		5583: Delta = 44'sb10111111111111111111111111111111111111111110;
		12: Delta = 44'sb00000000000000000000000000000000000000001100;
		17607: Delta = 44'sb11111111111111111111111111111111111111110100;
		20: Delta = 44'sb00000000000000000000000000000000000000010100;
		17599: Delta = 44'sb11111111111111111111111111111111111111101100;
		36: Delta = 44'sb00000000000000000000000000000000000000100100;
		17591: Delta = 44'sb11111111111111111111111111111111111111100100;
		28: Delta = 44'sb00000000000000000000000000000000000000011100;
		17583: Delta = 44'sb11111111111111111111111111111111111111011100;
		68: Delta = 44'sb00000000000000000000000000000000000001000100;
		17559: Delta = 44'sb11111111111111111111111111111111111111000100;
		60: Delta = 44'sb00000000000000000000000000000000000000111100;
		17551: Delta = 44'sb11111111111111111111111111111111111110111100;
		132: Delta = 44'sb00000000000000000000000000000000000010000100;
		17495: Delta = 44'sb11111111111111111111111111111111111110000100;
		124: Delta = 44'sb00000000000000000000000000000000000001111100;
		17487: Delta = 44'sb11111111111111111111111111111111111101111100;
		260: Delta = 44'sb00000000000000000000000000000000000100000100;
		17367: Delta = 44'sb11111111111111111111111111111111111100000100;
		252: Delta = 44'sb00000000000000000000000000000000000011111100;
		17359: Delta = 44'sb11111111111111111111111111111111111011111100;
		516: Delta = 44'sb00000000000000000000000000000000001000000100;
		17111: Delta = 44'sb11111111111111111111111111111111111000000100;
		508: Delta = 44'sb00000000000000000000000000000000000111111100;
		17103: Delta = 44'sb11111111111111111111111111111111110111111100;
		1028: Delta = 44'sb00000000000000000000000000000000010000000100;
		16599: Delta = 44'sb11111111111111111111111111111111110000000100;
		1020: Delta = 44'sb00000000000000000000000000000000001111111100;
		16591: Delta = 44'sb11111111111111111111111111111111101111111100;
		2052: Delta = 44'sb00000000000000000000000000000000100000000100;
		15575: Delta = 44'sb11111111111111111111111111111111100000000100;
		2044: Delta = 44'sb00000000000000000000000000000000011111111100;
		15567: Delta = 44'sb11111111111111111111111111111111011111111100;
		4100: Delta = 44'sb00000000000000000000000000000001000000000100;
		13527: Delta = 44'sb11111111111111111111111111111111000000000100;
		4092: Delta = 44'sb00000000000000000000000000000000111111111100;
		13519: Delta = 44'sb11111111111111111111111111111110111111111100;
		8196: Delta = 44'sb00000000000000000000000000000010000000000100;
		9431: Delta = 44'sb11111111111111111111111111111110000000000100;
		8188: Delta = 44'sb00000000000000000000000000000001111111111100;
		9423: Delta = 44'sb11111111111111111111111111111101111111111100;
		16388: Delta = 44'sb00000000000000000000000000000100000000000100;
		1239: Delta = 44'sb11111111111111111111111111111100000000000100;
		16380: Delta = 44'sb00000000000000000000000000000011111111111100;
		1231: Delta = 44'sb11111111111111111111111111111011111111111100;
		15153: Delta = 44'sb00000000000000000000000000001000000000000100;
		2474: Delta = 44'sb11111111111111111111111111111000000000000100;
		15145: Delta = 44'sb00000000000000000000000000000111111111111100;
		2466: Delta = 44'sb11111111111111111111111111110111111111111100;
		12683: Delta = 44'sb00000000000000000000000000010000000000000100;
		4944: Delta = 44'sb11111111111111111111111111110000000000000100;
		12675: Delta = 44'sb00000000000000000000000000001111111111111100;
		4936: Delta = 44'sb11111111111111111111111111101111111111111100;
		7743: Delta = 44'sb00000000000000000000000000100000000000000100;
		9884: Delta = 44'sb11111111111111111111111111100000000000000100;
		7735: Delta = 44'sb00000000000000000000000000011111111111111100;
		9876: Delta = 44'sb11111111111111111111111111011111111111111100;
		15482: Delta = 44'sb00000000000000000000000001000000000000000100;
		2145: Delta = 44'sb11111111111111111111111111000000000000000100;
		15474: Delta = 44'sb00000000000000000000000000111111111111111100;
		2137: Delta = 44'sb11111111111111111111111110111111111111111100;
		13341: Delta = 44'sb00000000000000000000000010000000000000000100;
		4286: Delta = 44'sb11111111111111111111111110000000000000000100;
		13333: Delta = 44'sb00000000000000000000000001111111111111111100;
		4278: Delta = 44'sb11111111111111111111111101111111111111111100;
		9059: Delta = 44'sb00000000000000000000000100000000000000000100;
		8568: Delta = 44'sb11111111111111111111111100000000000000000100;
		9051: Delta = 44'sb00000000000000000000000011111111111111111100;
		8560: Delta = 44'sb11111111111111111111111011111111111111111100;
		495: Delta = 44'sb00000000000000000000001000000000000000000100;
		17132: Delta = 44'sb11111111111111111111111000000000000000000100;
		487: Delta = 44'sb00000000000000000000000111111111111111111100;
		17124: Delta = 44'sb11111111111111111111110111111111111111111100;
		986: Delta = 44'sb00000000000000000000010000000000000000000100;
		16641: Delta = 44'sb11111111111111111111110000000000000000000100;
		978: Delta = 44'sb00000000000000000000001111111111111111111100;
		16633: Delta = 44'sb11111111111111111111101111111111111111111100;
		1968: Delta = 44'sb00000000000000000000100000000000000000000100;
		15659: Delta = 44'sb11111111111111111111100000000000000000000100;
		1960: Delta = 44'sb00000000000000000000011111111111111111111100;
		15651: Delta = 44'sb11111111111111111111011111111111111111111100;
		3932: Delta = 44'sb00000000000000000001000000000000000000000100;
		13695: Delta = 44'sb11111111111111111111000000000000000000000100;
		3924: Delta = 44'sb00000000000000000000111111111111111111111100;
		13687: Delta = 44'sb11111111111111111110111111111111111111111100;
		7860: Delta = 44'sb00000000000000000010000000000000000000000100;
		9767: Delta = 44'sb11111111111111111110000000000000000000000100;
		7852: Delta = 44'sb00000000000000000001111111111111111111111100;
		9759: Delta = 44'sb11111111111111111101111111111111111111111100;
		15716: Delta = 44'sb00000000000000000100000000000000000000000100;
		1911: Delta = 44'sb11111111111111111100000000000000000000000100;
		15708: Delta = 44'sb00000000000000000011111111111111111111111100;
		1903: Delta = 44'sb11111111111111111011111111111111111111111100;
		13809: Delta = 44'sb00000000000000001000000000000000000000000100;
		3818: Delta = 44'sb11111111111111111000000000000000000000000100;
		13801: Delta = 44'sb00000000000000000111111111111111111111111100;
		3810: Delta = 44'sb11111111111111110111111111111111111111111100;
		9995: Delta = 44'sb00000000000000010000000000000000000000000100;
		7632: Delta = 44'sb11111111111111110000000000000000000000000100;
		9987: Delta = 44'sb00000000000000001111111111111111111111111100;
		7624: Delta = 44'sb11111111111111101111111111111111111111111100;
		2367: Delta = 44'sb00000000000000100000000000000000000000000100;
		15260: Delta = 44'sb11111111111111100000000000000000000000000100;
		2359: Delta = 44'sb00000000000000011111111111111111111111111100;
		15252: Delta = 44'sb11111111111111011111111111111111111111111100;
		4730: Delta = 44'sb00000000000001000000000000000000000000000100;
		12897: Delta = 44'sb11111111111111000000000000000000000000000100;
		4722: Delta = 44'sb00000000000000111111111111111111111111111100;
		12889: Delta = 44'sb11111111111110111111111111111111111111111100;
		9456: Delta = 44'sb00000000000010000000000000000000000000000100;
		8171: Delta = 44'sb11111111111110000000000000000000000000000100;
		9448: Delta = 44'sb00000000000001111111111111111111111111111100;
		8163: Delta = 44'sb11111111111101111111111111111111111111111100;
		1289: Delta = 44'sb00000000000100000000000000000000000000000100;
		16338: Delta = 44'sb11111111111100000000000000000000000000000100;
		1281: Delta = 44'sb00000000000011111111111111111111111111111100;
		16330: Delta = 44'sb11111111111011111111111111111111111111111100;
		2574: Delta = 44'sb00000000001000000000000000000000000000000100;
		15053: Delta = 44'sb11111111111000000000000000000000000000000100;
		2566: Delta = 44'sb00000000000111111111111111111111111111111100;
		15045: Delta = 44'sb11111111110111111111111111111111111111111100;
		5144: Delta = 44'sb00000000010000000000000000000000000000000100;
		12483: Delta = 44'sb11111111110000000000000000000000000000000100;
		5136: Delta = 44'sb00000000001111111111111111111111111111111100;
		12475: Delta = 44'sb11111111101111111111111111111111111111111100;
		10284: Delta = 44'sb00000000100000000000000000000000000000000100;
		7343: Delta = 44'sb11111111100000000000000000000000000000000100;
		10276: Delta = 44'sb00000000011111111111111111111111111111111100;
		7335: Delta = 44'sb11111111011111111111111111111111111111111100;
		2945: Delta = 44'sb00000001000000000000000000000000000000000100;
		14682: Delta = 44'sb11111111000000000000000000000000000000000100;
		2937: Delta = 44'sb00000000111111111111111111111111111111111100;
		14674: Delta = 44'sb11111110111111111111111111111111111111111100;
		5886: Delta = 44'sb00000010000000000000000000000000000000000100;
		11741: Delta = 44'sb11111110000000000000000000000000000000000100;
		5878: Delta = 44'sb00000001111111111111111111111111111111111100;
		11733: Delta = 44'sb11111101111111111111111111111111111111111100;
		11768: Delta = 44'sb00000100000000000000000000000000000000000100;
		5859: Delta = 44'sb11111100000000000000000000000000000000000100;
		11760: Delta = 44'sb00000011111111111111111111111111111111111100;
		5851: Delta = 44'sb11111011111111111111111111111111111111111100;
		5913: Delta = 44'sb00001000000000000000000000000000000000000100;
		11714: Delta = 44'sb11111000000000000000000000000000000000000100;
		5905: Delta = 44'sb00000111111111111111111111111111111111111100;
		11706: Delta = 44'sb11110111111111111111111111111111111111111100;
		11822: Delta = 44'sb00010000000000000000000000000000000000000100;
		5805: Delta = 44'sb11110000000000000000000000000000000000000100;
		11814: Delta = 44'sb00001111111111111111111111111111111111111100;
		5797: Delta = 44'sb11101111111111111111111111111111111111111100;
		6021: Delta = 44'sb00100000000000000000000000000000000000000100;
		11606: Delta = 44'sb11100000000000000000000000000000000000000100;
		6013: Delta = 44'sb00011111111111111111111111111111111111111100;
		11598: Delta = 44'sb11011111111111111111111111111111111111111100;
		12038: Delta = 44'sb01000000000000000000000000000000000000000100;
		5589: Delta = 44'sb11000000000000000000000000000000000000000100;
		12030: Delta = 44'sb00111111111111111111111111111111111111111100;
		5581: Delta = 44'sb10111111111111111111111111111111111111111100;
		24: Delta = 44'sb00000000000000000000000000000000000000011000;
		17595: Delta = 44'sb11111111111111111111111111111111111111101000;
		40: Delta = 44'sb00000000000000000000000000000000000000101000;
		17579: Delta = 44'sb11111111111111111111111111111111111111011000;
		72: Delta = 44'sb00000000000000000000000000000000000001001000;
		17563: Delta = 44'sb11111111111111111111111111111111111111001000;
		56: Delta = 44'sb00000000000000000000000000000000000000111000;
		17547: Delta = 44'sb11111111111111111111111111111111111110111000;
		136: Delta = 44'sb00000000000000000000000000000000000010001000;
		17499: Delta = 44'sb11111111111111111111111111111111111110001000;
		120: Delta = 44'sb00000000000000000000000000000000000001111000;
		17483: Delta = 44'sb11111111111111111111111111111111111101111000;
		264: Delta = 44'sb00000000000000000000000000000000000100001000;
		17371: Delta = 44'sb11111111111111111111111111111111111100001000;
		248: Delta = 44'sb00000000000000000000000000000000000011111000;
		17355: Delta = 44'sb11111111111111111111111111111111111011111000;
		520: Delta = 44'sb00000000000000000000000000000000001000001000;
		17115: Delta = 44'sb11111111111111111111111111111111111000001000;
		504: Delta = 44'sb00000000000000000000000000000000000111111000;
		17099: Delta = 44'sb11111111111111111111111111111111110111111000;
		1032: Delta = 44'sb00000000000000000000000000000000010000001000;
		16603: Delta = 44'sb11111111111111111111111111111111110000001000;
		1016: Delta = 44'sb00000000000000000000000000000000001111111000;
		16587: Delta = 44'sb11111111111111111111111111111111101111111000;
		2056: Delta = 44'sb00000000000000000000000000000000100000001000;
		15579: Delta = 44'sb11111111111111111111111111111111100000001000;
		2040: Delta = 44'sb00000000000000000000000000000000011111111000;
		15563: Delta = 44'sb11111111111111111111111111111111011111111000;
		4104: Delta = 44'sb00000000000000000000000000000001000000001000;
		13531: Delta = 44'sb11111111111111111111111111111111000000001000;
		4088: Delta = 44'sb00000000000000000000000000000000111111111000;
		13515: Delta = 44'sb11111111111111111111111111111110111111111000;
		8200: Delta = 44'sb00000000000000000000000000000010000000001000;
		9435: Delta = 44'sb11111111111111111111111111111110000000001000;
		8184: Delta = 44'sb00000000000000000000000000000001111111111000;
		9419: Delta = 44'sb11111111111111111111111111111101111111111000;
		16392: Delta = 44'sb00000000000000000000000000000100000000001000;
		1243: Delta = 44'sb11111111111111111111111111111100000000001000;
		16376: Delta = 44'sb00000000000000000000000000000011111111111000;
		1227: Delta = 44'sb11111111111111111111111111111011111111111000;
		15157: Delta = 44'sb00000000000000000000000000001000000000001000;
		2478: Delta = 44'sb11111111111111111111111111111000000000001000;
		15141: Delta = 44'sb00000000000000000000000000000111111111111000;
		2462: Delta = 44'sb11111111111111111111111111110111111111111000;
		12687: Delta = 44'sb00000000000000000000000000010000000000001000;
		4948: Delta = 44'sb11111111111111111111111111110000000000001000;
		12671: Delta = 44'sb00000000000000000000000000001111111111111000;
		4932: Delta = 44'sb11111111111111111111111111101111111111111000;
		7747: Delta = 44'sb00000000000000000000000000100000000000001000;
		9888: Delta = 44'sb11111111111111111111111111100000000000001000;
		7731: Delta = 44'sb00000000000000000000000000011111111111111000;
		9872: Delta = 44'sb11111111111111111111111111011111111111111000;
		15486: Delta = 44'sb00000000000000000000000001000000000000001000;
		2149: Delta = 44'sb11111111111111111111111111000000000000001000;
		15470: Delta = 44'sb00000000000000000000000000111111111111111000;
		2133: Delta = 44'sb11111111111111111111111110111111111111111000;
		13345: Delta = 44'sb00000000000000000000000010000000000000001000;
		4290: Delta = 44'sb11111111111111111111111110000000000000001000;
		13329: Delta = 44'sb00000000000000000000000001111111111111111000;
		4274: Delta = 44'sb11111111111111111111111101111111111111111000;
		9063: Delta = 44'sb00000000000000000000000100000000000000001000;
		8572: Delta = 44'sb11111111111111111111111100000000000000001000;
		9047: Delta = 44'sb00000000000000000000000011111111111111111000;
		8556: Delta = 44'sb11111111111111111111111011111111111111111000;
		499: Delta = 44'sb00000000000000000000001000000000000000001000;
		17136: Delta = 44'sb11111111111111111111111000000000000000001000;
		483: Delta = 44'sb00000000000000000000000111111111111111111000;
		17120: Delta = 44'sb11111111111111111111110111111111111111111000;
		990: Delta = 44'sb00000000000000000000010000000000000000001000;
		16645: Delta = 44'sb11111111111111111111110000000000000000001000;
		974: Delta = 44'sb00000000000000000000001111111111111111111000;
		16629: Delta = 44'sb11111111111111111111101111111111111111111000;
		1972: Delta = 44'sb00000000000000000000100000000000000000001000;
		15663: Delta = 44'sb11111111111111111111100000000000000000001000;
		1956: Delta = 44'sb00000000000000000000011111111111111111111000;
		15647: Delta = 44'sb11111111111111111111011111111111111111111000;
		3936: Delta = 44'sb00000000000000000001000000000000000000001000;
		13699: Delta = 44'sb11111111111111111111000000000000000000001000;
		3920: Delta = 44'sb00000000000000000000111111111111111111111000;
		13683: Delta = 44'sb11111111111111111110111111111111111111111000;
		7864: Delta = 44'sb00000000000000000010000000000000000000001000;
		9771: Delta = 44'sb11111111111111111110000000000000000000001000;
		7848: Delta = 44'sb00000000000000000001111111111111111111111000;
		9755: Delta = 44'sb11111111111111111101111111111111111111111000;
		15720: Delta = 44'sb00000000000000000100000000000000000000001000;
		1915: Delta = 44'sb11111111111111111100000000000000000000001000;
		15704: Delta = 44'sb00000000000000000011111111111111111111111000;
		1899: Delta = 44'sb11111111111111111011111111111111111111111000;
		13813: Delta = 44'sb00000000000000001000000000000000000000001000;
		3822: Delta = 44'sb11111111111111111000000000000000000000001000;
		13797: Delta = 44'sb00000000000000000111111111111111111111111000;
		3806: Delta = 44'sb11111111111111110111111111111111111111111000;
		9999: Delta = 44'sb00000000000000010000000000000000000000001000;
		7636: Delta = 44'sb11111111111111110000000000000000000000001000;
		9983: Delta = 44'sb00000000000000001111111111111111111111111000;
		7620: Delta = 44'sb11111111111111101111111111111111111111111000;
		2371: Delta = 44'sb00000000000000100000000000000000000000001000;
		15264: Delta = 44'sb11111111111111100000000000000000000000001000;
		2355: Delta = 44'sb00000000000000011111111111111111111111111000;
		15248: Delta = 44'sb11111111111111011111111111111111111111111000;
		4734: Delta = 44'sb00000000000001000000000000000000000000001000;
		12901: Delta = 44'sb11111111111111000000000000000000000000001000;
		4718: Delta = 44'sb00000000000000111111111111111111111111111000;
		12885: Delta = 44'sb11111111111110111111111111111111111111111000;
		9460: Delta = 44'sb00000000000010000000000000000000000000001000;
		8175: Delta = 44'sb11111111111110000000000000000000000000001000;
		9444: Delta = 44'sb00000000000001111111111111111111111111111000;
		8159: Delta = 44'sb11111111111101111111111111111111111111111000;
		1293: Delta = 44'sb00000000000100000000000000000000000000001000;
		16342: Delta = 44'sb11111111111100000000000000000000000000001000;
		1277: Delta = 44'sb00000000000011111111111111111111111111111000;
		16326: Delta = 44'sb11111111111011111111111111111111111111111000;
		2578: Delta = 44'sb00000000001000000000000000000000000000001000;
		15057: Delta = 44'sb11111111111000000000000000000000000000001000;
		2562: Delta = 44'sb00000000000111111111111111111111111111111000;
		15041: Delta = 44'sb11111111110111111111111111111111111111111000;
		5148: Delta = 44'sb00000000010000000000000000000000000000001000;
		12487: Delta = 44'sb11111111110000000000000000000000000000001000;
		5132: Delta = 44'sb00000000001111111111111111111111111111111000;
		12471: Delta = 44'sb11111111101111111111111111111111111111111000;
		10288: Delta = 44'sb00000000100000000000000000000000000000001000;
		7347: Delta = 44'sb11111111100000000000000000000000000000001000;
		10272: Delta = 44'sb00000000011111111111111111111111111111111000;
		7331: Delta = 44'sb11111111011111111111111111111111111111111000;
		2949: Delta = 44'sb00000001000000000000000000000000000000001000;
		14686: Delta = 44'sb11111111000000000000000000000000000000001000;
		2933: Delta = 44'sb00000000111111111111111111111111111111111000;
		14670: Delta = 44'sb11111110111111111111111111111111111111111000;
		5890: Delta = 44'sb00000010000000000000000000000000000000001000;
		11745: Delta = 44'sb11111110000000000000000000000000000000001000;
		5874: Delta = 44'sb00000001111111111111111111111111111111111000;
		11729: Delta = 44'sb11111101111111111111111111111111111111111000;
		11772: Delta = 44'sb00000100000000000000000000000000000000001000;
		5863: Delta = 44'sb11111100000000000000000000000000000000001000;
		11756: Delta = 44'sb00000011111111111111111111111111111111111000;
		5847: Delta = 44'sb11111011111111111111111111111111111111111000;
		5917: Delta = 44'sb00001000000000000000000000000000000000001000;
		11718: Delta = 44'sb11111000000000000000000000000000000000001000;
		5901: Delta = 44'sb00000111111111111111111111111111111111111000;
		11702: Delta = 44'sb11110111111111111111111111111111111111111000;
		11826: Delta = 44'sb00010000000000000000000000000000000000001000;
		5809: Delta = 44'sb11110000000000000000000000000000000000001000;
		11810: Delta = 44'sb00001111111111111111111111111111111111111000;
		5793: Delta = 44'sb11101111111111111111111111111111111111111000;
		6025: Delta = 44'sb00100000000000000000000000000000000000001000;
		11610: Delta = 44'sb11100000000000000000000000000000000000001000;
		6009: Delta = 44'sb00011111111111111111111111111111111111111000;
		11594: Delta = 44'sb11011111111111111111111111111111111111111000;
		12042: Delta = 44'sb01000000000000000000000000000000000000001000;
		5593: Delta = 44'sb11000000000000000000000000000000000000001000;
		12026: Delta = 44'sb00111111111111111111111111111111111111111000;
		5577: Delta = 44'sb10111111111111111111111111111111111111111000;
		48: Delta = 44'sb00000000000000000000000000000000000000110000;
		17571: Delta = 44'sb11111111111111111111111111111111111111010000;
		80: Delta = 44'sb00000000000000000000000000000000000001010000;
		17539: Delta = 44'sb11111111111111111111111111111111111110110000;
		144: Delta = 44'sb00000000000000000000000000000000000010010000;
		17507: Delta = 44'sb11111111111111111111111111111111111110010000;
		112: Delta = 44'sb00000000000000000000000000000000000001110000;
		17475: Delta = 44'sb11111111111111111111111111111111111101110000;
		272: Delta = 44'sb00000000000000000000000000000000000100010000;
		17379: Delta = 44'sb11111111111111111111111111111111111100010000;
		240: Delta = 44'sb00000000000000000000000000000000000011110000;
		17347: Delta = 44'sb11111111111111111111111111111111111011110000;
		528: Delta = 44'sb00000000000000000000000000000000001000010000;
		17123: Delta = 44'sb11111111111111111111111111111111111000010000;
		496: Delta = 44'sb00000000000000000000000000000000000111110000;
		17091: Delta = 44'sb11111111111111111111111111111111110111110000;
		1040: Delta = 44'sb00000000000000000000000000000000010000010000;
		16611: Delta = 44'sb11111111111111111111111111111111110000010000;
		1008: Delta = 44'sb00000000000000000000000000000000001111110000;
		16579: Delta = 44'sb11111111111111111111111111111111101111110000;
		2064: Delta = 44'sb00000000000000000000000000000000100000010000;
		15587: Delta = 44'sb11111111111111111111111111111111100000010000;
		2032: Delta = 44'sb00000000000000000000000000000000011111110000;
		15555: Delta = 44'sb11111111111111111111111111111111011111110000;
		4112: Delta = 44'sb00000000000000000000000000000001000000010000;
		13539: Delta = 44'sb11111111111111111111111111111111000000010000;
		4080: Delta = 44'sb00000000000000000000000000000000111111110000;
		13507: Delta = 44'sb11111111111111111111111111111110111111110000;
		8208: Delta = 44'sb00000000000000000000000000000010000000010000;
		9443: Delta = 44'sb11111111111111111111111111111110000000010000;
		8176: Delta = 44'sb00000000000000000000000000000001111111110000;
		9411: Delta = 44'sb11111111111111111111111111111101111111110000;
		16400: Delta = 44'sb00000000000000000000000000000100000000010000;
		1251: Delta = 44'sb11111111111111111111111111111100000000010000;
		16368: Delta = 44'sb00000000000000000000000000000011111111110000;
		1219: Delta = 44'sb11111111111111111111111111111011111111110000;
		15165: Delta = 44'sb00000000000000000000000000001000000000010000;
		2486: Delta = 44'sb11111111111111111111111111111000000000010000;
		15133: Delta = 44'sb00000000000000000000000000000111111111110000;
		2454: Delta = 44'sb11111111111111111111111111110111111111110000;
		12695: Delta = 44'sb00000000000000000000000000010000000000010000;
		4956: Delta = 44'sb11111111111111111111111111110000000000010000;
		12663: Delta = 44'sb00000000000000000000000000001111111111110000;
		4924: Delta = 44'sb11111111111111111111111111101111111111110000;
		7755: Delta = 44'sb00000000000000000000000000100000000000010000;
		9896: Delta = 44'sb11111111111111111111111111100000000000010000;
		7723: Delta = 44'sb00000000000000000000000000011111111111110000;
		9864: Delta = 44'sb11111111111111111111111111011111111111110000;
		15494: Delta = 44'sb00000000000000000000000001000000000000010000;
		2157: Delta = 44'sb11111111111111111111111111000000000000010000;
		15462: Delta = 44'sb00000000000000000000000000111111111111110000;
		2125: Delta = 44'sb11111111111111111111111110111111111111110000;
		13353: Delta = 44'sb00000000000000000000000010000000000000010000;
		4298: Delta = 44'sb11111111111111111111111110000000000000010000;
		13321: Delta = 44'sb00000000000000000000000001111111111111110000;
		4266: Delta = 44'sb11111111111111111111111101111111111111110000;
		9071: Delta = 44'sb00000000000000000000000100000000000000010000;
		8580: Delta = 44'sb11111111111111111111111100000000000000010000;
		9039: Delta = 44'sb00000000000000000000000011111111111111110000;
		8548: Delta = 44'sb11111111111111111111111011111111111111110000;
		507: Delta = 44'sb00000000000000000000001000000000000000010000;
		17144: Delta = 44'sb11111111111111111111111000000000000000010000;
		475: Delta = 44'sb00000000000000000000000111111111111111110000;
		17112: Delta = 44'sb11111111111111111111110111111111111111110000;
		998: Delta = 44'sb00000000000000000000010000000000000000010000;
		16653: Delta = 44'sb11111111111111111111110000000000000000010000;
		966: Delta = 44'sb00000000000000000000001111111111111111110000;
		16621: Delta = 44'sb11111111111111111111101111111111111111110000;
		1980: Delta = 44'sb00000000000000000000100000000000000000010000;
		15671: Delta = 44'sb11111111111111111111100000000000000000010000;
		1948: Delta = 44'sb00000000000000000000011111111111111111110000;
		15639: Delta = 44'sb11111111111111111111011111111111111111110000;
		3944: Delta = 44'sb00000000000000000001000000000000000000010000;
		13707: Delta = 44'sb11111111111111111111000000000000000000010000;
		3912: Delta = 44'sb00000000000000000000111111111111111111110000;
		13675: Delta = 44'sb11111111111111111110111111111111111111110000;
		7872: Delta = 44'sb00000000000000000010000000000000000000010000;
		9779: Delta = 44'sb11111111111111111110000000000000000000010000;
		7840: Delta = 44'sb00000000000000000001111111111111111111110000;
		9747: Delta = 44'sb11111111111111111101111111111111111111110000;
		15728: Delta = 44'sb00000000000000000100000000000000000000010000;
		1923: Delta = 44'sb11111111111111111100000000000000000000010000;
		15696: Delta = 44'sb00000000000000000011111111111111111111110000;
		1891: Delta = 44'sb11111111111111111011111111111111111111110000;
		13821: Delta = 44'sb00000000000000001000000000000000000000010000;
		3830: Delta = 44'sb11111111111111111000000000000000000000010000;
		13789: Delta = 44'sb00000000000000000111111111111111111111110000;
		3798: Delta = 44'sb11111111111111110111111111111111111111110000;
		10007: Delta = 44'sb00000000000000010000000000000000000000010000;
		7644: Delta = 44'sb11111111111111110000000000000000000000010000;
		9975: Delta = 44'sb00000000000000001111111111111111111111110000;
		7612: Delta = 44'sb11111111111111101111111111111111111111110000;
		2379: Delta = 44'sb00000000000000100000000000000000000000010000;
		15272: Delta = 44'sb11111111111111100000000000000000000000010000;
		2347: Delta = 44'sb00000000000000011111111111111111111111110000;
		15240: Delta = 44'sb11111111111111011111111111111111111111110000;
		4742: Delta = 44'sb00000000000001000000000000000000000000010000;
		12909: Delta = 44'sb11111111111111000000000000000000000000010000;
		4710: Delta = 44'sb00000000000000111111111111111111111111110000;
		12877: Delta = 44'sb11111111111110111111111111111111111111110000;
		9468: Delta = 44'sb00000000000010000000000000000000000000010000;
		8183: Delta = 44'sb11111111111110000000000000000000000000010000;
		9436: Delta = 44'sb00000000000001111111111111111111111111110000;
		8151: Delta = 44'sb11111111111101111111111111111111111111110000;
		1301: Delta = 44'sb00000000000100000000000000000000000000010000;
		16350: Delta = 44'sb11111111111100000000000000000000000000010000;
		1269: Delta = 44'sb00000000000011111111111111111111111111110000;
		16318: Delta = 44'sb11111111111011111111111111111111111111110000;
		2586: Delta = 44'sb00000000001000000000000000000000000000010000;
		15065: Delta = 44'sb11111111111000000000000000000000000000010000;
		2554: Delta = 44'sb00000000000111111111111111111111111111110000;
		15033: Delta = 44'sb11111111110111111111111111111111111111110000;
		5156: Delta = 44'sb00000000010000000000000000000000000000010000;
		12495: Delta = 44'sb11111111110000000000000000000000000000010000;
		5124: Delta = 44'sb00000000001111111111111111111111111111110000;
		12463: Delta = 44'sb11111111101111111111111111111111111111110000;
		10296: Delta = 44'sb00000000100000000000000000000000000000010000;
		7355: Delta = 44'sb11111111100000000000000000000000000000010000;
		10264: Delta = 44'sb00000000011111111111111111111111111111110000;
		7323: Delta = 44'sb11111111011111111111111111111111111111110000;
		2957: Delta = 44'sb00000001000000000000000000000000000000010000;
		14694: Delta = 44'sb11111111000000000000000000000000000000010000;
		2925: Delta = 44'sb00000000111111111111111111111111111111110000;
		14662: Delta = 44'sb11111110111111111111111111111111111111110000;
		5898: Delta = 44'sb00000010000000000000000000000000000000010000;
		11753: Delta = 44'sb11111110000000000000000000000000000000010000;
		5866: Delta = 44'sb00000001111111111111111111111111111111110000;
		11721: Delta = 44'sb11111101111111111111111111111111111111110000;
		11780: Delta = 44'sb00000100000000000000000000000000000000010000;
		5871: Delta = 44'sb11111100000000000000000000000000000000010000;
		11748: Delta = 44'sb00000011111111111111111111111111111111110000;
		5839: Delta = 44'sb11111011111111111111111111111111111111110000;
		5925: Delta = 44'sb00001000000000000000000000000000000000010000;
		11726: Delta = 44'sb11111000000000000000000000000000000000010000;
		5893: Delta = 44'sb00000111111111111111111111111111111111110000;
		11694: Delta = 44'sb11110111111111111111111111111111111111110000;
		11834: Delta = 44'sb00010000000000000000000000000000000000010000;
		5817: Delta = 44'sb11110000000000000000000000000000000000010000;
		11802: Delta = 44'sb00001111111111111111111111111111111111110000;
		5785: Delta = 44'sb11101111111111111111111111111111111111110000;
		6033: Delta = 44'sb00100000000000000000000000000000000000010000;
		11618: Delta = 44'sb11100000000000000000000000000000000000010000;
		6001: Delta = 44'sb00011111111111111111111111111111111111110000;
		11586: Delta = 44'sb11011111111111111111111111111111111111110000;
		12050: Delta = 44'sb01000000000000000000000000000000000000010000;
		5601: Delta = 44'sb11000000000000000000000000000000000000010000;
		12018: Delta = 44'sb00111111111111111111111111111111111111110000;
		5569: Delta = 44'sb10111111111111111111111111111111111111110000;
		96: Delta = 44'sb00000000000000000000000000000000000001100000;
		17523: Delta = 44'sb11111111111111111111111111111111111110100000;
		160: Delta = 44'sb00000000000000000000000000000000000010100000;
		17459: Delta = 44'sb11111111111111111111111111111111111101100000;
		288: Delta = 44'sb00000000000000000000000000000000000100100000;
		17395: Delta = 44'sb11111111111111111111111111111111111100100000;
		224: Delta = 44'sb00000000000000000000000000000000000011100000;
		17331: Delta = 44'sb11111111111111111111111111111111111011100000;
		544: Delta = 44'sb00000000000000000000000000000000001000100000;
		17139: Delta = 44'sb11111111111111111111111111111111111000100000;
		480: Delta = 44'sb00000000000000000000000000000000000111100000;
		17075: Delta = 44'sb11111111111111111111111111111111110111100000;
		1056: Delta = 44'sb00000000000000000000000000000000010000100000;
		16627: Delta = 44'sb11111111111111111111111111111111110000100000;
		992: Delta = 44'sb00000000000000000000000000000000001111100000;
		16563: Delta = 44'sb11111111111111111111111111111111101111100000;
		2080: Delta = 44'sb00000000000000000000000000000000100000100000;
		15603: Delta = 44'sb11111111111111111111111111111111100000100000;
		2016: Delta = 44'sb00000000000000000000000000000000011111100000;
		15539: Delta = 44'sb11111111111111111111111111111111011111100000;
		4128: Delta = 44'sb00000000000000000000000000000001000000100000;
		13555: Delta = 44'sb11111111111111111111111111111111000000100000;
		4064: Delta = 44'sb00000000000000000000000000000000111111100000;
		13491: Delta = 44'sb11111111111111111111111111111110111111100000;
		8224: Delta = 44'sb00000000000000000000000000000010000000100000;
		9459: Delta = 44'sb11111111111111111111111111111110000000100000;
		8160: Delta = 44'sb00000000000000000000000000000001111111100000;
		9395: Delta = 44'sb11111111111111111111111111111101111111100000;
		16416: Delta = 44'sb00000000000000000000000000000100000000100000;
		1267: Delta = 44'sb11111111111111111111111111111100000000100000;
		16352: Delta = 44'sb00000000000000000000000000000011111111100000;
		1203: Delta = 44'sb11111111111111111111111111111011111111100000;
		15181: Delta = 44'sb00000000000000000000000000001000000000100000;
		2502: Delta = 44'sb11111111111111111111111111111000000000100000;
		15117: Delta = 44'sb00000000000000000000000000000111111111100000;
		2438: Delta = 44'sb11111111111111111111111111110111111111100000;
		12711: Delta = 44'sb00000000000000000000000000010000000000100000;
		4972: Delta = 44'sb11111111111111111111111111110000000000100000;
		12647: Delta = 44'sb00000000000000000000000000001111111111100000;
		4908: Delta = 44'sb11111111111111111111111111101111111111100000;
		7771: Delta = 44'sb00000000000000000000000000100000000000100000;
		9912: Delta = 44'sb11111111111111111111111111100000000000100000;
		7707: Delta = 44'sb00000000000000000000000000011111111111100000;
		9848: Delta = 44'sb11111111111111111111111111011111111111100000;
		15510: Delta = 44'sb00000000000000000000000001000000000000100000;
		2173: Delta = 44'sb11111111111111111111111111000000000000100000;
		15446: Delta = 44'sb00000000000000000000000000111111111111100000;
		2109: Delta = 44'sb11111111111111111111111110111111111111100000;
		13369: Delta = 44'sb00000000000000000000000010000000000000100000;
		4314: Delta = 44'sb11111111111111111111111110000000000000100000;
		13305: Delta = 44'sb00000000000000000000000001111111111111100000;
		4250: Delta = 44'sb11111111111111111111111101111111111111100000;
		9087: Delta = 44'sb00000000000000000000000100000000000000100000;
		8596: Delta = 44'sb11111111111111111111111100000000000000100000;
		9023: Delta = 44'sb00000000000000000000000011111111111111100000;
		8532: Delta = 44'sb11111111111111111111111011111111111111100000;
		523: Delta = 44'sb00000000000000000000001000000000000000100000;
		17160: Delta = 44'sb11111111111111111111111000000000000000100000;
		459: Delta = 44'sb00000000000000000000000111111111111111100000;
		17096: Delta = 44'sb11111111111111111111110111111111111111100000;
		1014: Delta = 44'sb00000000000000000000010000000000000000100000;
		16669: Delta = 44'sb11111111111111111111110000000000000000100000;
		950: Delta = 44'sb00000000000000000000001111111111111111100000;
		16605: Delta = 44'sb11111111111111111111101111111111111111100000;
		1996: Delta = 44'sb00000000000000000000100000000000000000100000;
		15687: Delta = 44'sb11111111111111111111100000000000000000100000;
		1932: Delta = 44'sb00000000000000000000011111111111111111100000;
		15623: Delta = 44'sb11111111111111111111011111111111111111100000;
		3960: Delta = 44'sb00000000000000000001000000000000000000100000;
		13723: Delta = 44'sb11111111111111111111000000000000000000100000;
		3896: Delta = 44'sb00000000000000000000111111111111111111100000;
		13659: Delta = 44'sb11111111111111111110111111111111111111100000;
		7888: Delta = 44'sb00000000000000000010000000000000000000100000;
		9795: Delta = 44'sb11111111111111111110000000000000000000100000;
		7824: Delta = 44'sb00000000000000000001111111111111111111100000;
		9731: Delta = 44'sb11111111111111111101111111111111111111100000;
		15744: Delta = 44'sb00000000000000000100000000000000000000100000;
		1939: Delta = 44'sb11111111111111111100000000000000000000100000;
		15680: Delta = 44'sb00000000000000000011111111111111111111100000;
		1875: Delta = 44'sb11111111111111111011111111111111111111100000;
		13837: Delta = 44'sb00000000000000001000000000000000000000100000;
		3846: Delta = 44'sb11111111111111111000000000000000000000100000;
		13773: Delta = 44'sb00000000000000000111111111111111111111100000;
		3782: Delta = 44'sb11111111111111110111111111111111111111100000;
		10023: Delta = 44'sb00000000000000010000000000000000000000100000;
		7660: Delta = 44'sb11111111111111110000000000000000000000100000;
		9959: Delta = 44'sb00000000000000001111111111111111111111100000;
		7596: Delta = 44'sb11111111111111101111111111111111111111100000;
		2395: Delta = 44'sb00000000000000100000000000000000000000100000;
		15288: Delta = 44'sb11111111111111100000000000000000000000100000;
		2331: Delta = 44'sb00000000000000011111111111111111111111100000;
		15224: Delta = 44'sb11111111111111011111111111111111111111100000;
		4758: Delta = 44'sb00000000000001000000000000000000000000100000;
		12925: Delta = 44'sb11111111111111000000000000000000000000100000;
		4694: Delta = 44'sb00000000000000111111111111111111111111100000;
		12861: Delta = 44'sb11111111111110111111111111111111111111100000;
		9484: Delta = 44'sb00000000000010000000000000000000000000100000;
		8199: Delta = 44'sb11111111111110000000000000000000000000100000;
		9420: Delta = 44'sb00000000000001111111111111111111111111100000;
		8135: Delta = 44'sb11111111111101111111111111111111111111100000;
		1317: Delta = 44'sb00000000000100000000000000000000000000100000;
		16366: Delta = 44'sb11111111111100000000000000000000000000100000;
		1253: Delta = 44'sb00000000000011111111111111111111111111100000;
		16302: Delta = 44'sb11111111111011111111111111111111111111100000;
		2602: Delta = 44'sb00000000001000000000000000000000000000100000;
		15081: Delta = 44'sb11111111111000000000000000000000000000100000;
		2538: Delta = 44'sb00000000000111111111111111111111111111100000;
		15017: Delta = 44'sb11111111110111111111111111111111111111100000;
		5172: Delta = 44'sb00000000010000000000000000000000000000100000;
		12511: Delta = 44'sb11111111110000000000000000000000000000100000;
		5108: Delta = 44'sb00000000001111111111111111111111111111100000;
		12447: Delta = 44'sb11111111101111111111111111111111111111100000;
		10312: Delta = 44'sb00000000100000000000000000000000000000100000;
		7371: Delta = 44'sb11111111100000000000000000000000000000100000;
		10248: Delta = 44'sb00000000011111111111111111111111111111100000;
		7307: Delta = 44'sb11111111011111111111111111111111111111100000;
		2973: Delta = 44'sb00000001000000000000000000000000000000100000;
		14710: Delta = 44'sb11111111000000000000000000000000000000100000;
		2909: Delta = 44'sb00000000111111111111111111111111111111100000;
		14646: Delta = 44'sb11111110111111111111111111111111111111100000;
		5914: Delta = 44'sb00000010000000000000000000000000000000100000;
		11769: Delta = 44'sb11111110000000000000000000000000000000100000;
		5850: Delta = 44'sb00000001111111111111111111111111111111100000;
		11705: Delta = 44'sb11111101111111111111111111111111111111100000;
		11796: Delta = 44'sb00000100000000000000000000000000000000100000;
		5887: Delta = 44'sb11111100000000000000000000000000000000100000;
		11732: Delta = 44'sb00000011111111111111111111111111111111100000;
		5823: Delta = 44'sb11111011111111111111111111111111111111100000;
		5941: Delta = 44'sb00001000000000000000000000000000000000100000;
		11742: Delta = 44'sb11111000000000000000000000000000000000100000;
		5877: Delta = 44'sb00000111111111111111111111111111111111100000;
		11678: Delta = 44'sb11110111111111111111111111111111111111100000;
		11850: Delta = 44'sb00010000000000000000000000000000000000100000;
		5833: Delta = 44'sb11110000000000000000000000000000000000100000;
		11786: Delta = 44'sb00001111111111111111111111111111111111100000;
		5769: Delta = 44'sb11101111111111111111111111111111111111100000;
		6049: Delta = 44'sb00100000000000000000000000000000000000100000;
		11634: Delta = 44'sb11100000000000000000000000000000000000100000;
		5985: Delta = 44'sb00011111111111111111111111111111111111100000;
		11570: Delta = 44'sb11011111111111111111111111111111111111100000;
		12066: Delta = 44'sb01000000000000000000000000000000000000100000;
		5617: Delta = 44'sb11000000000000000000000000000000000000100000;
		12002: Delta = 44'sb00111111111111111111111111111111111111100000;
		5553: Delta = 44'sb10111111111111111111111111111111111111100000;
		192: Delta = 44'sb00000000000000000000000000000000000011000000;
		17427: Delta = 44'sb11111111111111111111111111111111111101000000;
		320: Delta = 44'sb00000000000000000000000000000000000101000000;
		17299: Delta = 44'sb11111111111111111111111111111111111011000000;
		576: Delta = 44'sb00000000000000000000000000000000001001000000;
		17171: Delta = 44'sb11111111111111111111111111111111111001000000;
		448: Delta = 44'sb00000000000000000000000000000000000111000000;
		17043: Delta = 44'sb11111111111111111111111111111111110111000000;
		1088: Delta = 44'sb00000000000000000000000000000000010001000000;
		16659: Delta = 44'sb11111111111111111111111111111111110001000000;
		960: Delta = 44'sb00000000000000000000000000000000001111000000;
		16531: Delta = 44'sb11111111111111111111111111111111101111000000;
		2112: Delta = 44'sb00000000000000000000000000000000100001000000;
		15635: Delta = 44'sb11111111111111111111111111111111100001000000;
		1984: Delta = 44'sb00000000000000000000000000000000011111000000;
		15507: Delta = 44'sb11111111111111111111111111111111011111000000;
		4160: Delta = 44'sb00000000000000000000000000000001000001000000;
		13587: Delta = 44'sb11111111111111111111111111111111000001000000;
		4032: Delta = 44'sb00000000000000000000000000000000111111000000;
		13459: Delta = 44'sb11111111111111111111111111111110111111000000;
		8256: Delta = 44'sb00000000000000000000000000000010000001000000;
		9491: Delta = 44'sb11111111111111111111111111111110000001000000;
		8128: Delta = 44'sb00000000000000000000000000000001111111000000;
		9363: Delta = 44'sb11111111111111111111111111111101111111000000;
		16448: Delta = 44'sb00000000000000000000000000000100000001000000;
		1299: Delta = 44'sb11111111111111111111111111111100000001000000;
		16320: Delta = 44'sb00000000000000000000000000000011111111000000;
		1171: Delta = 44'sb11111111111111111111111111111011111111000000;
		15213: Delta = 44'sb00000000000000000000000000001000000001000000;
		2534: Delta = 44'sb11111111111111111111111111111000000001000000;
		15085: Delta = 44'sb00000000000000000000000000000111111111000000;
		2406: Delta = 44'sb11111111111111111111111111110111111111000000;
		12743: Delta = 44'sb00000000000000000000000000010000000001000000;
		5004: Delta = 44'sb11111111111111111111111111110000000001000000;
		12615: Delta = 44'sb00000000000000000000000000001111111111000000;
		4876: Delta = 44'sb11111111111111111111111111101111111111000000;
		7803: Delta = 44'sb00000000000000000000000000100000000001000000;
		9944: Delta = 44'sb11111111111111111111111111100000000001000000;
		7675: Delta = 44'sb00000000000000000000000000011111111111000000;
		9816: Delta = 44'sb11111111111111111111111111011111111111000000;
		15542: Delta = 44'sb00000000000000000000000001000000000001000000;
		2205: Delta = 44'sb11111111111111111111111111000000000001000000;
		15414: Delta = 44'sb00000000000000000000000000111111111111000000;
		2077: Delta = 44'sb11111111111111111111111110111111111111000000;
		13401: Delta = 44'sb00000000000000000000000010000000000001000000;
		4346: Delta = 44'sb11111111111111111111111110000000000001000000;
		13273: Delta = 44'sb00000000000000000000000001111111111111000000;
		4218: Delta = 44'sb11111111111111111111111101111111111111000000;
		9119: Delta = 44'sb00000000000000000000000100000000000001000000;
		8628: Delta = 44'sb11111111111111111111111100000000000001000000;
		8991: Delta = 44'sb00000000000000000000000011111111111111000000;
		8500: Delta = 44'sb11111111111111111111111011111111111111000000;
		555: Delta = 44'sb00000000000000000000001000000000000001000000;
		17192: Delta = 44'sb11111111111111111111111000000000000001000000;
		427: Delta = 44'sb00000000000000000000000111111111111111000000;
		17064: Delta = 44'sb11111111111111111111110111111111111111000000;
		1046: Delta = 44'sb00000000000000000000010000000000000001000000;
		16701: Delta = 44'sb11111111111111111111110000000000000001000000;
		918: Delta = 44'sb00000000000000000000001111111111111111000000;
		16573: Delta = 44'sb11111111111111111111101111111111111111000000;
		2028: Delta = 44'sb00000000000000000000100000000000000001000000;
		15719: Delta = 44'sb11111111111111111111100000000000000001000000;
		1900: Delta = 44'sb00000000000000000000011111111111111111000000;
		15591: Delta = 44'sb11111111111111111111011111111111111111000000;
		3992: Delta = 44'sb00000000000000000001000000000000000001000000;
		13755: Delta = 44'sb11111111111111111111000000000000000001000000;
		3864: Delta = 44'sb00000000000000000000111111111111111111000000;
		13627: Delta = 44'sb11111111111111111110111111111111111111000000;
		7920: Delta = 44'sb00000000000000000010000000000000000001000000;
		9827: Delta = 44'sb11111111111111111110000000000000000001000000;
		7792: Delta = 44'sb00000000000000000001111111111111111111000000;
		9699: Delta = 44'sb11111111111111111101111111111111111111000000;
		15776: Delta = 44'sb00000000000000000100000000000000000001000000;
		1971: Delta = 44'sb11111111111111111100000000000000000001000000;
		15648: Delta = 44'sb00000000000000000011111111111111111111000000;
		1843: Delta = 44'sb11111111111111111011111111111111111111000000;
		13869: Delta = 44'sb00000000000000001000000000000000000001000000;
		3878: Delta = 44'sb11111111111111111000000000000000000001000000;
		13741: Delta = 44'sb00000000000000000111111111111111111111000000;
		3750: Delta = 44'sb11111111111111110111111111111111111111000000;
		10055: Delta = 44'sb00000000000000010000000000000000000001000000;
		7692: Delta = 44'sb11111111111111110000000000000000000001000000;
		9927: Delta = 44'sb00000000000000001111111111111111111111000000;
		7564: Delta = 44'sb11111111111111101111111111111111111111000000;
		2427: Delta = 44'sb00000000000000100000000000000000000001000000;
		15320: Delta = 44'sb11111111111111100000000000000000000001000000;
		2299: Delta = 44'sb00000000000000011111111111111111111111000000;
		15192: Delta = 44'sb11111111111111011111111111111111111111000000;
		4790: Delta = 44'sb00000000000001000000000000000000000001000000;
		12957: Delta = 44'sb11111111111111000000000000000000000001000000;
		4662: Delta = 44'sb00000000000000111111111111111111111111000000;
		12829: Delta = 44'sb11111111111110111111111111111111111111000000;
		9516: Delta = 44'sb00000000000010000000000000000000000001000000;
		8231: Delta = 44'sb11111111111110000000000000000000000001000000;
		9388: Delta = 44'sb00000000000001111111111111111111111111000000;
		8103: Delta = 44'sb11111111111101111111111111111111111111000000;
		1349: Delta = 44'sb00000000000100000000000000000000000001000000;
		16398: Delta = 44'sb11111111111100000000000000000000000001000000;
		1221: Delta = 44'sb00000000000011111111111111111111111111000000;
		16270: Delta = 44'sb11111111111011111111111111111111111111000000;
		2634: Delta = 44'sb00000000001000000000000000000000000001000000;
		15113: Delta = 44'sb11111111111000000000000000000000000001000000;
		2506: Delta = 44'sb00000000000111111111111111111111111111000000;
		14985: Delta = 44'sb11111111110111111111111111111111111111000000;
		5204: Delta = 44'sb00000000010000000000000000000000000001000000;
		12543: Delta = 44'sb11111111110000000000000000000000000001000000;
		5076: Delta = 44'sb00000000001111111111111111111111111111000000;
		12415: Delta = 44'sb11111111101111111111111111111111111111000000;
		10344: Delta = 44'sb00000000100000000000000000000000000001000000;
		7403: Delta = 44'sb11111111100000000000000000000000000001000000;
		10216: Delta = 44'sb00000000011111111111111111111111111111000000;
		7275: Delta = 44'sb11111111011111111111111111111111111111000000;
		3005: Delta = 44'sb00000001000000000000000000000000000001000000;
		14742: Delta = 44'sb11111111000000000000000000000000000001000000;
		2877: Delta = 44'sb00000000111111111111111111111111111111000000;
		14614: Delta = 44'sb11111110111111111111111111111111111111000000;
		5946: Delta = 44'sb00000010000000000000000000000000000001000000;
		11801: Delta = 44'sb11111110000000000000000000000000000001000000;
		5818: Delta = 44'sb00000001111111111111111111111111111111000000;
		11673: Delta = 44'sb11111101111111111111111111111111111111000000;
		11828: Delta = 44'sb00000100000000000000000000000000000001000000;
		5919: Delta = 44'sb11111100000000000000000000000000000001000000;
		11700: Delta = 44'sb00000011111111111111111111111111111111000000;
		5791: Delta = 44'sb11111011111111111111111111111111111111000000;
		5973: Delta = 44'sb00001000000000000000000000000000000001000000;
		11774: Delta = 44'sb11111000000000000000000000000000000001000000;
		5845: Delta = 44'sb00000111111111111111111111111111111111000000;
		11646: Delta = 44'sb11110111111111111111111111111111111111000000;
		11882: Delta = 44'sb00010000000000000000000000000000000001000000;
		5865: Delta = 44'sb11110000000000000000000000000000000001000000;
		11754: Delta = 44'sb00001111111111111111111111111111111111000000;
		5737: Delta = 44'sb11101111111111111111111111111111111111000000;
		6081: Delta = 44'sb00100000000000000000000000000000000001000000;
		11666: Delta = 44'sb11100000000000000000000000000000000001000000;
		5953: Delta = 44'sb00011111111111111111111111111111111111000000;
		11538: Delta = 44'sb11011111111111111111111111111111111111000000;
		12098: Delta = 44'sb01000000000000000000000000000000000001000000;
		5649: Delta = 44'sb11000000000000000000000000000000000001000000;
		11970: Delta = 44'sb00111111111111111111111111111111111111000000;
		5521: Delta = 44'sb10111111111111111111111111111111111111000000;
		384: Delta = 44'sb00000000000000000000000000000000000110000000;
		17235: Delta = 44'sb11111111111111111111111111111111111010000000;
		640: Delta = 44'sb00000000000000000000000000000000001010000000;
		16979: Delta = 44'sb11111111111111111111111111111111110110000000;
		1152: Delta = 44'sb00000000000000000000000000000000010010000000;
		16723: Delta = 44'sb11111111111111111111111111111111110010000000;
		896: Delta = 44'sb00000000000000000000000000000000001110000000;
		16467: Delta = 44'sb11111111111111111111111111111111101110000000;
		2176: Delta = 44'sb00000000000000000000000000000000100010000000;
		15699: Delta = 44'sb11111111111111111111111111111111100010000000;
		1920: Delta = 44'sb00000000000000000000000000000000011110000000;
		15443: Delta = 44'sb11111111111111111111111111111111011110000000;
		4224: Delta = 44'sb00000000000000000000000000000001000010000000;
		13651: Delta = 44'sb11111111111111111111111111111111000010000000;
		3968: Delta = 44'sb00000000000000000000000000000000111110000000;
		13395: Delta = 44'sb11111111111111111111111111111110111110000000;
		8320: Delta = 44'sb00000000000000000000000000000010000010000000;
		9555: Delta = 44'sb11111111111111111111111111111110000010000000;
		8064: Delta = 44'sb00000000000000000000000000000001111110000000;
		9299: Delta = 44'sb11111111111111111111111111111101111110000000;
		16512: Delta = 44'sb00000000000000000000000000000100000010000000;
		1363: Delta = 44'sb11111111111111111111111111111100000010000000;
		16256: Delta = 44'sb00000000000000000000000000000011111110000000;
		1107: Delta = 44'sb11111111111111111111111111111011111110000000;
		15277: Delta = 44'sb00000000000000000000000000001000000010000000;
		2598: Delta = 44'sb11111111111111111111111111111000000010000000;
		15021: Delta = 44'sb00000000000000000000000000000111111110000000;
		2342: Delta = 44'sb11111111111111111111111111110111111110000000;
		12807: Delta = 44'sb00000000000000000000000000010000000010000000;
		5068: Delta = 44'sb11111111111111111111111111110000000010000000;
		12551: Delta = 44'sb00000000000000000000000000001111111110000000;
		4812: Delta = 44'sb11111111111111111111111111101111111110000000;
		7867: Delta = 44'sb00000000000000000000000000100000000010000000;
		10008: Delta = 44'sb11111111111111111111111111100000000010000000;
		7611: Delta = 44'sb00000000000000000000000000011111111110000000;
		9752: Delta = 44'sb11111111111111111111111111011111111110000000;
		15606: Delta = 44'sb00000000000000000000000001000000000010000000;
		2269: Delta = 44'sb11111111111111111111111111000000000010000000;
		15350: Delta = 44'sb00000000000000000000000000111111111110000000;
		2013: Delta = 44'sb11111111111111111111111110111111111110000000;
		13465: Delta = 44'sb00000000000000000000000010000000000010000000;
		4410: Delta = 44'sb11111111111111111111111110000000000010000000;
		13209: Delta = 44'sb00000000000000000000000001111111111110000000;
		4154: Delta = 44'sb11111111111111111111111101111111111110000000;
		9183: Delta = 44'sb00000000000000000000000100000000000010000000;
		8692: Delta = 44'sb11111111111111111111111100000000000010000000;
		8927: Delta = 44'sb00000000000000000000000011111111111110000000;
		8436: Delta = 44'sb11111111111111111111111011111111111110000000;
		619: Delta = 44'sb00000000000000000000001000000000000010000000;
		17256: Delta = 44'sb11111111111111111111111000000000000010000000;
		363: Delta = 44'sb00000000000000000000000111111111111110000000;
		17000: Delta = 44'sb11111111111111111111110111111111111110000000;
		1110: Delta = 44'sb00000000000000000000010000000000000010000000;
		16765: Delta = 44'sb11111111111111111111110000000000000010000000;
		854: Delta = 44'sb00000000000000000000001111111111111110000000;
		16509: Delta = 44'sb11111111111111111111101111111111111110000000;
		2092: Delta = 44'sb00000000000000000000100000000000000010000000;
		15783: Delta = 44'sb11111111111111111111100000000000000010000000;
		1836: Delta = 44'sb00000000000000000000011111111111111110000000;
		15527: Delta = 44'sb11111111111111111111011111111111111110000000;
		4056: Delta = 44'sb00000000000000000001000000000000000010000000;
		13819: Delta = 44'sb11111111111111111111000000000000000010000000;
		3800: Delta = 44'sb00000000000000000000111111111111111110000000;
		13563: Delta = 44'sb11111111111111111110111111111111111110000000;
		7984: Delta = 44'sb00000000000000000010000000000000000010000000;
		9891: Delta = 44'sb11111111111111111110000000000000000010000000;
		7728: Delta = 44'sb00000000000000000001111111111111111110000000;
		9635: Delta = 44'sb11111111111111111101111111111111111110000000;
		15840: Delta = 44'sb00000000000000000100000000000000000010000000;
		2035: Delta = 44'sb11111111111111111100000000000000000010000000;
		15584: Delta = 44'sb00000000000000000011111111111111111110000000;
		1779: Delta = 44'sb11111111111111111011111111111111111110000000;
		13933: Delta = 44'sb00000000000000001000000000000000000010000000;
		3942: Delta = 44'sb11111111111111111000000000000000000010000000;
		13677: Delta = 44'sb00000000000000000111111111111111111110000000;
		3686: Delta = 44'sb11111111111111110111111111111111111110000000;
		10119: Delta = 44'sb00000000000000010000000000000000000010000000;
		7756: Delta = 44'sb11111111111111110000000000000000000010000000;
		9863: Delta = 44'sb00000000000000001111111111111111111110000000;
		7500: Delta = 44'sb11111111111111101111111111111111111110000000;
		2491: Delta = 44'sb00000000000000100000000000000000000010000000;
		15384: Delta = 44'sb11111111111111100000000000000000000010000000;
		2235: Delta = 44'sb00000000000000011111111111111111111110000000;
		15128: Delta = 44'sb11111111111111011111111111111111111110000000;
		4854: Delta = 44'sb00000000000001000000000000000000000010000000;
		13021: Delta = 44'sb11111111111111000000000000000000000010000000;
		4598: Delta = 44'sb00000000000000111111111111111111111110000000;
		12765: Delta = 44'sb11111111111110111111111111111111111110000000;
		9580: Delta = 44'sb00000000000010000000000000000000000010000000;
		8295: Delta = 44'sb11111111111110000000000000000000000010000000;
		9324: Delta = 44'sb00000000000001111111111111111111111110000000;
		8039: Delta = 44'sb11111111111101111111111111111111111110000000;
		1413: Delta = 44'sb00000000000100000000000000000000000010000000;
		16462: Delta = 44'sb11111111111100000000000000000000000010000000;
		1157: Delta = 44'sb00000000000011111111111111111111111110000000;
		16206: Delta = 44'sb11111111111011111111111111111111111110000000;
		2698: Delta = 44'sb00000000001000000000000000000000000010000000;
		15177: Delta = 44'sb11111111111000000000000000000000000010000000;
		2442: Delta = 44'sb00000000000111111111111111111111111110000000;
		14921: Delta = 44'sb11111111110111111111111111111111111110000000;
		5268: Delta = 44'sb00000000010000000000000000000000000010000000;
		12607: Delta = 44'sb11111111110000000000000000000000000010000000;
		5012: Delta = 44'sb00000000001111111111111111111111111110000000;
		12351: Delta = 44'sb11111111101111111111111111111111111110000000;
		10408: Delta = 44'sb00000000100000000000000000000000000010000000;
		7467: Delta = 44'sb11111111100000000000000000000000000010000000;
		10152: Delta = 44'sb00000000011111111111111111111111111110000000;
		7211: Delta = 44'sb11111111011111111111111111111111111110000000;
		3069: Delta = 44'sb00000001000000000000000000000000000010000000;
		14806: Delta = 44'sb11111111000000000000000000000000000010000000;
		2813: Delta = 44'sb00000000111111111111111111111111111110000000;
		14550: Delta = 44'sb11111110111111111111111111111111111110000000;
		6010: Delta = 44'sb00000010000000000000000000000000000010000000;
		11865: Delta = 44'sb11111110000000000000000000000000000010000000;
		5754: Delta = 44'sb00000001111111111111111111111111111110000000;
		11609: Delta = 44'sb11111101111111111111111111111111111110000000;
		11892: Delta = 44'sb00000100000000000000000000000000000010000000;
		5983: Delta = 44'sb11111100000000000000000000000000000010000000;
		11636: Delta = 44'sb00000011111111111111111111111111111110000000;
		5727: Delta = 44'sb11111011111111111111111111111111111110000000;
		6037: Delta = 44'sb00001000000000000000000000000000000010000000;
		11838: Delta = 44'sb11111000000000000000000000000000000010000000;
		5781: Delta = 44'sb00000111111111111111111111111111111110000000;
		11582: Delta = 44'sb11110111111111111111111111111111111110000000;
		11946: Delta = 44'sb00010000000000000000000000000000000010000000;
		5929: Delta = 44'sb11110000000000000000000000000000000010000000;
		11690: Delta = 44'sb00001111111111111111111111111111111110000000;
		5673: Delta = 44'sb11101111111111111111111111111111111110000000;
		6145: Delta = 44'sb00100000000000000000000000000000000010000000;
		11730: Delta = 44'sb11100000000000000000000000000000000010000000;
		5889: Delta = 44'sb00011111111111111111111111111111111110000000;
		11474: Delta = 44'sb11011111111111111111111111111111111110000000;
		12162: Delta = 44'sb01000000000000000000000000000000000010000000;
		5713: Delta = 44'sb11000000000000000000000000000000000010000000;
		11906: Delta = 44'sb00111111111111111111111111111111111110000000;
		5457: Delta = 44'sb10111111111111111111111111111111111110000000;
		768: Delta = 44'sb00000000000000000000000000000000001100000000;
		16851: Delta = 44'sb11111111111111111111111111111111110100000000;
		1280: Delta = 44'sb00000000000000000000000000000000010100000000;
		16339: Delta = 44'sb11111111111111111111111111111111101100000000;
		2304: Delta = 44'sb00000000000000000000000000000000100100000000;
		15827: Delta = 44'sb11111111111111111111111111111111100100000000;
		1792: Delta = 44'sb00000000000000000000000000000000011100000000;
		15315: Delta = 44'sb11111111111111111111111111111111011100000000;
		4352: Delta = 44'sb00000000000000000000000000000001000100000000;
		13779: Delta = 44'sb11111111111111111111111111111111000100000000;
		3840: Delta = 44'sb00000000000000000000000000000000111100000000;
		13267: Delta = 44'sb11111111111111111111111111111110111100000000;
		8448: Delta = 44'sb00000000000000000000000000000010000100000000;
		9683: Delta = 44'sb11111111111111111111111111111110000100000000;
		7936: Delta = 44'sb00000000000000000000000000000001111100000000;
		9171: Delta = 44'sb11111111111111111111111111111101111100000000;
		16640: Delta = 44'sb00000000000000000000000000000100000100000000;
		1491: Delta = 44'sb11111111111111111111111111111100000100000000;
		16128: Delta = 44'sb00000000000000000000000000000011111100000000;
		979: Delta = 44'sb11111111111111111111111111111011111100000000;
		15405: Delta = 44'sb00000000000000000000000000001000000100000000;
		2726: Delta = 44'sb11111111111111111111111111111000000100000000;
		14893: Delta = 44'sb00000000000000000000000000000111111100000000;
		2214: Delta = 44'sb11111111111111111111111111110111111100000000;
		12935: Delta = 44'sb00000000000000000000000000010000000100000000;
		5196: Delta = 44'sb11111111111111111111111111110000000100000000;
		12423: Delta = 44'sb00000000000000000000000000001111111100000000;
		4684: Delta = 44'sb11111111111111111111111111101111111100000000;
		7995: Delta = 44'sb00000000000000000000000000100000000100000000;
		10136: Delta = 44'sb11111111111111111111111111100000000100000000;
		7483: Delta = 44'sb00000000000000000000000000011111111100000000;
		9624: Delta = 44'sb11111111111111111111111111011111111100000000;
		15734: Delta = 44'sb00000000000000000000000001000000000100000000;
		2397: Delta = 44'sb11111111111111111111111111000000000100000000;
		15222: Delta = 44'sb00000000000000000000000000111111111100000000;
		1885: Delta = 44'sb11111111111111111111111110111111111100000000;
		13593: Delta = 44'sb00000000000000000000000010000000000100000000;
		4538: Delta = 44'sb11111111111111111111111110000000000100000000;
		13081: Delta = 44'sb00000000000000000000000001111111111100000000;
		4026: Delta = 44'sb11111111111111111111111101111111111100000000;
		9311: Delta = 44'sb00000000000000000000000100000000000100000000;
		8820: Delta = 44'sb11111111111111111111111100000000000100000000;
		8799: Delta = 44'sb00000000000000000000000011111111111100000000;
		8308: Delta = 44'sb11111111111111111111111011111111111100000000;
		747: Delta = 44'sb00000000000000000000001000000000000100000000;
		17384: Delta = 44'sb11111111111111111111111000000000000100000000;
		235: Delta = 44'sb00000000000000000000000111111111111100000000;
		16872: Delta = 44'sb11111111111111111111110111111111111100000000;
		1238: Delta = 44'sb00000000000000000000010000000000000100000000;
		16893: Delta = 44'sb11111111111111111111110000000000000100000000;
		726: Delta = 44'sb00000000000000000000001111111111111100000000;
		16381: Delta = 44'sb11111111111111111111101111111111111100000000;
		2220: Delta = 44'sb00000000000000000000100000000000000100000000;
		15911: Delta = 44'sb11111111111111111111100000000000000100000000;
		1708: Delta = 44'sb00000000000000000000011111111111111100000000;
		15399: Delta = 44'sb11111111111111111111011111111111111100000000;
		4184: Delta = 44'sb00000000000000000001000000000000000100000000;
		13947: Delta = 44'sb11111111111111111111000000000000000100000000;
		3672: Delta = 44'sb00000000000000000000111111111111111100000000;
		13435: Delta = 44'sb11111111111111111110111111111111111100000000;
		8112: Delta = 44'sb00000000000000000010000000000000000100000000;
		10019: Delta = 44'sb11111111111111111110000000000000000100000000;
		7600: Delta = 44'sb00000000000000000001111111111111111100000000;
		9507: Delta = 44'sb11111111111111111101111111111111111100000000;
		15968: Delta = 44'sb00000000000000000100000000000000000100000000;
		2163: Delta = 44'sb11111111111111111100000000000000000100000000;
		15456: Delta = 44'sb00000000000000000011111111111111111100000000;
		1651: Delta = 44'sb11111111111111111011111111111111111100000000;
		14061: Delta = 44'sb00000000000000001000000000000000000100000000;
		4070: Delta = 44'sb11111111111111111000000000000000000100000000;
		13549: Delta = 44'sb00000000000000000111111111111111111100000000;
		3558: Delta = 44'sb11111111111111110111111111111111111100000000;
		10247: Delta = 44'sb00000000000000010000000000000000000100000000;
		7884: Delta = 44'sb11111111111111110000000000000000000100000000;
		9735: Delta = 44'sb00000000000000001111111111111111111100000000;
		7372: Delta = 44'sb11111111111111101111111111111111111100000000;
		2619: Delta = 44'sb00000000000000100000000000000000000100000000;
		15512: Delta = 44'sb11111111111111100000000000000000000100000000;
		2107: Delta = 44'sb00000000000000011111111111111111111100000000;
		15000: Delta = 44'sb11111111111111011111111111111111111100000000;
		4982: Delta = 44'sb00000000000001000000000000000000000100000000;
		13149: Delta = 44'sb11111111111111000000000000000000000100000000;
		4470: Delta = 44'sb00000000000000111111111111111111111100000000;
		12637: Delta = 44'sb11111111111110111111111111111111111100000000;
		9708: Delta = 44'sb00000000000010000000000000000000000100000000;
		8423: Delta = 44'sb11111111111110000000000000000000000100000000;
		9196: Delta = 44'sb00000000000001111111111111111111111100000000;
		7911: Delta = 44'sb11111111111101111111111111111111111100000000;
		1541: Delta = 44'sb00000000000100000000000000000000000100000000;
		16590: Delta = 44'sb11111111111100000000000000000000000100000000;
		1029: Delta = 44'sb00000000000011111111111111111111111100000000;
		16078: Delta = 44'sb11111111111011111111111111111111111100000000;
		2826: Delta = 44'sb00000000001000000000000000000000000100000000;
		15305: Delta = 44'sb11111111111000000000000000000000000100000000;
		2314: Delta = 44'sb00000000000111111111111111111111111100000000;
		14793: Delta = 44'sb11111111110111111111111111111111111100000000;
		5396: Delta = 44'sb00000000010000000000000000000000000100000000;
		12735: Delta = 44'sb11111111110000000000000000000000000100000000;
		4884: Delta = 44'sb00000000001111111111111111111111111100000000;
		12223: Delta = 44'sb11111111101111111111111111111111111100000000;
		10536: Delta = 44'sb00000000100000000000000000000000000100000000;
		7595: Delta = 44'sb11111111100000000000000000000000000100000000;
		10024: Delta = 44'sb00000000011111111111111111111111111100000000;
		7083: Delta = 44'sb11111111011111111111111111111111111100000000;
		3197: Delta = 44'sb00000001000000000000000000000000000100000000;
		14934: Delta = 44'sb11111111000000000000000000000000000100000000;
		2685: Delta = 44'sb00000000111111111111111111111111111100000000;
		14422: Delta = 44'sb11111110111111111111111111111111111100000000;
		6138: Delta = 44'sb00000010000000000000000000000000000100000000;
		11993: Delta = 44'sb11111110000000000000000000000000000100000000;
		5626: Delta = 44'sb00000001111111111111111111111111111100000000;
		11481: Delta = 44'sb11111101111111111111111111111111111100000000;
		12020: Delta = 44'sb00000100000000000000000000000000000100000000;
		6111: Delta = 44'sb11111100000000000000000000000000000100000000;
		11508: Delta = 44'sb00000011111111111111111111111111111100000000;
		5599: Delta = 44'sb11111011111111111111111111111111111100000000;
		6165: Delta = 44'sb00001000000000000000000000000000000100000000;
		11966: Delta = 44'sb11111000000000000000000000000000000100000000;
		5653: Delta = 44'sb00000111111111111111111111111111111100000000;
		11454: Delta = 44'sb11110111111111111111111111111111111100000000;
		12074: Delta = 44'sb00010000000000000000000000000000000100000000;
		6057: Delta = 44'sb11110000000000000000000000000000000100000000;
		11562: Delta = 44'sb00001111111111111111111111111111111100000000;
		5545: Delta = 44'sb11101111111111111111111111111111111100000000;
		6273: Delta = 44'sb00100000000000000000000000000000000100000000;
		11858: Delta = 44'sb11100000000000000000000000000000000100000000;
		5761: Delta = 44'sb00011111111111111111111111111111111100000000;
		11346: Delta = 44'sb11011111111111111111111111111111111100000000;
		12290: Delta = 44'sb01000000000000000000000000000000000100000000;
		5841: Delta = 44'sb11000000000000000000000000000000000100000000;
		11778: Delta = 44'sb00111111111111111111111111111111111100000000;
		5329: Delta = 44'sb10111111111111111111111111111111111100000000;
		1536: Delta = 44'sb00000000000000000000000000000000011000000000;
		16083: Delta = 44'sb11111111111111111111111111111111101000000000;
		2560: Delta = 44'sb00000000000000000000000000000000101000000000;
		15059: Delta = 44'sb11111111111111111111111111111111011000000000;
		4608: Delta = 44'sb00000000000000000000000000000001001000000000;
		14035: Delta = 44'sb11111111111111111111111111111111001000000000;
		3584: Delta = 44'sb00000000000000000000000000000000111000000000;
		13011: Delta = 44'sb11111111111111111111111111111110111000000000;
		8704: Delta = 44'sb00000000000000000000000000000010001000000000;
		9939: Delta = 44'sb11111111111111111111111111111110001000000000;
		7680: Delta = 44'sb00000000000000000000000000000001111000000000;
		8915: Delta = 44'sb11111111111111111111111111111101111000000000;
		16896: Delta = 44'sb00000000000000000000000000000100001000000000;
		1747: Delta = 44'sb11111111111111111111111111111100001000000000;
		15872: Delta = 44'sb00000000000000000000000000000011111000000000;
		723: Delta = 44'sb11111111111111111111111111111011111000000000;
		15661: Delta = 44'sb00000000000000000000000000001000001000000000;
		2982: Delta = 44'sb11111111111111111111111111111000001000000000;
		14637: Delta = 44'sb00000000000000000000000000000111111000000000;
		1958: Delta = 44'sb11111111111111111111111111110111111000000000;
		13191: Delta = 44'sb00000000000000000000000000010000001000000000;
		5452: Delta = 44'sb11111111111111111111111111110000001000000000;
		12167: Delta = 44'sb00000000000000000000000000001111111000000000;
		4428: Delta = 44'sb11111111111111111111111111101111111000000000;
		8251: Delta = 44'sb00000000000000000000000000100000001000000000;
		10392: Delta = 44'sb11111111111111111111111111100000001000000000;
		7227: Delta = 44'sb00000000000000000000000000011111111000000000;
		9368: Delta = 44'sb11111111111111111111111111011111111000000000;
		15990: Delta = 44'sb00000000000000000000000001000000001000000000;
		2653: Delta = 44'sb11111111111111111111111111000000001000000000;
		14966: Delta = 44'sb00000000000000000000000000111111111000000000;
		1629: Delta = 44'sb11111111111111111111111110111111111000000000;
		13849: Delta = 44'sb00000000000000000000000010000000001000000000;
		4794: Delta = 44'sb11111111111111111111111110000000001000000000;
		12825: Delta = 44'sb00000000000000000000000001111111111000000000;
		3770: Delta = 44'sb11111111111111111111111101111111111000000000;
		9567: Delta = 44'sb00000000000000000000000100000000001000000000;
		9076: Delta = 44'sb11111111111111111111111100000000001000000000;
		8543: Delta = 44'sb00000000000000000000000011111111111000000000;
		8052: Delta = 44'sb11111111111111111111111011111111111000000000;
		1003: Delta = 44'sb00000000000000000000001000000000001000000000;
		21: Delta = 44'sb11111111111111111111111000000000001000000000;
		17598: Delta = 44'sb00000000000000000000000111111111111000000000;
		16616: Delta = 44'sb11111111111111111111110111111111111000000000;
		1494: Delta = 44'sb00000000000000000000010000000000001000000000;
		17149: Delta = 44'sb11111111111111111111110000000000001000000000;
		470: Delta = 44'sb00000000000000000000001111111111111000000000;
		16125: Delta = 44'sb11111111111111111111101111111111111000000000;
		2476: Delta = 44'sb00000000000000000000100000000000001000000000;
		16167: Delta = 44'sb11111111111111111111100000000000001000000000;
		1452: Delta = 44'sb00000000000000000000011111111111111000000000;
		15143: Delta = 44'sb11111111111111111111011111111111111000000000;
		4440: Delta = 44'sb00000000000000000001000000000000001000000000;
		14203: Delta = 44'sb11111111111111111111000000000000001000000000;
		3416: Delta = 44'sb00000000000000000000111111111111111000000000;
		13179: Delta = 44'sb11111111111111111110111111111111111000000000;
		8368: Delta = 44'sb00000000000000000010000000000000001000000000;
		10275: Delta = 44'sb11111111111111111110000000000000001000000000;
		7344: Delta = 44'sb00000000000000000001111111111111111000000000;
		9251: Delta = 44'sb11111111111111111101111111111111111000000000;
		16224: Delta = 44'sb00000000000000000100000000000000001000000000;
		2419: Delta = 44'sb11111111111111111100000000000000001000000000;
		15200: Delta = 44'sb00000000000000000011111111111111111000000000;
		1395: Delta = 44'sb11111111111111111011111111111111111000000000;
		14317: Delta = 44'sb00000000000000001000000000000000001000000000;
		4326: Delta = 44'sb11111111111111111000000000000000001000000000;
		13293: Delta = 44'sb00000000000000000111111111111111111000000000;
		3302: Delta = 44'sb11111111111111110111111111111111111000000000;
		10503: Delta = 44'sb00000000000000010000000000000000001000000000;
		8140: Delta = 44'sb11111111111111110000000000000000001000000000;
		9479: Delta = 44'sb00000000000000001111111111111111111000000000;
		7116: Delta = 44'sb11111111111111101111111111111111111000000000;
		2875: Delta = 44'sb00000000000000100000000000000000001000000000;
		15768: Delta = 44'sb11111111111111100000000000000000001000000000;
		1851: Delta = 44'sb00000000000000011111111111111111111000000000;
		14744: Delta = 44'sb11111111111111011111111111111111111000000000;
		5238: Delta = 44'sb00000000000001000000000000000000001000000000;
		13405: Delta = 44'sb11111111111111000000000000000000001000000000;
		4214: Delta = 44'sb00000000000000111111111111111111111000000000;
		12381: Delta = 44'sb11111111111110111111111111111111111000000000;
		9964: Delta = 44'sb00000000000010000000000000000000001000000000;
		8679: Delta = 44'sb11111111111110000000000000000000001000000000;
		8940: Delta = 44'sb00000000000001111111111111111111111000000000;
		7655: Delta = 44'sb11111111111101111111111111111111111000000000;
		1797: Delta = 44'sb00000000000100000000000000000000001000000000;
		16846: Delta = 44'sb11111111111100000000000000000000001000000000;
		773: Delta = 44'sb00000000000011111111111111111111111000000000;
		15822: Delta = 44'sb11111111111011111111111111111111111000000000;
		3082: Delta = 44'sb00000000001000000000000000000000001000000000;
		15561: Delta = 44'sb11111111111000000000000000000000001000000000;
		2058: Delta = 44'sb00000000000111111111111111111111111000000000;
		14537: Delta = 44'sb11111111110111111111111111111111111000000000;
		5652: Delta = 44'sb00000000010000000000000000000000001000000000;
		12991: Delta = 44'sb11111111110000000000000000000000001000000000;
		4628: Delta = 44'sb00000000001111111111111111111111111000000000;
		11967: Delta = 44'sb11111111101111111111111111111111111000000000;
		10792: Delta = 44'sb00000000100000000000000000000000001000000000;
		7851: Delta = 44'sb11111111100000000000000000000000001000000000;
		9768: Delta = 44'sb00000000011111111111111111111111111000000000;
		6827: Delta = 44'sb11111111011111111111111111111111111000000000;
		3453: Delta = 44'sb00000001000000000000000000000000001000000000;
		15190: Delta = 44'sb11111111000000000000000000000000001000000000;
		2429: Delta = 44'sb00000000111111111111111111111111111000000000;
		14166: Delta = 44'sb11111110111111111111111111111111111000000000;
		6394: Delta = 44'sb00000010000000000000000000000000001000000000;
		12249: Delta = 44'sb11111110000000000000000000000000001000000000;
		5370: Delta = 44'sb00000001111111111111111111111111111000000000;
		11225: Delta = 44'sb11111101111111111111111111111111111000000000;
		12276: Delta = 44'sb00000100000000000000000000000000001000000000;
		6367: Delta = 44'sb11111100000000000000000000000000001000000000;
		11252: Delta = 44'sb00000011111111111111111111111111111000000000;
		5343: Delta = 44'sb11111011111111111111111111111111111000000000;
		6421: Delta = 44'sb00001000000000000000000000000000001000000000;
		12222: Delta = 44'sb11111000000000000000000000000000001000000000;
		5397: Delta = 44'sb00000111111111111111111111111111111000000000;
		11198: Delta = 44'sb11110111111111111111111111111111111000000000;
		12330: Delta = 44'sb00010000000000000000000000000000001000000000;
		6313: Delta = 44'sb11110000000000000000000000000000001000000000;
		11306: Delta = 44'sb00001111111111111111111111111111111000000000;
		5289: Delta = 44'sb11101111111111111111111111111111111000000000;
		6529: Delta = 44'sb00100000000000000000000000000000001000000000;
		12114: Delta = 44'sb11100000000000000000000000000000001000000000;
		5505: Delta = 44'sb00011111111111111111111111111111111000000000;
		11090: Delta = 44'sb11011111111111111111111111111111111000000000;
		12546: Delta = 44'sb01000000000000000000000000000000001000000000;
		6097: Delta = 44'sb11000000000000000000000000000000001000000000;
		11522: Delta = 44'sb00111111111111111111111111111111111000000000;
		5073: Delta = 44'sb10111111111111111111111111111111111000000000;
		3072: Delta = 44'sb00000000000000000000000000000000110000000000;
		14547: Delta = 44'sb11111111111111111111111111111111010000000000;
		5120: Delta = 44'sb00000000000000000000000000000001010000000000;
		12499: Delta = 44'sb11111111111111111111111111111110110000000000;
		9216: Delta = 44'sb00000000000000000000000000000010010000000000;
		10451: Delta = 44'sb11111111111111111111111111111110010000000000;
		7168: Delta = 44'sb00000000000000000000000000000001110000000000;
		8403: Delta = 44'sb11111111111111111111111111111101110000000000;
		17408: Delta = 44'sb00000000000000000000000000000100010000000000;
		2259: Delta = 44'sb11111111111111111111111111111100010000000000;
		15360: Delta = 44'sb00000000000000000000000000000011110000000000;
		211: Delta = 44'sb11111111111111111111111111111011110000000000;
		16173: Delta = 44'sb00000000000000000000000000001000010000000000;
		3494: Delta = 44'sb11111111111111111111111111111000010000000000;
		14125: Delta = 44'sb00000000000000000000000000000111110000000000;
		1446: Delta = 44'sb11111111111111111111111111110111110000000000;
		13703: Delta = 44'sb00000000000000000000000000010000010000000000;
		5964: Delta = 44'sb11111111111111111111111111110000010000000000;
		11655: Delta = 44'sb00000000000000000000000000001111110000000000;
		3916: Delta = 44'sb11111111111111111111111111101111110000000000;
		8763: Delta = 44'sb00000000000000000000000000100000010000000000;
		10904: Delta = 44'sb11111111111111111111111111100000010000000000;
		6715: Delta = 44'sb00000000000000000000000000011111110000000000;
		8856: Delta = 44'sb11111111111111111111111111011111110000000000;
		16502: Delta = 44'sb00000000000000000000000001000000010000000000;
		3165: Delta = 44'sb11111111111111111111111111000000010000000000;
		14454: Delta = 44'sb00000000000000000000000000111111110000000000;
		1117: Delta = 44'sb11111111111111111111111110111111110000000000;
		14361: Delta = 44'sb00000000000000000000000010000000010000000000;
		5306: Delta = 44'sb11111111111111111111111110000000010000000000;
		12313: Delta = 44'sb00000000000000000000000001111111110000000000;
		3258: Delta = 44'sb11111111111111111111111101111111110000000000;
		10079: Delta = 44'sb00000000000000000000000100000000010000000000;
		9588: Delta = 44'sb11111111111111111111111100000000010000000000;
		8031: Delta = 44'sb00000000000000000000000011111111110000000000;
		7540: Delta = 44'sb11111111111111111111111011111111110000000000;
		1515: Delta = 44'sb00000000000000000000001000000000010000000000;
		533: Delta = 44'sb11111111111111111111111000000000010000000000;
		17086: Delta = 44'sb00000000000000000000000111111111110000000000;
		16104: Delta = 44'sb11111111111111111111110111111111110000000000;
		2006: Delta = 44'sb00000000000000000000010000000000010000000000;
		42: Delta = 44'sb11111111111111111111110000000000010000000000;
		17577: Delta = 44'sb00000000000000000000001111111111110000000000;
		15613: Delta = 44'sb11111111111111111111101111111111110000000000;
		2988: Delta = 44'sb00000000000000000000100000000000010000000000;
		16679: Delta = 44'sb11111111111111111111100000000000010000000000;
		940: Delta = 44'sb00000000000000000000011111111111110000000000;
		14631: Delta = 44'sb11111111111111111111011111111111110000000000;
		4952: Delta = 44'sb00000000000000000001000000000000010000000000;
		14715: Delta = 44'sb11111111111111111111000000000000010000000000;
		2904: Delta = 44'sb00000000000000000000111111111111110000000000;
		12667: Delta = 44'sb11111111111111111110111111111111110000000000;
		8880: Delta = 44'sb00000000000000000010000000000000010000000000;
		10787: Delta = 44'sb11111111111111111110000000000000010000000000;
		6832: Delta = 44'sb00000000000000000001111111111111110000000000;
		8739: Delta = 44'sb11111111111111111101111111111111110000000000;
		16736: Delta = 44'sb00000000000000000100000000000000010000000000;
		2931: Delta = 44'sb11111111111111111100000000000000010000000000;
		14688: Delta = 44'sb00000000000000000011111111111111110000000000;
		883: Delta = 44'sb11111111111111111011111111111111110000000000;
		14829: Delta = 44'sb00000000000000001000000000000000010000000000;
		4838: Delta = 44'sb11111111111111111000000000000000010000000000;
		12781: Delta = 44'sb00000000000000000111111111111111110000000000;
		2790: Delta = 44'sb11111111111111110111111111111111110000000000;
		11015: Delta = 44'sb00000000000000010000000000000000010000000000;
		8652: Delta = 44'sb11111111111111110000000000000000010000000000;
		8967: Delta = 44'sb00000000000000001111111111111111110000000000;
		6604: Delta = 44'sb11111111111111101111111111111111110000000000;
		3387: Delta = 44'sb00000000000000100000000000000000010000000000;
		16280: Delta = 44'sb11111111111111100000000000000000010000000000;
		1339: Delta = 44'sb00000000000000011111111111111111110000000000;
		14232: Delta = 44'sb11111111111111011111111111111111110000000000;
		5750: Delta = 44'sb00000000000001000000000000000000010000000000;
		13917: Delta = 44'sb11111111111111000000000000000000010000000000;
		3702: Delta = 44'sb00000000000000111111111111111111110000000000;
		11869: Delta = 44'sb11111111111110111111111111111111110000000000;
		10476: Delta = 44'sb00000000000010000000000000000000010000000000;
		9191: Delta = 44'sb11111111111110000000000000000000010000000000;
		8428: Delta = 44'sb00000000000001111111111111111111110000000000;
		7143: Delta = 44'sb11111111111101111111111111111111110000000000;
		2309: Delta = 44'sb00000000000100000000000000000000010000000000;
		17358: Delta = 44'sb11111111111100000000000000000000010000000000;
		261: Delta = 44'sb00000000000011111111111111111111110000000000;
		15310: Delta = 44'sb11111111111011111111111111111111110000000000;
		3594: Delta = 44'sb00000000001000000000000000000000010000000000;
		16073: Delta = 44'sb11111111111000000000000000000000010000000000;
		1546: Delta = 44'sb00000000000111111111111111111111110000000000;
		14025: Delta = 44'sb11111111110111111111111111111111110000000000;
		6164: Delta = 44'sb00000000010000000000000000000000010000000000;
		13503: Delta = 44'sb11111111110000000000000000000000010000000000;
		4116: Delta = 44'sb00000000001111111111111111111111110000000000;
		11455: Delta = 44'sb11111111101111111111111111111111110000000000;
		11304: Delta = 44'sb00000000100000000000000000000000010000000000;
		8363: Delta = 44'sb11111111100000000000000000000000010000000000;
		9256: Delta = 44'sb00000000011111111111111111111111110000000000;
		6315: Delta = 44'sb11111111011111111111111111111111110000000000;
		3965: Delta = 44'sb00000001000000000000000000000000010000000000;
		15702: Delta = 44'sb11111111000000000000000000000000010000000000;
		1917: Delta = 44'sb00000000111111111111111111111111110000000000;
		13654: Delta = 44'sb11111110111111111111111111111111110000000000;
		6906: Delta = 44'sb00000010000000000000000000000000010000000000;
		12761: Delta = 44'sb11111110000000000000000000000000010000000000;
		4858: Delta = 44'sb00000001111111111111111111111111110000000000;
		10713: Delta = 44'sb11111101111111111111111111111111110000000000;
		12788: Delta = 44'sb00000100000000000000000000000000010000000000;
		6879: Delta = 44'sb11111100000000000000000000000000010000000000;
		10740: Delta = 44'sb00000011111111111111111111111111110000000000;
		4831: Delta = 44'sb11111011111111111111111111111111110000000000;
		6933: Delta = 44'sb00001000000000000000000000000000010000000000;
		12734: Delta = 44'sb11111000000000000000000000000000010000000000;
		4885: Delta = 44'sb00000111111111111111111111111111110000000000;
		10686: Delta = 44'sb11110111111111111111111111111111110000000000;
		12842: Delta = 44'sb00010000000000000000000000000000010000000000;
		6825: Delta = 44'sb11110000000000000000000000000000010000000000;
		10794: Delta = 44'sb00001111111111111111111111111111110000000000;
		4777: Delta = 44'sb11101111111111111111111111111111110000000000;
		7041: Delta = 44'sb00100000000000000000000000000000010000000000;
		12626: Delta = 44'sb11100000000000000000000000000000010000000000;
		4993: Delta = 44'sb00011111111111111111111111111111110000000000;
		10578: Delta = 44'sb11011111111111111111111111111111110000000000;
		13058: Delta = 44'sb01000000000000000000000000000000010000000000;
		6609: Delta = 44'sb11000000000000000000000000000000010000000000;
		11010: Delta = 44'sb00111111111111111111111111111111110000000000;
		4561: Delta = 44'sb10111111111111111111111111111111110000000000;
		6144: Delta = 44'sb00000000000000000000000000000001100000000000;
		11475: Delta = 44'sb11111111111111111111111111111110100000000000;
		10240: Delta = 44'sb00000000000000000000000000000010100000000000;
		7379: Delta = 44'sb11111111111111111111111111111101100000000000;
		813: Delta = 44'sb00000000000000000000000000000100100000000000;
		3283: Delta = 44'sb11111111111111111111111111111100100000000000;
		14336: Delta = 44'sb00000000000000000000000000000011100000000000;
		16806: Delta = 44'sb11111111111111111111111111111011100000000000;
		17197: Delta = 44'sb00000000000000000000000000001000100000000000;
		4518: Delta = 44'sb11111111111111111111111111111000100000000000;
		13101: Delta = 44'sb00000000000000000000000000000111100000000000;
		422: Delta = 44'sb11111111111111111111111111110111100000000000;
		14727: Delta = 44'sb00000000000000000000000000010000100000000000;
		6988: Delta = 44'sb11111111111111111111111111110000100000000000;
		10631: Delta = 44'sb00000000000000000000000000001111100000000000;
		2892: Delta = 44'sb11111111111111111111111111101111100000000000;
		9787: Delta = 44'sb00000000000000000000000000100000100000000000;
		11928: Delta = 44'sb11111111111111111111111111100000100000000000;
		5691: Delta = 44'sb00000000000000000000000000011111100000000000;
		7832: Delta = 44'sb11111111111111111111111111011111100000000000;
		17526: Delta = 44'sb00000000000000000000000001000000100000000000;
		4189: Delta = 44'sb11111111111111111111111111000000100000000000;
		13430: Delta = 44'sb00000000000000000000000000111111100000000000;
		93: Delta = 44'sb11111111111111111111111110111111100000000000;
		15385: Delta = 44'sb00000000000000000000000010000000100000000000;
		6330: Delta = 44'sb11111111111111111111111110000000100000000000;
		11289: Delta = 44'sb00000000000000000000000001111111100000000000;
		2234: Delta = 44'sb11111111111111111111111101111111100000000000;
		11103: Delta = 44'sb00000000000000000000000100000000100000000000;
		10612: Delta = 44'sb11111111111111111111111100000000100000000000;
		7007: Delta = 44'sb00000000000000000000000011111111100000000000;
		6516: Delta = 44'sb11111111111111111111111011111111100000000000;
		2539: Delta = 44'sb00000000000000000000001000000000100000000000;
		1557: Delta = 44'sb11111111111111111111111000000000100000000000;
		16062: Delta = 44'sb00000000000000000000000111111111100000000000;
		15080: Delta = 44'sb11111111111111111111110111111111100000000000;
		3030: Delta = 44'sb00000000000000000000010000000000100000000000;
		1066: Delta = 44'sb11111111111111111111110000000000100000000000;
		16553: Delta = 44'sb00000000000000000000001111111111100000000000;
		14589: Delta = 44'sb11111111111111111111101111111111100000000000;
		4012: Delta = 44'sb00000000000000000000100000000000100000000000;
		84: Delta = 44'sb11111111111111111111100000000000100000000000;
		17535: Delta = 44'sb00000000000000000000011111111111100000000000;
		13607: Delta = 44'sb11111111111111111111011111111111100000000000;
		5976: Delta = 44'sb00000000000000000001000000000000100000000000;
		15739: Delta = 44'sb11111111111111111111000000000000100000000000;
		1880: Delta = 44'sb00000000000000000000111111111111100000000000;
		11643: Delta = 44'sb11111111111111111110111111111111100000000000;
		9904: Delta = 44'sb00000000000000000010000000000000100000000000;
		11811: Delta = 44'sb11111111111111111110000000000000100000000000;
		5808: Delta = 44'sb00000000000000000001111111111111100000000000;
		7715: Delta = 44'sb11111111111111111101111111111111100000000000;
		141: Delta = 44'sb00000000000000000100000000000000100000000000;
		3955: Delta = 44'sb11111111111111111100000000000000100000000000;
		13664: Delta = 44'sb00000000000000000011111111111111100000000000;
		17478: Delta = 44'sb11111111111111111011111111111111100000000000;
		15853: Delta = 44'sb00000000000000001000000000000000100000000000;
		5862: Delta = 44'sb11111111111111111000000000000000100000000000;
		11757: Delta = 44'sb00000000000000000111111111111111100000000000;
		1766: Delta = 44'sb11111111111111110111111111111111100000000000;
		12039: Delta = 44'sb00000000000000010000000000000000100000000000;
		9676: Delta = 44'sb11111111111111110000000000000000100000000000;
		7943: Delta = 44'sb00000000000000001111111111111111100000000000;
		5580: Delta = 44'sb11111111111111101111111111111111100000000000;
		4411: Delta = 44'sb00000000000000100000000000000000100000000000;
		17304: Delta = 44'sb11111111111111100000000000000000100000000000;
		315: Delta = 44'sb00000000000000011111111111111111100000000000;
		13208: Delta = 44'sb11111111111111011111111111111111100000000000;
		6774: Delta = 44'sb00000000000001000000000000000000100000000000;
		14941: Delta = 44'sb11111111111111000000000000000000100000000000;
		2678: Delta = 44'sb00000000000000111111111111111111100000000000;
		10845: Delta = 44'sb11111111111110111111111111111111100000000000;
		11500: Delta = 44'sb00000000000010000000000000000000100000000000;
		10215: Delta = 44'sb11111111111110000000000000000000100000000000;
		7404: Delta = 44'sb00000000000001111111111111111111100000000000;
		6119: Delta = 44'sb11111111111101111111111111111111100000000000;
		3333: Delta = 44'sb00000000000100000000000000000000100000000000;
		763: Delta = 44'sb11111111111100000000000000000000100000000000;
		16856: Delta = 44'sb00000000000011111111111111111111100000000000;
		14286: Delta = 44'sb11111111111011111111111111111111100000000000;
		4618: Delta = 44'sb00000000001000000000000000000000100000000000;
		17097: Delta = 44'sb11111111111000000000000000000000100000000000;
		522: Delta = 44'sb00000000000111111111111111111111100000000000;
		13001: Delta = 44'sb11111111110111111111111111111111100000000000;
		7188: Delta = 44'sb00000000010000000000000000000000100000000000;
		14527: Delta = 44'sb11111111110000000000000000000000100000000000;
		3092: Delta = 44'sb00000000001111111111111111111111100000000000;
		10431: Delta = 44'sb11111111101111111111111111111111100000000000;
		12328: Delta = 44'sb00000000100000000000000000000000100000000000;
		9387: Delta = 44'sb11111111100000000000000000000000100000000000;
		8232: Delta = 44'sb00000000011111111111111111111111100000000000;
		5291: Delta = 44'sb11111111011111111111111111111111100000000000;
		4989: Delta = 44'sb00000001000000000000000000000000100000000000;
		16726: Delta = 44'sb11111111000000000000000000000000100000000000;
		893: Delta = 44'sb00000000111111111111111111111111100000000000;
		12630: Delta = 44'sb11111110111111111111111111111111100000000000;
		7930: Delta = 44'sb00000010000000000000000000000000100000000000;
		13785: Delta = 44'sb11111110000000000000000000000000100000000000;
		3834: Delta = 44'sb00000001111111111111111111111111100000000000;
		9689: Delta = 44'sb11111101111111111111111111111111100000000000;
		13812: Delta = 44'sb00000100000000000000000000000000100000000000;
		7903: Delta = 44'sb11111100000000000000000000000000100000000000;
		9716: Delta = 44'sb00000011111111111111111111111111100000000000;
		3807: Delta = 44'sb11111011111111111111111111111111100000000000;
		7957: Delta = 44'sb00001000000000000000000000000000100000000000;
		13758: Delta = 44'sb11111000000000000000000000000000100000000000;
		3861: Delta = 44'sb00000111111111111111111111111111100000000000;
		9662: Delta = 44'sb11110111111111111111111111111111100000000000;
		13866: Delta = 44'sb00010000000000000000000000000000100000000000;
		7849: Delta = 44'sb11110000000000000000000000000000100000000000;
		9770: Delta = 44'sb00001111111111111111111111111111100000000000;
		3753: Delta = 44'sb11101111111111111111111111111111100000000000;
		8065: Delta = 44'sb00100000000000000000000000000000100000000000;
		13650: Delta = 44'sb11100000000000000000000000000000100000000000;
		3969: Delta = 44'sb00011111111111111111111111111111100000000000;
		9554: Delta = 44'sb11011111111111111111111111111111100000000000;
		14082: Delta = 44'sb01000000000000000000000000000000100000000000;
		7633: Delta = 44'sb11000000000000000000000000000000100000000000;
		9986: Delta = 44'sb00111111111111111111111111111111100000000000;
		3537: Delta = 44'sb10111111111111111111111111111111100000000000;
		12288: Delta = 44'sb00000000000000000000000000000011000000000000;
		5331: Delta = 44'sb11111111111111111111111111111101000000000000;
		2861: Delta = 44'sb00000000000000000000000000000101000000000000;
		14758: Delta = 44'sb11111111111111111111111111111011000000000000;
		1626: Delta = 44'sb00000000000000000000000000001001000000000000;
		6566: Delta = 44'sb11111111111111111111111111111001000000000000;
		11053: Delta = 44'sb00000000000000000000000000000111000000000000;
		15993: Delta = 44'sb11111111111111111111111111110111000000000000;
		16775: Delta = 44'sb00000000000000000000000000010001000000000000;
		9036: Delta = 44'sb11111111111111111111111111110001000000000000;
		8583: Delta = 44'sb00000000000000000000000000001111000000000000;
		844: Delta = 44'sb11111111111111111111111111101111000000000000;
		11835: Delta = 44'sb00000000000000000000000000100001000000000000;
		13976: Delta = 44'sb11111111111111111111111111100001000000000000;
		3643: Delta = 44'sb00000000000000000000000000011111000000000000;
		5784: Delta = 44'sb11111111111111111111111111011111000000000000;
		1955: Delta = 44'sb00000000000000000000000001000001000000000000;
		6237: Delta = 44'sb11111111111111111111111111000001000000000000;
		11382: Delta = 44'sb00000000000000000000000000111111000000000000;
		15664: Delta = 44'sb11111111111111111111111110111111000000000000;
		17433: Delta = 44'sb00000000000000000000000010000001000000000000;
		8378: Delta = 44'sb11111111111111111111111110000001000000000000;
		9241: Delta = 44'sb00000000000000000000000001111111000000000000;
		186: Delta = 44'sb11111111111111111111111101111111000000000000;
		13151: Delta = 44'sb00000000000000000000000100000001000000000000;
		12660: Delta = 44'sb11111111111111111111111100000001000000000000;
		4959: Delta = 44'sb00000000000000000000000011111111000000000000;
		4468: Delta = 44'sb11111111111111111111111011111111000000000000;
		4587: Delta = 44'sb00000000000000000000001000000001000000000000;
		3605: Delta = 44'sb11111111111111111111111000000001000000000000;
		14014: Delta = 44'sb00000000000000000000000111111111000000000000;
		13032: Delta = 44'sb11111111111111111111110111111111000000000000;
		5078: Delta = 44'sb00000000000000000000010000000001000000000000;
		3114: Delta = 44'sb11111111111111111111110000000001000000000000;
		14505: Delta = 44'sb00000000000000000000001111111111000000000000;
		12541: Delta = 44'sb11111111111111111111101111111111000000000000;
		6060: Delta = 44'sb00000000000000000000100000000001000000000000;
		2132: Delta = 44'sb11111111111111111111100000000001000000000000;
		15487: Delta = 44'sb00000000000000000000011111111111000000000000;
		11559: Delta = 44'sb11111111111111111111011111111111000000000000;
		8024: Delta = 44'sb00000000000000000001000000000001000000000000;
		168: Delta = 44'sb11111111111111111111000000000001000000000000;
		17451: Delta = 44'sb00000000000000000000111111111111000000000000;
		9595: Delta = 44'sb11111111111111111110111111111111000000000000;
		11952: Delta = 44'sb00000000000000000010000000000001000000000000;
		13859: Delta = 44'sb11111111111111111110000000000001000000000000;
		3760: Delta = 44'sb00000000000000000001111111111111000000000000;
		5667: Delta = 44'sb11111111111111111101111111111111000000000000;
		2189: Delta = 44'sb00000000000000000100000000000001000000000000;
		6003: Delta = 44'sb11111111111111111100000000000001000000000000;
		11616: Delta = 44'sb00000000000000000011111111111111000000000000;
		15430: Delta = 44'sb11111111111111111011111111111111000000000000;
		282: Delta = 44'sb00000000000000001000000000000001000000000000;
		7910: Delta = 44'sb11111111111111111000000000000001000000000000;
		9709: Delta = 44'sb00000000000000000111111111111111000000000000;
		17337: Delta = 44'sb11111111111111110111111111111111000000000000;
		14087: Delta = 44'sb00000000000000010000000000000001000000000000;
		11724: Delta = 44'sb11111111111111110000000000000001000000000000;
		5895: Delta = 44'sb00000000000000001111111111111111000000000000;
		3532: Delta = 44'sb11111111111111101111111111111111000000000000;
		6459: Delta = 44'sb00000000000000100000000000000001000000000000;
		1733: Delta = 44'sb11111111111111100000000000000001000000000000;
		15886: Delta = 44'sb00000000000000011111111111111111000000000000;
		11160: Delta = 44'sb11111111111111011111111111111111000000000000;
		8822: Delta = 44'sb00000000000001000000000000000001000000000000;
		16989: Delta = 44'sb11111111111111000000000000000001000000000000;
		630: Delta = 44'sb00000000000000111111111111111111000000000000;
		8797: Delta = 44'sb11111111111110111111111111111111000000000000;
		13548: Delta = 44'sb00000000000010000000000000000001000000000000;
		12263: Delta = 44'sb11111111111110000000000000000001000000000000;
		5356: Delta = 44'sb00000000000001111111111111111111000000000000;
		4071: Delta = 44'sb11111111111101111111111111111111000000000000;
		5381: Delta = 44'sb00000000000100000000000000000001000000000000;
		2811: Delta = 44'sb11111111111100000000000000000001000000000000;
		14808: Delta = 44'sb00000000000011111111111111111111000000000000;
		12238: Delta = 44'sb11111111111011111111111111111111000000000000;
		6666: Delta = 44'sb00000000001000000000000000000001000000000000;
		1526: Delta = 44'sb11111111111000000000000000000001000000000000;
		16093: Delta = 44'sb00000000000111111111111111111111000000000000;
		10953: Delta = 44'sb11111111110111111111111111111111000000000000;
		9236: Delta = 44'sb00000000010000000000000000000001000000000000;
		16575: Delta = 44'sb11111111110000000000000000000001000000000000;
		1044: Delta = 44'sb00000000001111111111111111111111000000000000;
		8383: Delta = 44'sb11111111101111111111111111111111000000000000;
		14376: Delta = 44'sb00000000100000000000000000000001000000000000;
		11435: Delta = 44'sb11111111100000000000000000000001000000000000;
		6184: Delta = 44'sb00000000011111111111111111111111000000000000;
		3243: Delta = 44'sb11111111011111111111111111111111000000000000;
		7037: Delta = 44'sb00000001000000000000000000000001000000000000;
		1155: Delta = 44'sb11111111000000000000000000000001000000000000;
		16464: Delta = 44'sb00000000111111111111111111111111000000000000;
		10582: Delta = 44'sb11111110111111111111111111111111000000000000;
		9978: Delta = 44'sb00000010000000000000000000000001000000000000;
		15833: Delta = 44'sb11111110000000000000000000000001000000000000;
		1786: Delta = 44'sb00000001111111111111111111111111000000000000;
		7641: Delta = 44'sb11111101111111111111111111111111000000000000;
		15860: Delta = 44'sb00000100000000000000000000000001000000000000;
		9951: Delta = 44'sb11111100000000000000000000000001000000000000;
		7668: Delta = 44'sb00000011111111111111111111111111000000000000;
		1759: Delta = 44'sb11111011111111111111111111111111000000000000;
		10005: Delta = 44'sb00001000000000000000000000000001000000000000;
		15806: Delta = 44'sb11111000000000000000000000000001000000000000;
		1813: Delta = 44'sb00000111111111111111111111111111000000000000;
		7614: Delta = 44'sb11110111111111111111111111111111000000000000;
		15914: Delta = 44'sb00010000000000000000000000000001000000000000;
		9897: Delta = 44'sb11110000000000000000000000000001000000000000;
		7722: Delta = 44'sb00001111111111111111111111111111000000000000;
		1705: Delta = 44'sb11101111111111111111111111111111000000000000;
		10113: Delta = 44'sb00100000000000000000000000000001000000000000;
		15698: Delta = 44'sb11100000000000000000000000000001000000000000;
		1921: Delta = 44'sb00011111111111111111111111111111000000000000;
		7506: Delta = 44'sb11011111111111111111111111111111000000000000;
		16130: Delta = 44'sb01000000000000000000000000000001000000000000;
		9681: Delta = 44'sb11000000000000000000000000000001000000000000;
		7938: Delta = 44'sb00111111111111111111111111111111000000000000;
		1489: Delta = 44'sb10111111111111111111111111111111000000000000;
		6957: Delta = 44'sb00000000000000000000000000000110000000000000;
		10662: Delta = 44'sb11111111111111111111111111111010000000000000;
		5722: Delta = 44'sb00000000000000000000000000001010000000000000;
		11897: Delta = 44'sb11111111111111111111111111110110000000000000;
		3252: Delta = 44'sb00000000000000000000000000010010000000000000;
		13132: Delta = 44'sb11111111111111111111111111110010000000000000;
		4487: Delta = 44'sb00000000000000000000000000001110000000000000;
		14367: Delta = 44'sb11111111111111111111111111101110000000000000;
		15931: Delta = 44'sb00000000000000000000000000100010000000000000;
		453: Delta = 44'sb11111111111111111111111111100010000000000000;
		17166: Delta = 44'sb00000000000000000000000000011110000000000000;
		1688: Delta = 44'sb11111111111111111111111111011110000000000000;
		6051: Delta = 44'sb00000000000000000000000001000010000000000000;
		10333: Delta = 44'sb11111111111111111111111111000010000000000000;
		7286: Delta = 44'sb00000000000000000000000000111110000000000000;
		11568: Delta = 44'sb11111111111111111111111110111110000000000000;
		3910: Delta = 44'sb00000000000000000000000010000010000000000000;
		12474: Delta = 44'sb11111111111111111111111110000010000000000000;
		5145: Delta = 44'sb00000000000000000000000001111110000000000000;
		13709: Delta = 44'sb11111111111111111111111101111110000000000000;
		17247: Delta = 44'sb00000000000000000000000100000010000000000000;
		16756: Delta = 44'sb11111111111111111111111100000010000000000000;
		863: Delta = 44'sb00000000000000000000000011111110000000000000;
		372: Delta = 44'sb11111111111111111111111011111110000000000000;
		8683: Delta = 44'sb00000000000000000000001000000010000000000000;
		7701: Delta = 44'sb11111111111111111111111000000010000000000000;
		9918: Delta = 44'sb00000000000000000000000111111110000000000000;
		8936: Delta = 44'sb11111111111111111111110111111110000000000000;
		9174: Delta = 44'sb00000000000000000000010000000010000000000000;
		7210: Delta = 44'sb11111111111111111111110000000010000000000000;
		10409: Delta = 44'sb00000000000000000000001111111110000000000000;
		8445: Delta = 44'sb11111111111111111111101111111110000000000000;
		10156: Delta = 44'sb00000000000000000000100000000010000000000000;
		6228: Delta = 44'sb11111111111111111111100000000010000000000000;
		11391: Delta = 44'sb00000000000000000000011111111110000000000000;
		7463: Delta = 44'sb11111111111111111111011111111110000000000000;
		12120: Delta = 44'sb00000000000000000001000000000010000000000000;
		4264: Delta = 44'sb11111111111111111111000000000010000000000000;
		13355: Delta = 44'sb00000000000000000000111111111110000000000000;
		5499: Delta = 44'sb11111111111111111110111111111110000000000000;
		16048: Delta = 44'sb00000000000000000010000000000010000000000000;
		336: Delta = 44'sb11111111111111111110000000000010000000000000;
		17283: Delta = 44'sb00000000000000000001111111111110000000000000;
		1571: Delta = 44'sb11111111111111111101111111111110000000000000;
		6285: Delta = 44'sb00000000000000000100000000000010000000000000;
		10099: Delta = 44'sb11111111111111111100000000000010000000000000;
		7520: Delta = 44'sb00000000000000000011111111111110000000000000;
		11334: Delta = 44'sb11111111111111111011111111111110000000000000;
		4378: Delta = 44'sb00000000000000001000000000000010000000000000;
		12006: Delta = 44'sb11111111111111111000000000000010000000000000;
		5613: Delta = 44'sb00000000000000000111111111111110000000000000;
		13241: Delta = 44'sb11111111111111110111111111111110000000000000;
		564: Delta = 44'sb00000000000000010000000000000010000000000000;
		15820: Delta = 44'sb11111111111111110000000000000010000000000000;
		1799: Delta = 44'sb00000000000000001111111111111110000000000000;
		17055: Delta = 44'sb11111111111111101111111111111110000000000000;
		10555: Delta = 44'sb00000000000000100000000000000010000000000000;
		5829: Delta = 44'sb11111111111111100000000000000010000000000000;
		11790: Delta = 44'sb00000000000000011111111111111110000000000000;
		7064: Delta = 44'sb11111111111111011111111111111110000000000000;
		12918: Delta = 44'sb00000000000001000000000000000010000000000000;
		3466: Delta = 44'sb11111111111111000000000000000010000000000000;
		14153: Delta = 44'sb00000000000000111111111111111110000000000000;
		4701: Delta = 44'sb11111111111110111111111111111110000000000000;
		25: Delta = 44'sb00000000000010000000000000000010000000000000;
		16359: Delta = 44'sb11111111111110000000000000000010000000000000;
		1260: Delta = 44'sb00000000000001111111111111111110000000000000;
		17594: Delta = 44'sb11111111111101111111111111111110000000000000;
		9477: Delta = 44'sb00000000000100000000000000000010000000000000;
		6907: Delta = 44'sb11111111111100000000000000000010000000000000;
		10712: Delta = 44'sb00000000000011111111111111111110000000000000;
		8142: Delta = 44'sb11111111111011111111111111111110000000000000;
		10762: Delta = 44'sb00000000001000000000000000000010000000000000;
		5622: Delta = 44'sb11111111111000000000000000000010000000000000;
		11997: Delta = 44'sb00000000000111111111111111111110000000000000;
		6857: Delta = 44'sb11111111110111111111111111111110000000000000;
		13332: Delta = 44'sb00000000010000000000000000000010000000000000;
		3052: Delta = 44'sb11111111110000000000000000000010000000000000;
		14567: Delta = 44'sb00000000001111111111111111111110000000000000;
		4287: Delta = 44'sb11111111101111111111111111111110000000000000;
		853: Delta = 44'sb00000000100000000000000000000010000000000000;
		15531: Delta = 44'sb11111111100000000000000000000010000000000000;
		2088: Delta = 44'sb00000000011111111111111111111110000000000000;
		16766: Delta = 44'sb11111111011111111111111111111110000000000000;
		11133: Delta = 44'sb00000001000000000000000000000010000000000000;
		5251: Delta = 44'sb11111111000000000000000000000010000000000000;
		12368: Delta = 44'sb00000000111111111111111111111110000000000000;
		6486: Delta = 44'sb11111110111111111111111111111110000000000000;
		14074: Delta = 44'sb00000010000000000000000000000010000000000000;
		2310: Delta = 44'sb11111110000000000000000000000010000000000000;
		15309: Delta = 44'sb00000001111111111111111111111110000000000000;
		3545: Delta = 44'sb11111101111111111111111111111110000000000000;
		2337: Delta = 44'sb00000100000000000000000000000010000000000000;
		14047: Delta = 44'sb11111100000000000000000000000010000000000000;
		3572: Delta = 44'sb00000011111111111111111111111110000000000000;
		15282: Delta = 44'sb11111011111111111111111111111110000000000000;
		14101: Delta = 44'sb00001000000000000000000000000010000000000000;
		2283: Delta = 44'sb11111000000000000000000000000010000000000000;
		15336: Delta = 44'sb00000111111111111111111111111110000000000000;
		3518: Delta = 44'sb11110111111111111111111111111110000000000000;
		2391: Delta = 44'sb00010000000000000000000000000010000000000000;
		13993: Delta = 44'sb11110000000000000000000000000010000000000000;
		3626: Delta = 44'sb00001111111111111111111111111110000000000000;
		15228: Delta = 44'sb11101111111111111111111111111110000000000000;
		14209: Delta = 44'sb00100000000000000000000000000010000000000000;
		2175: Delta = 44'sb11100000000000000000000000000010000000000000;
		15444: Delta = 44'sb00011111111111111111111111111110000000000000;
		3410: Delta = 44'sb11011111111111111111111111111110000000000000;
		2607: Delta = 44'sb01000000000000000000000000000010000000000000;
		13777: Delta = 44'sb11000000000000000000000000000010000000000000;
		3842: Delta = 44'sb00111111111111111111111111111110000000000000;
		15012: Delta = 44'sb10111111111111111111111111111110000000000000;
		13914: Delta = 44'sb00000000000000000000000000001100000000000000;
		3705: Delta = 44'sb11111111111111111111111111110100000000000000;
		11444: Delta = 44'sb00000000000000000000000000010100000000000000;
		6175: Delta = 44'sb11111111111111111111111111101100000000000000;
		6504: Delta = 44'sb00000000000000000000000000100100000000000000;
		8645: Delta = 44'sb11111111111111111111111111100100000000000000;
		8974: Delta = 44'sb00000000000000000000000000011100000000000000;
		11115: Delta = 44'sb11111111111111111111111111011100000000000000;
		14243: Delta = 44'sb00000000000000000000000001000100000000000000;
		906: Delta = 44'sb11111111111111111111111111000100000000000000;
		16713: Delta = 44'sb00000000000000000000000000111100000000000000;
		3376: Delta = 44'sb11111111111111111111111110111100000000000000;
		12102: Delta = 44'sb00000000000000000000000010000100000000000000;
		3047: Delta = 44'sb11111111111111111111111110000100000000000000;
		14572: Delta = 44'sb00000000000000000000000001111100000000000000;
		5517: Delta = 44'sb11111111111111111111111101111100000000000000;
		7820: Delta = 44'sb00000000000000000000000100000100000000000000;
		7329: Delta = 44'sb11111111111111111111111100000100000000000000;
		10290: Delta = 44'sb00000000000000000000000011111100000000000000;
		9799: Delta = 44'sb11111111111111111111111011111100000000000000;
		16875: Delta = 44'sb00000000000000000000001000000100000000000000;
		15893: Delta = 44'sb11111111111111111111111000000100000000000000;
		1726: Delta = 44'sb00000000000000000000000111111100000000000000;
		744: Delta = 44'sb11111111111111111111110111111100000000000000;
		17366: Delta = 44'sb00000000000000000000010000000100000000000000;
		15402: Delta = 44'sb11111111111111111111110000000100000000000000;
		2217: Delta = 44'sb00000000000000000000001111111100000000000000;
		253: Delta = 44'sb11111111111111111111101111111100000000000000;
		729: Delta = 44'sb00000000000000000000100000000100000000000000;
		14420: Delta = 44'sb11111111111111111111100000000100000000000000;
		3199: Delta = 44'sb00000000000000000000011111111100000000000000;
		16890: Delta = 44'sb11111111111111111111011111111100000000000000;
		2693: Delta = 44'sb00000000000000000001000000000100000000000000;
		12456: Delta = 44'sb11111111111111111111000000000100000000000000;
		5163: Delta = 44'sb00000000000000000000111111111100000000000000;
		14926: Delta = 44'sb11111111111111111110111111111100000000000000;
		6621: Delta = 44'sb00000000000000000010000000000100000000000000;
		8528: Delta = 44'sb11111111111111111110000000000100000000000000;
		9091: Delta = 44'sb00000000000000000001111111111100000000000000;
		10998: Delta = 44'sb11111111111111111101111111111100000000000000;
		14477: Delta = 44'sb00000000000000000100000000000100000000000000;
		672: Delta = 44'sb11111111111111111100000000000100000000000000;
		16947: Delta = 44'sb00000000000000000011111111111100000000000000;
		3142: Delta = 44'sb11111111111111111011111111111100000000000000;
		12570: Delta = 44'sb00000000000000001000000000000100000000000000;
		2579: Delta = 44'sb11111111111111111000000000000100000000000000;
		15040: Delta = 44'sb00000000000000000111111111111100000000000000;
		5049: Delta = 44'sb11111111111111110111111111111100000000000000;
		8756: Delta = 44'sb00000000000000010000000000000100000000000000;
		6393: Delta = 44'sb11111111111111110000000000000100000000000000;
		11226: Delta = 44'sb00000000000000001111111111111100000000000000;
		8863: Delta = 44'sb11111111111111101111111111111100000000000000;
		1128: Delta = 44'sb00000000000000100000000000000100000000000000;
		14021: Delta = 44'sb11111111111111100000000000000100000000000000;
		3598: Delta = 44'sb00000000000000011111111111111100000000000000;
		16491: Delta = 44'sb11111111111111011111111111111100000000000000;
		3491: Delta = 44'sb00000000000001000000000000000100000000000000;
		11658: Delta = 44'sb11111111111111000000000000000100000000000000;
		5961: Delta = 44'sb00000000000000111111111111111100000000000000;
		14128: Delta = 44'sb11111111111110111111111111111100000000000000;
		8217: Delta = 44'sb00000000000010000000000000000100000000000000;
		6932: Delta = 44'sb11111111111110000000000000000100000000000000;
		10687: Delta = 44'sb00000000000001111111111111111100000000000000;
		9402: Delta = 44'sb11111111111101111111111111111100000000000000;
		50: Delta = 44'sb00000000000100000000000000000100000000000000;
		15099: Delta = 44'sb11111111111100000000000000000100000000000000;
		2520: Delta = 44'sb00000000000011111111111111111100000000000000;
		17569: Delta = 44'sb11111111111011111111111111111100000000000000;
		1335: Delta = 44'sb00000000001000000000000000000100000000000000;
		13814: Delta = 44'sb11111111111000000000000000000100000000000000;
		3805: Delta = 44'sb00000000000111111111111111111100000000000000;
		16284: Delta = 44'sb11111111110111111111111111111100000000000000;
		3905: Delta = 44'sb00000000010000000000000000000100000000000000;
		11244: Delta = 44'sb11111111110000000000000000000100000000000000;
		6375: Delta = 44'sb00000000001111111111111111111100000000000000;
		13714: Delta = 44'sb11111111101111111111111111111100000000000000;
		9045: Delta = 44'sb00000000100000000000000000000100000000000000;
		6104: Delta = 44'sb11111111100000000000000000000100000000000000;
		11515: Delta = 44'sb00000000011111111111111111111100000000000000;
		8574: Delta = 44'sb11111111011111111111111111111100000000000000;
		1706: Delta = 44'sb00000001000000000000000000000100000000000000;
		13443: Delta = 44'sb11111111000000000000000000000100000000000000;
		4176: Delta = 44'sb00000000111111111111111111111100000000000000;
		15913: Delta = 44'sb11111110111111111111111111111100000000000000;
		4647: Delta = 44'sb00000010000000000000000000000100000000000000;
		10502: Delta = 44'sb11111110000000000000000000000100000000000000;
		7117: Delta = 44'sb00000001111111111111111111111100000000000000;
		12972: Delta = 44'sb11111101111111111111111111111100000000000000;
		10529: Delta = 44'sb00000100000000000000000000000100000000000000;
		4620: Delta = 44'sb11111100000000000000000000000100000000000000;
		12999: Delta = 44'sb00000011111111111111111111111100000000000000;
		7090: Delta = 44'sb11111011111111111111111111111100000000000000;
		4674: Delta = 44'sb00001000000000000000000000000100000000000000;
		10475: Delta = 44'sb11111000000000000000000000000100000000000000;
		7144: Delta = 44'sb00000111111111111111111111111100000000000000;
		12945: Delta = 44'sb11110111111111111111111111111100000000000000;
		10583: Delta = 44'sb00010000000000000000000000000100000000000000;
		4566: Delta = 44'sb11110000000000000000000000000100000000000000;
		13053: Delta = 44'sb00001111111111111111111111111100000000000000;
		7036: Delta = 44'sb11101111111111111111111111111100000000000000;
		4782: Delta = 44'sb00100000000000000000000000000100000000000000;
		10367: Delta = 44'sb11100000000000000000000000000100000000000000;
		7252: Delta = 44'sb00011111111111111111111111111100000000000000;
		12837: Delta = 44'sb11011111111111111111111111111100000000000000;
		10799: Delta = 44'sb01000000000000000000000000000100000000000000;
		4350: Delta = 44'sb11000000000000000000000000000100000000000000;
		13269: Delta = 44'sb00111111111111111111111111111100000000000000;
		6820: Delta = 44'sb10111111111111111111111111111100000000000000;
		10209: Delta = 44'sb00000000000000000000000000011000000000000000;
		7410: Delta = 44'sb11111111111111111111111111101000000000000000;
		5269: Delta = 44'sb00000000000000000000000000101000000000000000;
		12350: Delta = 44'sb11111111111111111111111111011000000000000000;
		13008: Delta = 44'sb00000000000000000000000001001000000000000000;
		17290: Delta = 44'sb11111111111111111111111111001000000000000000;
		329: Delta = 44'sb00000000000000000000000000111000000000000000;
		4611: Delta = 44'sb11111111111111111111111110111000000000000000;
		10867: Delta = 44'sb00000000000000000000000010001000000000000000;
		1812: Delta = 44'sb11111111111111111111111110001000000000000000;
		15807: Delta = 44'sb00000000000000000000000001111000000000000000;
		6752: Delta = 44'sb11111111111111111111111101111000000000000000;
		6585: Delta = 44'sb00000000000000000000000100001000000000000000;
		6094: Delta = 44'sb11111111111111111111111100001000000000000000;
		11525: Delta = 44'sb00000000000000000000000011111000000000000000;
		11034: Delta = 44'sb11111111111111111111111011111000000000000000;
		15640: Delta = 44'sb00000000000000000000001000001000000000000000;
		14658: Delta = 44'sb11111111111111111111111000001000000000000000;
		2961: Delta = 44'sb00000000000000000000000111111000000000000000;
		1979: Delta = 44'sb11111111111111111111110111111000000000000000;
		16131: Delta = 44'sb00000000000000000000010000001000000000000000;
		14167: Delta = 44'sb11111111111111111111110000001000000000000000;
		3452: Delta = 44'sb00000000000000000000001111111000000000000000;
		1488: Delta = 44'sb11111111111111111111101111111000000000000000;
		17113: Delta = 44'sb00000000000000000000100000001000000000000000;
		13185: Delta = 44'sb11111111111111111111100000001000000000000000;
		4434: Delta = 44'sb00000000000000000000011111111000000000000000;
		506: Delta = 44'sb11111111111111111111011111111000000000000000;
		1458: Delta = 44'sb00000000000000000001000000001000000000000000;
		11221: Delta = 44'sb11111111111111111111000000001000000000000000;
		6398: Delta = 44'sb00000000000000000000111111111000000000000000;
		16161: Delta = 44'sb11111111111111111110111111111000000000000000;
		5386: Delta = 44'sb00000000000000000010000000001000000000000000;
		7293: Delta = 44'sb11111111111111111110000000001000000000000000;
		10326: Delta = 44'sb00000000000000000001111111111000000000000000;
		12233: Delta = 44'sb11111111111111111101111111111000000000000000;
		13242: Delta = 44'sb00000000000000000100000000001000000000000000;
		17056: Delta = 44'sb11111111111111111100000000001000000000000000;
		563: Delta = 44'sb00000000000000000011111111111000000000000000;
		4377: Delta = 44'sb11111111111111111011111111111000000000000000;
		11335: Delta = 44'sb00000000000000001000000000001000000000000000;
		1344: Delta = 44'sb11111111111111111000000000001000000000000000;
		16275: Delta = 44'sb00000000000000000111111111111000000000000000;
		6284: Delta = 44'sb11111111111111110111111111111000000000000000;
		7521: Delta = 44'sb00000000000000010000000000001000000000000000;
		5158: Delta = 44'sb11111111111111110000000000001000000000000000;
		12461: Delta = 44'sb00000000000000001111111111111000000000000000;
		10098: Delta = 44'sb11111111111111101111111111111000000000000000;
		17512: Delta = 44'sb00000000000000100000000000001000000000000000;
		12786: Delta = 44'sb11111111111111100000000000001000000000000000;
		4833: Delta = 44'sb00000000000000011111111111111000000000000000;
		107: Delta = 44'sb11111111111111011111111111111000000000000000;
		2256: Delta = 44'sb00000000000001000000000000001000000000000000;
		10423: Delta = 44'sb11111111111111000000000000001000000000000000;
		7196: Delta = 44'sb00000000000000111111111111111000000000000000;
		15363: Delta = 44'sb11111111111110111111111111111000000000000000;
		6982: Delta = 44'sb00000000000010000000000000001000000000000000;
		5697: Delta = 44'sb11111111111110000000000000001000000000000000;
		11922: Delta = 44'sb00000000000001111111111111111000000000000000;
		10637: Delta = 44'sb11111111111101111111111111111000000000000000;
		16434: Delta = 44'sb00000000000100000000000000001000000000000000;
		13864: Delta = 44'sb11111111111100000000000000001000000000000000;
		3755: Delta = 44'sb00000000000011111111111111111000000000000000;
		1185: Delta = 44'sb11111111111011111111111111111000000000000000;
		100: Delta = 44'sb00000000001000000000000000001000000000000000;
		12579: Delta = 44'sb11111111111000000000000000001000000000000000;
		5040: Delta = 44'sb00000000000111111111111111111000000000000000;
		17519: Delta = 44'sb11111111110111111111111111111000000000000000;
		2670: Delta = 44'sb00000000010000000000000000001000000000000000;
		10009: Delta = 44'sb11111111110000000000000000001000000000000000;
		7610: Delta = 44'sb00000000001111111111111111111000000000000000;
		14949: Delta = 44'sb11111111101111111111111111111000000000000000;
		7810: Delta = 44'sb00000000100000000000000000001000000000000000;
		4869: Delta = 44'sb11111111100000000000000000001000000000000000;
		12750: Delta = 44'sb00000000011111111111111111111000000000000000;
		9809: Delta = 44'sb11111111011111111111111111111000000000000000;
		471: Delta = 44'sb00000001000000000000000000001000000000000000;
		12208: Delta = 44'sb11111111000000000000000000001000000000000000;
		5411: Delta = 44'sb00000000111111111111111111111000000000000000;
		17148: Delta = 44'sb11111110111111111111111111111000000000000000;
		3412: Delta = 44'sb00000010000000000000000000001000000000000000;
		9267: Delta = 44'sb11111110000000000000000000001000000000000000;
		8352: Delta = 44'sb00000001111111111111111111111000000000000000;
		14207: Delta = 44'sb11111101111111111111111111111000000000000000;
		9294: Delta = 44'sb00000100000000000000000000001000000000000000;
		3385: Delta = 44'sb11111100000000000000000000001000000000000000;
		14234: Delta = 44'sb00000011111111111111111111111000000000000000;
		8325: Delta = 44'sb11111011111111111111111111111000000000000000;
		3439: Delta = 44'sb00001000000000000000000000001000000000000000;
		9240: Delta = 44'sb11111000000000000000000000001000000000000000;
		8379: Delta = 44'sb00000111111111111111111111111000000000000000;
		14180: Delta = 44'sb11110111111111111111111111111000000000000000;
		9348: Delta = 44'sb00010000000000000000000000001000000000000000;
		3331: Delta = 44'sb11110000000000000000000000001000000000000000;
		14288: Delta = 44'sb00001111111111111111111111111000000000000000;
		8271: Delta = 44'sb11101111111111111111111111111000000000000000;
		3547: Delta = 44'sb00100000000000000000000000001000000000000000;
		9132: Delta = 44'sb11100000000000000000000000001000000000000000;
		8487: Delta = 44'sb00011111111111111111111111111000000000000000;
		14072: Delta = 44'sb11011111111111111111111111111000000000000000;
		9564: Delta = 44'sb01000000000000000000000000001000000000000000;
		3115: Delta = 44'sb11000000000000000000000000001000000000000000;
		14504: Delta = 44'sb00111111111111111111111111111000000000000000;
		8055: Delta = 44'sb10111111111111111111111111111000000000000000;
		2799: Delta = 44'sb00000000000000000000000000110000000000000000;
		14820: Delta = 44'sb11111111111111111111111111010000000000000000;
		10538: Delta = 44'sb00000000000000000000000001010000000000000000;
		7081: Delta = 44'sb11111111111111111111111110110000000000000000;
		8397: Delta = 44'sb00000000000000000000000010010000000000000000;
		16961: Delta = 44'sb11111111111111111111111110010000000000000000;
		658: Delta = 44'sb00000000000000000000000001110000000000000000;
		9222: Delta = 44'sb11111111111111111111111101110000000000000000;
		4115: Delta = 44'sb00000000000000000000000100010000000000000000;
		3624: Delta = 44'sb11111111111111111111111100010000000000000000;
		13995: Delta = 44'sb00000000000000000000000011110000000000000000;
		13504: Delta = 44'sb11111111111111111111111011110000000000000000;
		13170: Delta = 44'sb00000000000000000000001000010000000000000000;
		12188: Delta = 44'sb11111111111111111111111000010000000000000000;
		5431: Delta = 44'sb00000000000000000000000111110000000000000000;
		4449: Delta = 44'sb11111111111111111111110111110000000000000000;
		13661: Delta = 44'sb00000000000000000000010000010000000000000000;
		11697: Delta = 44'sb11111111111111111111110000010000000000000000;
		5922: Delta = 44'sb00000000000000000000001111110000000000000000;
		3958: Delta = 44'sb11111111111111111111101111110000000000000000;
		14643: Delta = 44'sb00000000000000000000100000010000000000000000;
		10715: Delta = 44'sb11111111111111111111100000010000000000000000;
		6904: Delta = 44'sb00000000000000000000011111110000000000000000;
		2976: Delta = 44'sb11111111111111111111011111110000000000000000;
		16607: Delta = 44'sb00000000000000000001000000010000000000000000;
		8751: Delta = 44'sb11111111111111111111000000010000000000000000;
		8868: Delta = 44'sb00000000000000000000111111110000000000000000;
		1012: Delta = 44'sb11111111111111111110111111110000000000000000;
		2916: Delta = 44'sb00000000000000000010000000010000000000000000;
		4823: Delta = 44'sb11111111111111111110000000010000000000000000;
		12796: Delta = 44'sb00000000000000000001111111110000000000000000;
		14703: Delta = 44'sb11111111111111111101111111110000000000000000;
		10772: Delta = 44'sb00000000000000000100000000010000000000000000;
		14586: Delta = 44'sb11111111111111111100000000010000000000000000;
		3033: Delta = 44'sb00000000000000000011111111110000000000000000;
		6847: Delta = 44'sb11111111111111111011111111110000000000000000;
		8865: Delta = 44'sb00000000000000001000000000010000000000000000;
		16493: Delta = 44'sb11111111111111111000000000010000000000000000;
		1126: Delta = 44'sb00000000000000000111111111110000000000000000;
		8754: Delta = 44'sb11111111111111110111111111110000000000000000;
		5051: Delta = 44'sb00000000000000010000000000010000000000000000;
		2688: Delta = 44'sb11111111111111110000000000010000000000000000;
		14931: Delta = 44'sb00000000000000001111111111110000000000000000;
		12568: Delta = 44'sb11111111111111101111111111110000000000000000;
		15042: Delta = 44'sb00000000000000100000000000010000000000000000;
		10316: Delta = 44'sb11111111111111100000000000010000000000000000;
		7303: Delta = 44'sb00000000000000011111111111110000000000000000;
		2577: Delta = 44'sb11111111111111011111111111110000000000000000;
		17405: Delta = 44'sb00000000000001000000000000010000000000000000;
		7953: Delta = 44'sb11111111111111000000000000010000000000000000;
		9666: Delta = 44'sb00000000000000111111111111110000000000000000;
		214: Delta = 44'sb11111111111110111111111111110000000000000000;
		4512: Delta = 44'sb00000000000010000000000000010000000000000000;
		3227: Delta = 44'sb11111111111110000000000000010000000000000000;
		14392: Delta = 44'sb00000000000001111111111111110000000000000000;
		13107: Delta = 44'sb11111111111101111111111111110000000000000000;
		13964: Delta = 44'sb00000000000100000000000000010000000000000000;
		11394: Delta = 44'sb11111111111100000000000000010000000000000000;
		6225: Delta = 44'sb00000000000011111111111111110000000000000000;
		3655: Delta = 44'sb11111111111011111111111111110000000000000000;
		15249: Delta = 44'sb00000000001000000000000000010000000000000000;
		10109: Delta = 44'sb11111111111000000000000000010000000000000000;
		7510: Delta = 44'sb00000000000111111111111111110000000000000000;
		2370: Delta = 44'sb11111111110111111111111111110000000000000000;
		200: Delta = 44'sb00000000010000000000000000010000000000000000;
		7539: Delta = 44'sb11111111110000000000000000010000000000000000;
		10080: Delta = 44'sb00000000001111111111111111110000000000000000;
		17419: Delta = 44'sb11111111101111111111111111110000000000000000;
		5340: Delta = 44'sb00000000100000000000000000010000000000000000;
		2399: Delta = 44'sb11111111100000000000000000010000000000000000;
		15220: Delta = 44'sb00000000011111111111111111110000000000000000;
		12279: Delta = 44'sb11111111011111111111111111110000000000000000;
		15620: Delta = 44'sb00000001000000000000000000010000000000000000;
		9738: Delta = 44'sb11111111000000000000000000010000000000000000;
		7881: Delta = 44'sb00000000111111111111111111110000000000000000;
		1999: Delta = 44'sb11111110111111111111111111110000000000000000;
		942: Delta = 44'sb00000010000000000000000000010000000000000000;
		6797: Delta = 44'sb11111110000000000000000000010000000000000000;
		10822: Delta = 44'sb00000001111111111111111111110000000000000000;
		16677: Delta = 44'sb11111101111111111111111111110000000000000000;
		6824: Delta = 44'sb00000100000000000000000000010000000000000000;
		915: Delta = 44'sb11111100000000000000000000010000000000000000;
		16704: Delta = 44'sb00000011111111111111111111110000000000000000;
		10795: Delta = 44'sb11111011111111111111111111110000000000000000;
		969: Delta = 44'sb00001000000000000000000000010000000000000000;
		6770: Delta = 44'sb11111000000000000000000000010000000000000000;
		10849: Delta = 44'sb00000111111111111111111111110000000000000000;
		16650: Delta = 44'sb11110111111111111111111111110000000000000000;
		6878: Delta = 44'sb00010000000000000000000000010000000000000000;
		861: Delta = 44'sb11110000000000000000000000010000000000000000;
		16758: Delta = 44'sb00001111111111111111111111110000000000000000;
		10741: Delta = 44'sb11101111111111111111111111110000000000000000;
		1077: Delta = 44'sb00100000000000000000000000010000000000000000;
		6662: Delta = 44'sb11100000000000000000000000010000000000000000;
		10957: Delta = 44'sb00011111111111111111111111110000000000000000;
		16542: Delta = 44'sb11011111111111111111111111110000000000000000;
		7094: Delta = 44'sb01000000000000000000000000010000000000000000;
		645: Delta = 44'sb11000000000000000000000000010000000000000000;
		16974: Delta = 44'sb00111111111111111111111111110000000000000000;
		10525: Delta = 44'sb10111111111111111111111111110000000000000000;
		5598: Delta = 44'sb00000000000000000000000001100000000000000000;
		12021: Delta = 44'sb11111111111111111111111110100000000000000000;
		3457: Delta = 44'sb00000000000000000000000010100000000000000000;
		14162: Delta = 44'sb11111111111111111111111101100000000000000000;
		16794: Delta = 44'sb00000000000000000000000100100000000000000000;
		16303: Delta = 44'sb11111111111111111111111100100000000000000000;
		1316: Delta = 44'sb00000000000000000000000011100000000000000000;
		825: Delta = 44'sb11111111111111111111111011100000000000000000;
		8230: Delta = 44'sb00000000000000000000001000100000000000000000;
		7248: Delta = 44'sb11111111111111111111111000100000000000000000;
		10371: Delta = 44'sb00000000000000000000000111100000000000000000;
		9389: Delta = 44'sb11111111111111111111110111100000000000000000;
		8721: Delta = 44'sb00000000000000000000010000100000000000000000;
		6757: Delta = 44'sb11111111111111111111110000100000000000000000;
		10862: Delta = 44'sb00000000000000000000001111100000000000000000;
		8898: Delta = 44'sb11111111111111111111101111100000000000000000;
		9703: Delta = 44'sb00000000000000000000100000100000000000000000;
		5775: Delta = 44'sb11111111111111111111100000100000000000000000;
		11844: Delta = 44'sb00000000000000000000011111100000000000000000;
		7916: Delta = 44'sb11111111111111111111011111100000000000000000;
		11667: Delta = 44'sb00000000000000000001000000100000000000000000;
		3811: Delta = 44'sb11111111111111111111000000100000000000000000;
		13808: Delta = 44'sb00000000000000000000111111100000000000000000;
		5952: Delta = 44'sb11111111111111111110111111100000000000000000;
		15595: Delta = 44'sb00000000000000000010000000100000000000000000;
		17502: Delta = 44'sb11111111111111111110000000100000000000000000;
		117: Delta = 44'sb00000000000000000001111111100000000000000000;
		2024: Delta = 44'sb11111111111111111101111111100000000000000000;
		5832: Delta = 44'sb00000000000000000100000000100000000000000000;
		9646: Delta = 44'sb11111111111111111100000000100000000000000000;
		7973: Delta = 44'sb00000000000000000011111111100000000000000000;
		11787: Delta = 44'sb11111111111111111011111111100000000000000000;
		3925: Delta = 44'sb00000000000000001000000000100000000000000000;
		11553: Delta = 44'sb11111111111111111000000000100000000000000000;
		6066: Delta = 44'sb00000000000000000111111111100000000000000000;
		13694: Delta = 44'sb11111111111111110111111111100000000000000000;
		111: Delta = 44'sb00000000000000010000000000100000000000000000;
		15367: Delta = 44'sb11111111111111110000000000100000000000000000;
		2252: Delta = 44'sb00000000000000001111111111100000000000000000;
		17508: Delta = 44'sb11111111111111101111111111100000000000000000;
		10102: Delta = 44'sb00000000000000100000000000100000000000000000;
		5376: Delta = 44'sb11111111111111100000000000100000000000000000;
		12243: Delta = 44'sb00000000000000011111111111100000000000000000;
		7517: Delta = 44'sb11111111111111011111111111100000000000000000;
		12465: Delta = 44'sb00000000000001000000000000100000000000000000;
		3013: Delta = 44'sb11111111111111000000000000100000000000000000;
		14606: Delta = 44'sb00000000000000111111111111100000000000000000;
		5154: Delta = 44'sb11111111111110111111111111100000000000000000;
		17191: Delta = 44'sb00000000000010000000000000100000000000000000;
		15906: Delta = 44'sb11111111111110000000000000100000000000000000;
		1713: Delta = 44'sb00000000000001111111111111100000000000000000;
		428: Delta = 44'sb11111111111101111111111111100000000000000000;
		9024: Delta = 44'sb00000000000100000000000000100000000000000000;
		6454: Delta = 44'sb11111111111100000000000000100000000000000000;
		11165: Delta = 44'sb00000000000011111111111111100000000000000000;
		8595: Delta = 44'sb11111111111011111111111111100000000000000000;
		10309: Delta = 44'sb00000000001000000000000000100000000000000000;
		5169: Delta = 44'sb11111111111000000000000000100000000000000000;
		12450: Delta = 44'sb00000000000111111111111111100000000000000000;
		7310: Delta = 44'sb11111111110111111111111111100000000000000000;
		12879: Delta = 44'sb00000000010000000000000000100000000000000000;
		2599: Delta = 44'sb11111111110000000000000000100000000000000000;
		15020: Delta = 44'sb00000000001111111111111111100000000000000000;
		4740: Delta = 44'sb11111111101111111111111111100000000000000000;
		400: Delta = 44'sb00000000100000000000000000100000000000000000;
		15078: Delta = 44'sb11111111100000000000000000100000000000000000;
		2541: Delta = 44'sb00000000011111111111111111100000000000000000;
		17219: Delta = 44'sb11111111011111111111111111100000000000000000;
		10680: Delta = 44'sb00000001000000000000000000100000000000000000;
		4798: Delta = 44'sb11111111000000000000000000100000000000000000;
		12821: Delta = 44'sb00000000111111111111111111100000000000000000;
		6939: Delta = 44'sb11111110111111111111111111100000000000000000;
		13621: Delta = 44'sb00000010000000000000000000100000000000000000;
		1857: Delta = 44'sb11111110000000000000000000100000000000000000;
		15762: Delta = 44'sb00000001111111111111111111100000000000000000;
		3998: Delta = 44'sb11111101111111111111111111100000000000000000;
		1884: Delta = 44'sb00000100000000000000000000100000000000000000;
		13594: Delta = 44'sb11111100000000000000000000100000000000000000;
		4025: Delta = 44'sb00000011111111111111111111100000000000000000;
		15735: Delta = 44'sb11111011111111111111111111100000000000000000;
		13648: Delta = 44'sb00001000000000000000000000100000000000000000;
		1830: Delta = 44'sb11111000000000000000000000100000000000000000;
		15789: Delta = 44'sb00000111111111111111111111100000000000000000;
		3971: Delta = 44'sb11110111111111111111111111100000000000000000;
		1938: Delta = 44'sb00010000000000000000000000100000000000000000;
		13540: Delta = 44'sb11110000000000000000000000100000000000000000;
		4079: Delta = 44'sb00001111111111111111111111100000000000000000;
		15681: Delta = 44'sb11101111111111111111111111100000000000000000;
		13756: Delta = 44'sb00100000000000000000000000100000000000000000;
		1722: Delta = 44'sb11100000000000000000000000100000000000000000;
		15897: Delta = 44'sb00011111111111111111111111100000000000000000;
		3863: Delta = 44'sb11011111111111111111111111100000000000000000;
		2154: Delta = 44'sb01000000000000000000000000100000000000000000;
		13324: Delta = 44'sb11000000000000000000000000100000000000000000;
		4295: Delta = 44'sb00111111111111111111111111100000000000000000;
		15465: Delta = 44'sb10111111111111111111111111100000000000000000;
		11196: Delta = 44'sb00000000000000000000000011000000000000000000;
		6423: Delta = 44'sb11111111111111111111111101000000000000000000;
		6914: Delta = 44'sb00000000000000000000000101000000000000000000;
		10705: Delta = 44'sb11111111111111111111111011000000000000000000;
		15969: Delta = 44'sb00000000000000000000001001000000000000000000;
		14987: Delta = 44'sb11111111111111111111111001000000000000000000;
		2632: Delta = 44'sb00000000000000000000000111000000000000000000;
		1650: Delta = 44'sb11111111111111111111110111000000000000000000;
		16460: Delta = 44'sb00000000000000000000010001000000000000000000;
		14496: Delta = 44'sb11111111111111111111110001000000000000000000;
		3123: Delta = 44'sb00000000000000000000001111000000000000000000;
		1159: Delta = 44'sb11111111111111111111101111000000000000000000;
		17442: Delta = 44'sb00000000000000000000100001000000000000000000;
		13514: Delta = 44'sb11111111111111111111100001000000000000000000;
		4105: Delta = 44'sb00000000000000000000011111000000000000000000;
		177: Delta = 44'sb11111111111111111111011111000000000000000000;
		1787: Delta = 44'sb00000000000000000001000001000000000000000000;
		11550: Delta = 44'sb11111111111111111111000001000000000000000000;
		6069: Delta = 44'sb00000000000000000000111111000000000000000000;
		15832: Delta = 44'sb11111111111111111110111111000000000000000000;
		5715: Delta = 44'sb00000000000000000010000001000000000000000000;
		7622: Delta = 44'sb11111111111111111110000001000000000000000000;
		9997: Delta = 44'sb00000000000000000001111111000000000000000000;
		11904: Delta = 44'sb11111111111111111101111111000000000000000000;
		13571: Delta = 44'sb00000000000000000100000001000000000000000000;
		17385: Delta = 44'sb11111111111111111100000001000000000000000000;
		234: Delta = 44'sb00000000000000000011111111000000000000000000;
		4048: Delta = 44'sb11111111111111111011111111000000000000000000;
		11664: Delta = 44'sb00000000000000001000000001000000000000000000;
		1673: Delta = 44'sb11111111111111111000000001000000000000000000;
		15946: Delta = 44'sb00000000000000000111111111000000000000000000;
		5955: Delta = 44'sb11111111111111110111111111000000000000000000;
		7850: Delta = 44'sb00000000000000010000000001000000000000000000;
		5487: Delta = 44'sb11111111111111110000000001000000000000000000;
		12132: Delta = 44'sb00000000000000001111111111000000000000000000;
		9769: Delta = 44'sb11111111111111101111111111000000000000000000;
		222: Delta = 44'sb00000000000000100000000001000000000000000000;
		13115: Delta = 44'sb11111111111111100000000001000000000000000000;
		4504: Delta = 44'sb00000000000000011111111111000000000000000000;
		17397: Delta = 44'sb11111111111111011111111111000000000000000000;
		2585: Delta = 44'sb00000000000001000000000001000000000000000000;
		10752: Delta = 44'sb11111111111111000000000001000000000000000000;
		6867: Delta = 44'sb00000000000000111111111111000000000000000000;
		15034: Delta = 44'sb11111111111110111111111111000000000000000000;
		7311: Delta = 44'sb00000000000010000000000001000000000000000000;
		6026: Delta = 44'sb11111111111110000000000001000000000000000000;
		11593: Delta = 44'sb00000000000001111111111111000000000000000000;
		10308: Delta = 44'sb11111111111101111111111111000000000000000000;
		16763: Delta = 44'sb00000000000100000000000001000000000000000000;
		14193: Delta = 44'sb11111111111100000000000001000000000000000000;
		3426: Delta = 44'sb00000000000011111111111111000000000000000000;
		856: Delta = 44'sb11111111111011111111111111000000000000000000;
		429: Delta = 44'sb00000000001000000000000001000000000000000000;
		12908: Delta = 44'sb11111111111000000000000001000000000000000000;
		4711: Delta = 44'sb00000000000111111111111111000000000000000000;
		17190: Delta = 44'sb11111111110111111111111111000000000000000000;
		2999: Delta = 44'sb00000000010000000000000001000000000000000000;
		10338: Delta = 44'sb11111111110000000000000001000000000000000000;
		7281: Delta = 44'sb00000000001111111111111111000000000000000000;
		14620: Delta = 44'sb11111111101111111111111111000000000000000000;
		8139: Delta = 44'sb00000000100000000000000001000000000000000000;
		5198: Delta = 44'sb11111111100000000000000001000000000000000000;
		12421: Delta = 44'sb00000000011111111111111111000000000000000000;
		9480: Delta = 44'sb11111111011111111111111111000000000000000000;
		800: Delta = 44'sb00000001000000000000000001000000000000000000;
		12537: Delta = 44'sb11111111000000000000000001000000000000000000;
		5082: Delta = 44'sb00000000111111111111111111000000000000000000;
		16819: Delta = 44'sb11111110111111111111111111000000000000000000;
		3741: Delta = 44'sb00000010000000000000000001000000000000000000;
		9596: Delta = 44'sb11111110000000000000000001000000000000000000;
		8023: Delta = 44'sb00000001111111111111111111000000000000000000;
		13878: Delta = 44'sb11111101111111111111111111000000000000000000;
		9623: Delta = 44'sb00000100000000000000000001000000000000000000;
		3714: Delta = 44'sb11111100000000000000000001000000000000000000;
		13905: Delta = 44'sb00000011111111111111111111000000000000000000;
		7996: Delta = 44'sb11111011111111111111111111000000000000000000;
		3768: Delta = 44'sb00001000000000000000000001000000000000000000;
		9569: Delta = 44'sb11111000000000000000000001000000000000000000;
		8050: Delta = 44'sb00000111111111111111111111000000000000000000;
		13851: Delta = 44'sb11110111111111111111111111000000000000000000;
		9677: Delta = 44'sb00010000000000000000000001000000000000000000;
		3660: Delta = 44'sb11110000000000000000000001000000000000000000;
		13959: Delta = 44'sb00001111111111111111111111000000000000000000;
		7942: Delta = 44'sb11101111111111111111111111000000000000000000;
		3876: Delta = 44'sb00100000000000000000000001000000000000000000;
		9461: Delta = 44'sb11100000000000000000000001000000000000000000;
		8158: Delta = 44'sb00011111111111111111111111000000000000000000;
		13743: Delta = 44'sb11011111111111111111111111000000000000000000;
		9893: Delta = 44'sb01000000000000000000000001000000000000000000;
		3444: Delta = 44'sb11000000000000000000000001000000000000000000;
		14175: Delta = 44'sb00111111111111111111111111000000000000000000;
		7726: Delta = 44'sb10111111111111111111111111000000000000000000;
		4773: Delta = 44'sb00000000000000000000000110000000000000000000;
		12846: Delta = 44'sb11111111111111111111111010000000000000000000;
		13828: Delta = 44'sb00000000000000000000001010000000000000000000;
		3791: Delta = 44'sb11111111111111111111110110000000000000000000;
		14319: Delta = 44'sb00000000000000000000010010000000000000000000;
		12355: Delta = 44'sb11111111111111111111110010000000000000000000;
		5264: Delta = 44'sb00000000000000000000001110000000000000000000;
		3300: Delta = 44'sb11111111111111111111101110000000000000000000;
		15301: Delta = 44'sb00000000000000000000100010000000000000000000;
		11373: Delta = 44'sb11111111111111111111100010000000000000000000;
		6246: Delta = 44'sb00000000000000000000011110000000000000000000;
		2318: Delta = 44'sb11111111111111111111011110000000000000000000;
		17265: Delta = 44'sb00000000000000000001000010000000000000000000;
		9409: Delta = 44'sb11111111111111111111000010000000000000000000;
		8210: Delta = 44'sb00000000000000000000111110000000000000000000;
		354: Delta = 44'sb11111111111111111110111110000000000000000000;
		3574: Delta = 44'sb00000000000000000010000010000000000000000000;
		5481: Delta = 44'sb11111111111111111110000010000000000000000000;
		12138: Delta = 44'sb00000000000000000001111110000000000000000000;
		14045: Delta = 44'sb11111111111111111101111110000000000000000000;
		11430: Delta = 44'sb00000000000000000100000010000000000000000000;
		15244: Delta = 44'sb11111111111111111100000010000000000000000000;
		2375: Delta = 44'sb00000000000000000011111110000000000000000000;
		6189: Delta = 44'sb11111111111111111011111110000000000000000000;
		9523: Delta = 44'sb00000000000000001000000010000000000000000000;
		17151: Delta = 44'sb11111111111111111000000010000000000000000000;
		468: Delta = 44'sb00000000000000000111111110000000000000000000;
		8096: Delta = 44'sb11111111111111110111111110000000000000000000;
		5709: Delta = 44'sb00000000000000010000000010000000000000000000;
		3346: Delta = 44'sb11111111111111110000000010000000000000000000;
		14273: Delta = 44'sb00000000000000001111111110000000000000000000;
		11910: Delta = 44'sb11111111111111101111111110000000000000000000;
		15700: Delta = 44'sb00000000000000100000000010000000000000000000;
		10974: Delta = 44'sb11111111111111100000000010000000000000000000;
		6645: Delta = 44'sb00000000000000011111111110000000000000000000;
		1919: Delta = 44'sb11111111111111011111111110000000000000000000;
		444: Delta = 44'sb00000000000001000000000010000000000000000000;
		8611: Delta = 44'sb11111111111111000000000010000000000000000000;
		9008: Delta = 44'sb00000000000000111111111110000000000000000000;
		17175: Delta = 44'sb11111111111110111111111110000000000000000000;
		5170: Delta = 44'sb00000000000010000000000010000000000000000000;
		3885: Delta = 44'sb11111111111110000000000010000000000000000000;
		13734: Delta = 44'sb00000000000001111111111110000000000000000000;
		12449: Delta = 44'sb11111111111101111111111110000000000000000000;
		14622: Delta = 44'sb00000000000100000000000010000000000000000000;
		12052: Delta = 44'sb11111111111100000000000010000000000000000000;
		5567: Delta = 44'sb00000000000011111111111110000000000000000000;
		2997: Delta = 44'sb11111111111011111111111110000000000000000000;
		15907: Delta = 44'sb00000000001000000000000010000000000000000000;
		10767: Delta = 44'sb11111111111000000000000010000000000000000000;
		6852: Delta = 44'sb00000000000111111111111110000000000000000000;
		1712: Delta = 44'sb11111111110111111111111110000000000000000000;
		858: Delta = 44'sb00000000010000000000000010000000000000000000;
		8197: Delta = 44'sb11111111110000000000000010000000000000000000;
		9422: Delta = 44'sb00000000001111111111111110000000000000000000;
		16761: Delta = 44'sb11111111101111111111111110000000000000000000;
		5998: Delta = 44'sb00000000100000000000000010000000000000000000;
		3057: Delta = 44'sb11111111100000000000000010000000000000000000;
		14562: Delta = 44'sb00000000011111111111111110000000000000000000;
		11621: Delta = 44'sb11111111011111111111111110000000000000000000;
		16278: Delta = 44'sb00000001000000000000000010000000000000000000;
		10396: Delta = 44'sb11111111000000000000000010000000000000000000;
		7223: Delta = 44'sb00000000111111111111111110000000000000000000;
		1341: Delta = 44'sb11111110111111111111111110000000000000000000;
		1600: Delta = 44'sb00000010000000000000000010000000000000000000;
		7455: Delta = 44'sb11111110000000000000000010000000000000000000;
		10164: Delta = 44'sb00000001111111111111111110000000000000000000;
		16019: Delta = 44'sb11111101111111111111111110000000000000000000;
		7482: Delta = 44'sb00000100000000000000000010000000000000000000;
		1573: Delta = 44'sb11111100000000000000000010000000000000000000;
		16046: Delta = 44'sb00000011111111111111111110000000000000000000;
		10137: Delta = 44'sb11111011111111111111111110000000000000000000;
		1627: Delta = 44'sb00001000000000000000000010000000000000000000;
		7428: Delta = 44'sb11111000000000000000000010000000000000000000;
		10191: Delta = 44'sb00000111111111111111111110000000000000000000;
		15992: Delta = 44'sb11110111111111111111111110000000000000000000;
		7536: Delta = 44'sb00010000000000000000000010000000000000000000;
		1519: Delta = 44'sb11110000000000000000000010000000000000000000;
		16100: Delta = 44'sb00001111111111111111111110000000000000000000;
		10083: Delta = 44'sb11101111111111111111111110000000000000000000;
		1735: Delta = 44'sb00100000000000000000000010000000000000000000;
		7320: Delta = 44'sb11100000000000000000000010000000000000000000;
		10299: Delta = 44'sb00011111111111111111111110000000000000000000;
		15884: Delta = 44'sb11011111111111111111111110000000000000000000;
		7752: Delta = 44'sb01000000000000000000000010000000000000000000;
		1303: Delta = 44'sb11000000000000000000000010000000000000000000;
		16316: Delta = 44'sb00111111111111111111111110000000000000000000;
		9867: Delta = 44'sb10111111111111111111111110000000000000000000;
		9546: Delta = 44'sb00000000000000000000001100000000000000000000;
		8073: Delta = 44'sb11111111111111111111110100000000000000000000;
		10037: Delta = 44'sb00000000000000000000010100000000000000000000;
		7582: Delta = 44'sb11111111111111111111101100000000000000000000;
		11019: Delta = 44'sb00000000000000000000100100000000000000000000;
		7091: Delta = 44'sb11111111111111111111100100000000000000000000;
		10528: Delta = 44'sb00000000000000000000011100000000000000000000;
		6600: Delta = 44'sb11111111111111111111011100000000000000000000;
		12983: Delta = 44'sb00000000000000000001000100000000000000000000;
		5127: Delta = 44'sb11111111111111111111000100000000000000000000;
		12492: Delta = 44'sb00000000000000000000111100000000000000000000;
		4636: Delta = 44'sb11111111111111111110111100000000000000000000;
		16911: Delta = 44'sb00000000000000000010000100000000000000000000;
		1199: Delta = 44'sb11111111111111111110000100000000000000000000;
		16420: Delta = 44'sb00000000000000000001111100000000000000000000;
		708: Delta = 44'sb11111111111111111101111100000000000000000000;
		7148: Delta = 44'sb00000000000000000100000100000000000000000000;
		10962: Delta = 44'sb11111111111111111100000100000000000000000000;
		6657: Delta = 44'sb00000000000000000011111100000000000000000000;
		10471: Delta = 44'sb11111111111111111011111100000000000000000000;
		5241: Delta = 44'sb00000000000000001000000100000000000000000000;
		12869: Delta = 44'sb11111111111111111000000100000000000000000000;
		4750: Delta = 44'sb00000000000000000111111100000000000000000000;
		12378: Delta = 44'sb11111111111111110111111100000000000000000000;
		1427: Delta = 44'sb00000000000000010000000100000000000000000000;
		16683: Delta = 44'sb11111111111111110000000100000000000000000000;
		936: Delta = 44'sb00000000000000001111111100000000000000000000;
		16192: Delta = 44'sb11111111111111101111111100000000000000000000;
		11418: Delta = 44'sb00000000000000100000000100000000000000000000;
		6692: Delta = 44'sb11111111111111100000000100000000000000000000;
		10927: Delta = 44'sb00000000000000011111111100000000000000000000;
		6201: Delta = 44'sb11111111111111011111111100000000000000000000;
		13781: Delta = 44'sb00000000000001000000000100000000000000000000;
		4329: Delta = 44'sb11111111111111000000000100000000000000000000;
		13290: Delta = 44'sb00000000000000111111111100000000000000000000;
		3838: Delta = 44'sb11111111111110111111111100000000000000000000;
		888: Delta = 44'sb00000000000010000000000100000000000000000000;
		17222: Delta = 44'sb11111111111110000000000100000000000000000000;
		397: Delta = 44'sb00000000000001111111111100000000000000000000;
		16731: Delta = 44'sb11111111111101111111111100000000000000000000;
		10340: Delta = 44'sb00000000000100000000000100000000000000000000;
		7770: Delta = 44'sb11111111111100000000000100000000000000000000;
		9849: Delta = 44'sb00000000000011111111111100000000000000000000;
		7279: Delta = 44'sb11111111111011111111111100000000000000000000;
		11625: Delta = 44'sb00000000001000000000000100000000000000000000;
		6485: Delta = 44'sb11111111111000000000000100000000000000000000;
		11134: Delta = 44'sb00000000000111111111111100000000000000000000;
		5994: Delta = 44'sb11111111110111111111111100000000000000000000;
		14195: Delta = 44'sb00000000010000000000000100000000000000000000;
		3915: Delta = 44'sb11111111110000000000000100000000000000000000;
		13704: Delta = 44'sb00000000001111111111111100000000000000000000;
		3424: Delta = 44'sb11111111101111111111111100000000000000000000;
		1716: Delta = 44'sb00000000100000000000000100000000000000000000;
		16394: Delta = 44'sb11111111100000000000000100000000000000000000;
		1225: Delta = 44'sb00000000011111111111111100000000000000000000;
		15903: Delta = 44'sb11111111011111111111111100000000000000000000;
		11996: Delta = 44'sb00000001000000000000000100000000000000000000;
		6114: Delta = 44'sb11111111000000000000000100000000000000000000;
		11505: Delta = 44'sb00000000111111111111111100000000000000000000;
		5623: Delta = 44'sb11111110111111111111111100000000000000000000;
		14937: Delta = 44'sb00000010000000000000000100000000000000000000;
		3173: Delta = 44'sb11111110000000000000000100000000000000000000;
		14446: Delta = 44'sb00000001111111111111111100000000000000000000;
		2682: Delta = 44'sb11111101111111111111111100000000000000000000;
		3200: Delta = 44'sb00000100000000000000000100000000000000000000;
		14910: Delta = 44'sb11111100000000000000000100000000000000000000;
		2709: Delta = 44'sb00000011111111111111111100000000000000000000;
		14419: Delta = 44'sb11111011111111111111111100000000000000000000;
		14964: Delta = 44'sb00001000000000000000000100000000000000000000;
		3146: Delta = 44'sb11111000000000000000000100000000000000000000;
		14473: Delta = 44'sb00000111111111111111111100000000000000000000;
		2655: Delta = 44'sb11110111111111111111111100000000000000000000;
		3254: Delta = 44'sb00010000000000000000000100000000000000000000;
		14856: Delta = 44'sb11110000000000000000000100000000000000000000;
		2763: Delta = 44'sb00001111111111111111111100000000000000000000;
		14365: Delta = 44'sb11101111111111111111111100000000000000000000;
		15072: Delta = 44'sb00100000000000000000000100000000000000000000;
		3038: Delta = 44'sb11100000000000000000000100000000000000000000;
		14581: Delta = 44'sb00011111111111111111111100000000000000000000;
		2547: Delta = 44'sb11011111111111111111111100000000000000000000;
		3470: Delta = 44'sb01000000000000000000000100000000000000000000;
		14640: Delta = 44'sb11000000000000000000000100000000000000000000;
		2979: Delta = 44'sb00111111111111111111111100000000000000000000;
		14149: Delta = 44'sb10111111111111111111111100000000000000000000;
		1473: Delta = 44'sb00000000000000000000011000000000000000000000;
		16146: Delta = 44'sb11111111111111111111101000000000000000000000;
		2455: Delta = 44'sb00000000000000000000101000000000000000000000;
		15164: Delta = 44'sb11111111111111111111011000000000000000000000;
		4419: Delta = 44'sb00000000000000000001001000000000000000000000;
		14182: Delta = 44'sb11111111111111111111001000000000000000000000;
		3437: Delta = 44'sb00000000000000000000111000000000000000000000;
		13200: Delta = 44'sb11111111111111111110111000000000000000000000;
		8347: Delta = 44'sb00000000000000000010001000000000000000000000;
		10254: Delta = 44'sb11111111111111111110001000000000000000000000;
		7365: Delta = 44'sb00000000000000000001111000000000000000000000;
		9272: Delta = 44'sb11111111111111111101111000000000000000000000;
		16203: Delta = 44'sb00000000000000000100001000000000000000000000;
		2398: Delta = 44'sb11111111111111111100001000000000000000000000;
		15221: Delta = 44'sb00000000000000000011111000000000000000000000;
		1416: Delta = 44'sb11111111111111111011111000000000000000000000;
		14296: Delta = 44'sb00000000000000001000001000000000000000000000;
		4305: Delta = 44'sb11111111111111111000001000000000000000000000;
		13314: Delta = 44'sb00000000000000000111111000000000000000000000;
		3323: Delta = 44'sb11111111111111110111111000000000000000000000;
		10482: Delta = 44'sb00000000000000010000001000000000000000000000;
		8119: Delta = 44'sb11111111111111110000001000000000000000000000;
		9500: Delta = 44'sb00000000000000001111111000000000000000000000;
		7137: Delta = 44'sb11111111111111101111111000000000000000000000;
		2854: Delta = 44'sb00000000000000100000001000000000000000000000;
		15747: Delta = 44'sb11111111111111100000001000000000000000000000;
		1872: Delta = 44'sb00000000000000011111111000000000000000000000;
		14765: Delta = 44'sb11111111111111011111111000000000000000000000;
		5217: Delta = 44'sb00000000000001000000001000000000000000000000;
		13384: Delta = 44'sb11111111111111000000001000000000000000000000;
		4235: Delta = 44'sb00000000000000111111111000000000000000000000;
		12402: Delta = 44'sb11111111111110111111111000000000000000000000;
		9943: Delta = 44'sb00000000000010000000001000000000000000000000;
		8658: Delta = 44'sb11111111111110000000001000000000000000000000;
		8961: Delta = 44'sb00000000000001111111111000000000000000000000;
		7676: Delta = 44'sb11111111111101111111111000000000000000000000;
		1776: Delta = 44'sb00000000000100000000001000000000000000000000;
		16825: Delta = 44'sb11111111111100000000001000000000000000000000;
		794: Delta = 44'sb00000000000011111111111000000000000000000000;
		15843: Delta = 44'sb11111111111011111111111000000000000000000000;
		3061: Delta = 44'sb00000000001000000000001000000000000000000000;
		15540: Delta = 44'sb11111111111000000000001000000000000000000000;
		2079: Delta = 44'sb00000000000111111111111000000000000000000000;
		14558: Delta = 44'sb11111111110111111111111000000000000000000000;
		5631: Delta = 44'sb00000000010000000000001000000000000000000000;
		12970: Delta = 44'sb11111111110000000000001000000000000000000000;
		4649: Delta = 44'sb00000000001111111111111000000000000000000000;
		11988: Delta = 44'sb11111111101111111111111000000000000000000000;
		10771: Delta = 44'sb00000000100000000000001000000000000000000000;
		7830: Delta = 44'sb11111111100000000000001000000000000000000000;
		9789: Delta = 44'sb00000000011111111111111000000000000000000000;
		6848: Delta = 44'sb11111111011111111111111000000000000000000000;
		3432: Delta = 44'sb00000001000000000000001000000000000000000000;
		15169: Delta = 44'sb11111111000000000000001000000000000000000000;
		2450: Delta = 44'sb00000000111111111111111000000000000000000000;
		14187: Delta = 44'sb11111110111111111111111000000000000000000000;
		6373: Delta = 44'sb00000010000000000000001000000000000000000000;
		12228: Delta = 44'sb11111110000000000000001000000000000000000000;
		5391: Delta = 44'sb00000001111111111111111000000000000000000000;
		11246: Delta = 44'sb11111101111111111111111000000000000000000000;
		12255: Delta = 44'sb00000100000000000000001000000000000000000000;
		6346: Delta = 44'sb11111100000000000000001000000000000000000000;
		11273: Delta = 44'sb00000011111111111111111000000000000000000000;
		5364: Delta = 44'sb11111011111111111111111000000000000000000000;
		6400: Delta = 44'sb00001000000000000000001000000000000000000000;
		12201: Delta = 44'sb11111000000000000000001000000000000000000000;
		5418: Delta = 44'sb00000111111111111111111000000000000000000000;
		11219: Delta = 44'sb11110111111111111111111000000000000000000000;
		12309: Delta = 44'sb00010000000000000000001000000000000000000000;
		6292: Delta = 44'sb11110000000000000000001000000000000000000000;
		11327: Delta = 44'sb00001111111111111111111000000000000000000000;
		5310: Delta = 44'sb11101111111111111111111000000000000000000000;
		6508: Delta = 44'sb00100000000000000000001000000000000000000000;
		12093: Delta = 44'sb11100000000000000000001000000000000000000000;
		5526: Delta = 44'sb00011111111111111111111000000000000000000000;
		11111: Delta = 44'sb11011111111111111111111000000000000000000000;
		12525: Delta = 44'sb01000000000000000000001000000000000000000000;
		6076: Delta = 44'sb11000000000000000000001000000000000000000000;
		11543: Delta = 44'sb00111111111111111111111000000000000000000000;
		5094: Delta = 44'sb10111111111111111111111000000000000000000000;
		2946: Delta = 44'sb00000000000000000000110000000000000000000000;
		14673: Delta = 44'sb11111111111111111111010000000000000000000000;
		4910: Delta = 44'sb00000000000000000001010000000000000000000000;
		12709: Delta = 44'sb11111111111111111110110000000000000000000000;
		8838: Delta = 44'sb00000000000000000010010000000000000000000000;
		10745: Delta = 44'sb11111111111111111110010000000000000000000000;
		6874: Delta = 44'sb00000000000000000001110000000000000000000000;
		8781: Delta = 44'sb11111111111111111101110000000000000000000000;
		16694: Delta = 44'sb00000000000000000100010000000000000000000000;
		2889: Delta = 44'sb11111111111111111100010000000000000000000000;
		14730: Delta = 44'sb00000000000000000011110000000000000000000000;
		925: Delta = 44'sb11111111111111111011110000000000000000000000;
		14787: Delta = 44'sb00000000000000001000010000000000000000000000;
		4796: Delta = 44'sb11111111111111111000010000000000000000000000;
		12823: Delta = 44'sb00000000000000000111110000000000000000000000;
		2832: Delta = 44'sb11111111111111110111110000000000000000000000;
		10973: Delta = 44'sb00000000000000010000010000000000000000000000;
		8610: Delta = 44'sb11111111111111110000010000000000000000000000;
		9009: Delta = 44'sb00000000000000001111110000000000000000000000;
		6646: Delta = 44'sb11111111111111101111110000000000000000000000;
		3345: Delta = 44'sb00000000000000100000010000000000000000000000;
		16238: Delta = 44'sb11111111111111100000010000000000000000000000;
		1381: Delta = 44'sb00000000000000011111110000000000000000000000;
		14274: Delta = 44'sb11111111111111011111110000000000000000000000;
		5708: Delta = 44'sb00000000000001000000010000000000000000000000;
		13875: Delta = 44'sb11111111111111000000010000000000000000000000;
		3744: Delta = 44'sb00000000000000111111110000000000000000000000;
		11911: Delta = 44'sb11111111111110111111110000000000000000000000;
		10434: Delta = 44'sb00000000000010000000010000000000000000000000;
		9149: Delta = 44'sb11111111111110000000010000000000000000000000;
		8470: Delta = 44'sb00000000000001111111110000000000000000000000;
		7185: Delta = 44'sb11111111111101111111110000000000000000000000;
		2267: Delta = 44'sb00000000000100000000010000000000000000000000;
		17316: Delta = 44'sb11111111111100000000010000000000000000000000;
		303: Delta = 44'sb00000000000011111111110000000000000000000000;
		15352: Delta = 44'sb11111111111011111111110000000000000000000000;
		3552: Delta = 44'sb00000000001000000000010000000000000000000000;
		16031: Delta = 44'sb11111111111000000000010000000000000000000000;
		1588: Delta = 44'sb00000000000111111111110000000000000000000000;
		14067: Delta = 44'sb11111111110111111111110000000000000000000000;
		6122: Delta = 44'sb00000000010000000000010000000000000000000000;
		13461: Delta = 44'sb11111111110000000000010000000000000000000000;
		4158: Delta = 44'sb00000000001111111111110000000000000000000000;
		11497: Delta = 44'sb11111111101111111111110000000000000000000000;
		11262: Delta = 44'sb00000000100000000000010000000000000000000000;
		8321: Delta = 44'sb11111111100000000000010000000000000000000000;
		9298: Delta = 44'sb00000000011111111111110000000000000000000000;
		6357: Delta = 44'sb11111111011111111111110000000000000000000000;
		3923: Delta = 44'sb00000001000000000000010000000000000000000000;
		15660: Delta = 44'sb11111111000000000000010000000000000000000000;
		1959: Delta = 44'sb00000000111111111111110000000000000000000000;
		13696: Delta = 44'sb11111110111111111111110000000000000000000000;
		6864: Delta = 44'sb00000010000000000000010000000000000000000000;
		12719: Delta = 44'sb11111110000000000000010000000000000000000000;
		4900: Delta = 44'sb00000001111111111111110000000000000000000000;
		10755: Delta = 44'sb11111101111111111111110000000000000000000000;
		12746: Delta = 44'sb00000100000000000000010000000000000000000000;
		6837: Delta = 44'sb11111100000000000000010000000000000000000000;
		10782: Delta = 44'sb00000011111111111111110000000000000000000000;
		4873: Delta = 44'sb11111011111111111111110000000000000000000000;
		6891: Delta = 44'sb00001000000000000000010000000000000000000000;
		12692: Delta = 44'sb11111000000000000000010000000000000000000000;
		4927: Delta = 44'sb00000111111111111111110000000000000000000000;
		10728: Delta = 44'sb11110111111111111111110000000000000000000000;
		12800: Delta = 44'sb00010000000000000000010000000000000000000000;
		6783: Delta = 44'sb11110000000000000000010000000000000000000000;
		10836: Delta = 44'sb00001111111111111111110000000000000000000000;
		4819: Delta = 44'sb11101111111111111111110000000000000000000000;
		6999: Delta = 44'sb00100000000000000000010000000000000000000000;
		12584: Delta = 44'sb11100000000000000000010000000000000000000000;
		5035: Delta = 44'sb00011111111111111111110000000000000000000000;
		10620: Delta = 44'sb11011111111111111111110000000000000000000000;
		13016: Delta = 44'sb01000000000000000000010000000000000000000000;
		6567: Delta = 44'sb11000000000000000000010000000000000000000000;
		11052: Delta = 44'sb00111111111111111111110000000000000000000000;
		4603: Delta = 44'sb10111111111111111111110000000000000000000000;
		5892: Delta = 44'sb00000000000000000001100000000000000000000000;
		11727: Delta = 44'sb11111111111111111110100000000000000000000000;
		9820: Delta = 44'sb00000000000000000010100000000000000000000000;
		7799: Delta = 44'sb11111111111111111101100000000000000000000000;
		57: Delta = 44'sb00000000000000000100100000000000000000000000;
		3871: Delta = 44'sb11111111111111111100100000000000000000000000;
		13748: Delta = 44'sb00000000000000000011100000000000000000000000;
		17562: Delta = 44'sb11111111111111111011100000000000000000000000;
		15769: Delta = 44'sb00000000000000001000100000000000000000000000;
		5778: Delta = 44'sb11111111111111111000100000000000000000000000;
		11841: Delta = 44'sb00000000000000000111100000000000000000000000;
		1850: Delta = 44'sb11111111111111110111100000000000000000000000;
		11955: Delta = 44'sb00000000000000010000100000000000000000000000;
		9592: Delta = 44'sb11111111111111110000100000000000000000000000;
		8027: Delta = 44'sb00000000000000001111100000000000000000000000;
		5664: Delta = 44'sb11111111111111101111100000000000000000000000;
		4327: Delta = 44'sb00000000000000100000100000000000000000000000;
		17220: Delta = 44'sb11111111111111100000100000000000000000000000;
		399: Delta = 44'sb00000000000000011111100000000000000000000000;
		13292: Delta = 44'sb11111111111111011111100000000000000000000000;
		6690: Delta = 44'sb00000000000001000000100000000000000000000000;
		14857: Delta = 44'sb11111111111111000000100000000000000000000000;
		2762: Delta = 44'sb00000000000000111111100000000000000000000000;
		10929: Delta = 44'sb11111111111110111111100000000000000000000000;
		11416: Delta = 44'sb00000000000010000000100000000000000000000000;
		10131: Delta = 44'sb11111111111110000000100000000000000000000000;
		7488: Delta = 44'sb00000000000001111111100000000000000000000000;
		6203: Delta = 44'sb11111111111101111111100000000000000000000000;
		3249: Delta = 44'sb00000000000100000000100000000000000000000000;
		679: Delta = 44'sb11111111111100000000100000000000000000000000;
		16940: Delta = 44'sb00000000000011111111100000000000000000000000;
		14370: Delta = 44'sb11111111111011111111100000000000000000000000;
		4534: Delta = 44'sb00000000001000000000100000000000000000000000;
		17013: Delta = 44'sb11111111111000000000100000000000000000000000;
		606: Delta = 44'sb00000000000111111111100000000000000000000000;
		13085: Delta = 44'sb11111111110111111111100000000000000000000000;
		7104: Delta = 44'sb00000000010000000000100000000000000000000000;
		14443: Delta = 44'sb11111111110000000000100000000000000000000000;
		3176: Delta = 44'sb00000000001111111111100000000000000000000000;
		10515: Delta = 44'sb11111111101111111111100000000000000000000000;
		12244: Delta = 44'sb00000000100000000000100000000000000000000000;
		9303: Delta = 44'sb11111111100000000000100000000000000000000000;
		8316: Delta = 44'sb00000000011111111111100000000000000000000000;
		5375: Delta = 44'sb11111111011111111111100000000000000000000000;
		4905: Delta = 44'sb00000001000000000000100000000000000000000000;
		16642: Delta = 44'sb11111111000000000000100000000000000000000000;
		977: Delta = 44'sb00000000111111111111100000000000000000000000;
		12714: Delta = 44'sb11111110111111111111100000000000000000000000;
		7846: Delta = 44'sb00000010000000000000100000000000000000000000;
		13701: Delta = 44'sb11111110000000000000100000000000000000000000;
		3918: Delta = 44'sb00000001111111111111100000000000000000000000;
		9773: Delta = 44'sb11111101111111111111100000000000000000000000;
		13728: Delta = 44'sb00000100000000000000100000000000000000000000;
		7819: Delta = 44'sb11111100000000000000100000000000000000000000;
		9800: Delta = 44'sb00000011111111111111100000000000000000000000;
		3891: Delta = 44'sb11111011111111111111100000000000000000000000;
		7873: Delta = 44'sb00001000000000000000100000000000000000000000;
		13674: Delta = 44'sb11111000000000000000100000000000000000000000;
		3945: Delta = 44'sb00000111111111111111100000000000000000000000;
		9746: Delta = 44'sb11110111111111111111100000000000000000000000;
		13782: Delta = 44'sb00010000000000000000100000000000000000000000;
		7765: Delta = 44'sb11110000000000000000100000000000000000000000;
		9854: Delta = 44'sb00001111111111111111100000000000000000000000;
		3837: Delta = 44'sb11101111111111111111100000000000000000000000;
		7981: Delta = 44'sb00100000000000000000100000000000000000000000;
		13566: Delta = 44'sb11100000000000000000100000000000000000000000;
		4053: Delta = 44'sb00011111111111111111100000000000000000000000;
		9638: Delta = 44'sb11011111111111111111100000000000000000000000;
		13998: Delta = 44'sb01000000000000000000100000000000000000000000;
		7549: Delta = 44'sb11000000000000000000100000000000000000000000;
		10070: Delta = 44'sb00111111111111111111100000000000000000000000;
		3621: Delta = 44'sb10111111111111111111100000000000000000000000;
		11784: Delta = 44'sb00000000000000000011000000000000000000000000;
		5835: Delta = 44'sb11111111111111111101000000000000000000000000;
		2021: Delta = 44'sb00000000000000000101000000000000000000000000;
		15598: Delta = 44'sb11111111111111111011000000000000000000000000;
		114: Delta = 44'sb00000000000000001001000000000000000000000000;
		7742: Delta = 44'sb11111111111111111001000000000000000000000000;
		9877: Delta = 44'sb00000000000000000111000000000000000000000000;
		17505: Delta = 44'sb11111111111111110111000000000000000000000000;
		13919: Delta = 44'sb00000000000000010001000000000000000000000000;
		11556: Delta = 44'sb11111111111111110001000000000000000000000000;
		6063: Delta = 44'sb00000000000000001111000000000000000000000000;
		3700: Delta = 44'sb11111111111111101111000000000000000000000000;
		6291: Delta = 44'sb00000000000000100001000000000000000000000000;
		1565: Delta = 44'sb11111111111111100001000000000000000000000000;
		16054: Delta = 44'sb00000000000000011111000000000000000000000000;
		11328: Delta = 44'sb11111111111111011111000000000000000000000000;
		8654: Delta = 44'sb00000000000001000001000000000000000000000000;
		16821: Delta = 44'sb11111111111111000001000000000000000000000000;
		798: Delta = 44'sb00000000000000111111000000000000000000000000;
		8965: Delta = 44'sb11111111111110111111000000000000000000000000;
		13380: Delta = 44'sb00000000000010000001000000000000000000000000;
		12095: Delta = 44'sb11111111111110000001000000000000000000000000;
		5524: Delta = 44'sb00000000000001111111000000000000000000000000;
		4239: Delta = 44'sb11111111111101111111000000000000000000000000;
		5213: Delta = 44'sb00000000000100000001000000000000000000000000;
		2643: Delta = 44'sb11111111111100000001000000000000000000000000;
		14976: Delta = 44'sb00000000000011111111000000000000000000000000;
		12406: Delta = 44'sb11111111111011111111000000000000000000000000;
		6498: Delta = 44'sb00000000001000000001000000000000000000000000;
		1358: Delta = 44'sb11111111111000000001000000000000000000000000;
		16261: Delta = 44'sb00000000000111111111000000000000000000000000;
		11121: Delta = 44'sb11111111110111111111000000000000000000000000;
		9068: Delta = 44'sb00000000010000000001000000000000000000000000;
		16407: Delta = 44'sb11111111110000000001000000000000000000000000;
		1212: Delta = 44'sb00000000001111111111000000000000000000000000;
		8551: Delta = 44'sb11111111101111111111000000000000000000000000;
		14208: Delta = 44'sb00000000100000000001000000000000000000000000;
		11267: Delta = 44'sb11111111100000000001000000000000000000000000;
		6352: Delta = 44'sb00000000011111111111000000000000000000000000;
		3411: Delta = 44'sb11111111011111111111000000000000000000000000;
		6869: Delta = 44'sb00000001000000000001000000000000000000000000;
		987: Delta = 44'sb11111111000000000001000000000000000000000000;
		16632: Delta = 44'sb00000000111111111111000000000000000000000000;
		10750: Delta = 44'sb11111110111111111111000000000000000000000000;
		9810: Delta = 44'sb00000010000000000001000000000000000000000000;
		15665: Delta = 44'sb11111110000000000001000000000000000000000000;
		1954: Delta = 44'sb00000001111111111111000000000000000000000000;
		7809: Delta = 44'sb11111101111111111111000000000000000000000000;
		15692: Delta = 44'sb00000100000000000001000000000000000000000000;
		9783: Delta = 44'sb11111100000000000001000000000000000000000000;
		7836: Delta = 44'sb00000011111111111111000000000000000000000000;
		1927: Delta = 44'sb11111011111111111111000000000000000000000000;
		9837: Delta = 44'sb00001000000000000001000000000000000000000000;
		15638: Delta = 44'sb11111000000000000001000000000000000000000000;
		1981: Delta = 44'sb00000111111111111111000000000000000000000000;
		7782: Delta = 44'sb11110111111111111111000000000000000000000000;
		15746: Delta = 44'sb00010000000000000001000000000000000000000000;
		9729: Delta = 44'sb11110000000000000001000000000000000000000000;
		7890: Delta = 44'sb00001111111111111111000000000000000000000000;
		1873: Delta = 44'sb11101111111111111111000000000000000000000000;
		9945: Delta = 44'sb00100000000000000001000000000000000000000000;
		15530: Delta = 44'sb11100000000000000001000000000000000000000000;
		2089: Delta = 44'sb00011111111111111111000000000000000000000000;
		7674: Delta = 44'sb11011111111111111111000000000000000000000000;
		15962: Delta = 44'sb01000000000000000001000000000000000000000000;
		9513: Delta = 44'sb11000000000000000001000000000000000000000000;
		8106: Delta = 44'sb00111111111111111111000000000000000000000000;
		1657: Delta = 44'sb10111111111111111111000000000000000000000000;
		5949: Delta = 44'sb00000000000000000110000000000000000000000000;
		11670: Delta = 44'sb11111111111111111010000000000000000000000000;
		4042: Delta = 44'sb00000000000000001010000000000000000000000000;
		13577: Delta = 44'sb11111111111111110110000000000000000000000000;
		228: Delta = 44'sb00000000000000010010000000000000000000000000;
		15484: Delta = 44'sb11111111111111110010000000000000000000000000;
		2135: Delta = 44'sb00000000000000001110000000000000000000000000;
		17391: Delta = 44'sb11111111111111101110000000000000000000000000;
		10219: Delta = 44'sb00000000000000100010000000000000000000000000;
		5493: Delta = 44'sb11111111111111100010000000000000000000000000;
		12126: Delta = 44'sb00000000000000011110000000000000000000000000;
		7400: Delta = 44'sb11111111111111011110000000000000000000000000;
		12582: Delta = 44'sb00000000000001000010000000000000000000000000;
		3130: Delta = 44'sb11111111111111000010000000000000000000000000;
		14489: Delta = 44'sb00000000000000111110000000000000000000000000;
		5037: Delta = 44'sb11111111111110111110000000000000000000000000;
		17308: Delta = 44'sb00000000000010000010000000000000000000000000;
		16023: Delta = 44'sb11111111111110000010000000000000000000000000;
		1596: Delta = 44'sb00000000000001111110000000000000000000000000;
		311: Delta = 44'sb11111111111101111110000000000000000000000000;
		9141: Delta = 44'sb00000000000100000010000000000000000000000000;
		6571: Delta = 44'sb11111111111100000010000000000000000000000000;
		11048: Delta = 44'sb00000000000011111110000000000000000000000000;
		8478: Delta = 44'sb11111111111011111110000000000000000000000000;
		10426: Delta = 44'sb00000000001000000010000000000000000000000000;
		5286: Delta = 44'sb11111111111000000010000000000000000000000000;
		12333: Delta = 44'sb00000000000111111110000000000000000000000000;
		7193: Delta = 44'sb11111111110111111110000000000000000000000000;
		12996: Delta = 44'sb00000000010000000010000000000000000000000000;
		2716: Delta = 44'sb11111111110000000010000000000000000000000000;
		14903: Delta = 44'sb00000000001111111110000000000000000000000000;
		4623: Delta = 44'sb11111111101111111110000000000000000000000000;
		517: Delta = 44'sb00000000100000000010000000000000000000000000;
		15195: Delta = 44'sb11111111100000000010000000000000000000000000;
		2424: Delta = 44'sb00000000011111111110000000000000000000000000;
		17102: Delta = 44'sb11111111011111111110000000000000000000000000;
		10797: Delta = 44'sb00000001000000000010000000000000000000000000;
		4915: Delta = 44'sb11111111000000000010000000000000000000000000;
		12704: Delta = 44'sb00000000111111111110000000000000000000000000;
		6822: Delta = 44'sb11111110111111111110000000000000000000000000;
		13738: Delta = 44'sb00000010000000000010000000000000000000000000;
		1974: Delta = 44'sb11111110000000000010000000000000000000000000;
		15645: Delta = 44'sb00000001111111111110000000000000000000000000;
		3881: Delta = 44'sb11111101111111111110000000000000000000000000;
		2001: Delta = 44'sb00000100000000000010000000000000000000000000;
		13711: Delta = 44'sb11111100000000000010000000000000000000000000;
		3908: Delta = 44'sb00000011111111111110000000000000000000000000;
		15618: Delta = 44'sb11111011111111111110000000000000000000000000;
		13765: Delta = 44'sb00001000000000000010000000000000000000000000;
		1947: Delta = 44'sb11111000000000000010000000000000000000000000;
		15672: Delta = 44'sb00000111111111111110000000000000000000000000;
		3854: Delta = 44'sb11110111111111111110000000000000000000000000;
		2055: Delta = 44'sb00010000000000000010000000000000000000000000;
		13657: Delta = 44'sb11110000000000000010000000000000000000000000;
		3962: Delta = 44'sb00001111111111111110000000000000000000000000;
		15564: Delta = 44'sb11101111111111111110000000000000000000000000;
		13873: Delta = 44'sb00100000000000000010000000000000000000000000;
		1839: Delta = 44'sb11100000000000000010000000000000000000000000;
		15780: Delta = 44'sb00011111111111111110000000000000000000000000;
		3746: Delta = 44'sb11011111111111111110000000000000000000000000;
		2271: Delta = 44'sb01000000000000000010000000000000000000000000;
		13441: Delta = 44'sb11000000000000000010000000000000000000000000;
		4178: Delta = 44'sb00111111111111111110000000000000000000000000;
		15348: Delta = 44'sb10111111111111111110000000000000000000000000;
		11898: Delta = 44'sb00000000000000001100000000000000000000000000;
		5721: Delta = 44'sb11111111111111110100000000000000000000000000;
		8084: Delta = 44'sb00000000000000010100000000000000000000000000;
		9535: Delta = 44'sb11111111111111101100000000000000000000000000;
		456: Delta = 44'sb00000000000000100100000000000000000000000000;
		13349: Delta = 44'sb11111111111111100100000000000000000000000000;
		4270: Delta = 44'sb00000000000000011100000000000000000000000000;
		17163: Delta = 44'sb11111111111111011100000000000000000000000000;
		2819: Delta = 44'sb00000000000001000100000000000000000000000000;
		10986: Delta = 44'sb11111111111111000100000000000000000000000000;
		6633: Delta = 44'sb00000000000000111100000000000000000000000000;
		14800: Delta = 44'sb11111111111110111100000000000000000000000000;
		7545: Delta = 44'sb00000000000010000100000000000000000000000000;
		6260: Delta = 44'sb11111111111110000100000000000000000000000000;
		11359: Delta = 44'sb00000000000001111100000000000000000000000000;
		10074: Delta = 44'sb11111111111101111100000000000000000000000000;
		16997: Delta = 44'sb00000000000100000100000000000000000000000000;
		14427: Delta = 44'sb11111111111100000100000000000000000000000000;
		3192: Delta = 44'sb00000000000011111100000000000000000000000000;
		622: Delta = 44'sb11111111111011111100000000000000000000000000;
		663: Delta = 44'sb00000000001000000100000000000000000000000000;
		13142: Delta = 44'sb11111111111000000100000000000000000000000000;
		4477: Delta = 44'sb00000000000111111100000000000000000000000000;
		16956: Delta = 44'sb11111111110111111100000000000000000000000000;
		3233: Delta = 44'sb00000000010000000100000000000000000000000000;
		10572: Delta = 44'sb11111111110000000100000000000000000000000000;
		7047: Delta = 44'sb00000000001111111100000000000000000000000000;
		14386: Delta = 44'sb11111111101111111100000000000000000000000000;
		8373: Delta = 44'sb00000000100000000100000000000000000000000000;
		5432: Delta = 44'sb11111111100000000100000000000000000000000000;
		12187: Delta = 44'sb00000000011111111100000000000000000000000000;
		9246: Delta = 44'sb11111111011111111100000000000000000000000000;
		1034: Delta = 44'sb00000001000000000100000000000000000000000000;
		12771: Delta = 44'sb11111111000000000100000000000000000000000000;
		4848: Delta = 44'sb00000000111111111100000000000000000000000000;
		16585: Delta = 44'sb11111110111111111100000000000000000000000000;
		3975: Delta = 44'sb00000010000000000100000000000000000000000000;
		9830: Delta = 44'sb11111110000000000100000000000000000000000000;
		7789: Delta = 44'sb00000001111111111100000000000000000000000000;
		13644: Delta = 44'sb11111101111111111100000000000000000000000000;
		9857: Delta = 44'sb00000100000000000100000000000000000000000000;
		3948: Delta = 44'sb11111100000000000100000000000000000000000000;
		13671: Delta = 44'sb00000011111111111100000000000000000000000000;
		7762: Delta = 44'sb11111011111111111100000000000000000000000000;
		4002: Delta = 44'sb00001000000000000100000000000000000000000000;
		9803: Delta = 44'sb11111000000000000100000000000000000000000000;
		7816: Delta = 44'sb00000111111111111100000000000000000000000000;
		13617: Delta = 44'sb11110111111111111100000000000000000000000000;
		9911: Delta = 44'sb00010000000000000100000000000000000000000000;
		3894: Delta = 44'sb11110000000000000100000000000000000000000000;
		13725: Delta = 44'sb00001111111111111100000000000000000000000000;
		7708: Delta = 44'sb11101111111111111100000000000000000000000000;
		4110: Delta = 44'sb00100000000000000100000000000000000000000000;
		9695: Delta = 44'sb11100000000000000100000000000000000000000000;
		7924: Delta = 44'sb00011111111111111100000000000000000000000000;
		13509: Delta = 44'sb11011111111111111100000000000000000000000000;
		10127: Delta = 44'sb01000000000000000100000000000000000000000000;
		3678: Delta = 44'sb11000000000000000100000000000000000000000000;
		13941: Delta = 44'sb00111111111111111100000000000000000000000000;
		7492: Delta = 44'sb10111111111111111100000000000000000000000000;
		6177: Delta = 44'sb00000000000000011000000000000000000000000000;
		11442: Delta = 44'sb11111111111111101000000000000000000000000000;
		16168: Delta = 44'sb00000000000000101000000000000000000000000000;
		1451: Delta = 44'sb11111111111111011000000000000000000000000000;
		912: Delta = 44'sb00000000000001001000000000000000000000000000;
		9079: Delta = 44'sb11111111111111001000000000000000000000000000;
		8540: Delta = 44'sb00000000000000111000000000000000000000000000;
		16707: Delta = 44'sb11111111111110111000000000000000000000000000;
		5638: Delta = 44'sb00000000000010001000000000000000000000000000;
		4353: Delta = 44'sb11111111111110001000000000000000000000000000;
		13266: Delta = 44'sb00000000000001111000000000000000000000000000;
		11981: Delta = 44'sb11111111111101111000000000000000000000000000;
		15090: Delta = 44'sb00000000000100001000000000000000000000000000;
		12520: Delta = 44'sb11111111111100001000000000000000000000000000;
		5099: Delta = 44'sb00000000000011111000000000000000000000000000;
		2529: Delta = 44'sb11111111111011111000000000000000000000000000;
		16375: Delta = 44'sb00000000001000001000000000000000000000000000;
		11235: Delta = 44'sb11111111111000001000000000000000000000000000;
		6384: Delta = 44'sb00000000000111111000000000000000000000000000;
		1244: Delta = 44'sb11111111110111111000000000000000000000000000;
		1326: Delta = 44'sb00000000010000001000000000000000000000000000;
		8665: Delta = 44'sb11111111110000001000000000000000000000000000;
		8954: Delta = 44'sb00000000001111111000000000000000000000000000;
		16293: Delta = 44'sb11111111101111111000000000000000000000000000;
		6466: Delta = 44'sb00000000100000001000000000000000000000000000;
		3525: Delta = 44'sb11111111100000001000000000000000000000000000;
		14094: Delta = 44'sb00000000011111111000000000000000000000000000;
		11153: Delta = 44'sb11111111011111111000000000000000000000000000;
		16746: Delta = 44'sb00000001000000001000000000000000000000000000;
		10864: Delta = 44'sb11111111000000001000000000000000000000000000;
		6755: Delta = 44'sb00000000111111111000000000000000000000000000;
		873: Delta = 44'sb11111110111111111000000000000000000000000000;
		2068: Delta = 44'sb00000010000000001000000000000000000000000000;
		7923: Delta = 44'sb11111110000000001000000000000000000000000000;
		9696: Delta = 44'sb00000001111111111000000000000000000000000000;
		15551: Delta = 44'sb11111101111111111000000000000000000000000000;
		7950: Delta = 44'sb00000100000000001000000000000000000000000000;
		2041: Delta = 44'sb11111100000000001000000000000000000000000000;
		15578: Delta = 44'sb00000011111111111000000000000000000000000000;
		9669: Delta = 44'sb11111011111111111000000000000000000000000000;
		2095: Delta = 44'sb00001000000000001000000000000000000000000000;
		7896: Delta = 44'sb11111000000000001000000000000000000000000000;
		9723: Delta = 44'sb00000111111111111000000000000000000000000000;
		15524: Delta = 44'sb11110111111111111000000000000000000000000000;
		8004: Delta = 44'sb00010000000000001000000000000000000000000000;
		1987: Delta = 44'sb11110000000000001000000000000000000000000000;
		15632: Delta = 44'sb00001111111111111000000000000000000000000000;
		9615: Delta = 44'sb11101111111111111000000000000000000000000000;
		2203: Delta = 44'sb00100000000000001000000000000000000000000000;
		7788: Delta = 44'sb11100000000000001000000000000000000000000000;
		9831: Delta = 44'sb00011111111111111000000000000000000000000000;
		15416: Delta = 44'sb11011111111111111000000000000000000000000000;
		8220: Delta = 44'sb01000000000000001000000000000000000000000000;
		1771: Delta = 44'sb11000000000000001000000000000000000000000000;
		15848: Delta = 44'sb00111111111111111000000000000000000000000000;
		9399: Delta = 44'sb10111111111111111000000000000000000000000000;
		12354: Delta = 44'sb00000000000000110000000000000000000000000000;
		5265: Delta = 44'sb11111111111111010000000000000000000000000000;
		14717: Delta = 44'sb00000000000001010000000000000000000000000000;
		2902: Delta = 44'sb11111111111110110000000000000000000000000000;
		1824: Delta = 44'sb00000000000010010000000000000000000000000000;
		539: Delta = 44'sb11111111111110010000000000000000000000000000;
		17080: Delta = 44'sb00000000000001110000000000000000000000000000;
		15795: Delta = 44'sb11111111111101110000000000000000000000000000;
		11276: Delta = 44'sb00000000000100010000000000000000000000000000;
		8706: Delta = 44'sb11111111111100010000000000000000000000000000;
		8913: Delta = 44'sb00000000000011110000000000000000000000000000;
		6343: Delta = 44'sb11111111111011110000000000000000000000000000;
		12561: Delta = 44'sb00000000001000010000000000000000000000000000;
		7421: Delta = 44'sb11111111111000010000000000000000000000000000;
		10198: Delta = 44'sb00000000000111110000000000000000000000000000;
		5058: Delta = 44'sb11111111110111110000000000000000000000000000;
		15131: Delta = 44'sb00000000010000010000000000000000000000000000;
		4851: Delta = 44'sb11111111110000010000000000000000000000000000;
		12768: Delta = 44'sb00000000001111110000000000000000000000000000;
		2488: Delta = 44'sb11111111101111110000000000000000000000000000;
		2652: Delta = 44'sb00000000100000010000000000000000000000000000;
		17330: Delta = 44'sb11111111100000010000000000000000000000000000;
		289: Delta = 44'sb00000000011111110000000000000000000000000000;
		14967: Delta = 44'sb11111111011111110000000000000000000000000000;
		12932: Delta = 44'sb00000001000000010000000000000000000000000000;
		7050: Delta = 44'sb11111111000000010000000000000000000000000000;
		10569: Delta = 44'sb00000000111111110000000000000000000000000000;
		4687: Delta = 44'sb11111110111111110000000000000000000000000000;
		15873: Delta = 44'sb00000010000000010000000000000000000000000000;
		4109: Delta = 44'sb11111110000000010000000000000000000000000000;
		13510: Delta = 44'sb00000001111111110000000000000000000000000000;
		1746: Delta = 44'sb11111101111111110000000000000000000000000000;
		4136: Delta = 44'sb00000100000000010000000000000000000000000000;
		15846: Delta = 44'sb11111100000000010000000000000000000000000000;
		1773: Delta = 44'sb00000011111111110000000000000000000000000000;
		13483: Delta = 44'sb11111011111111110000000000000000000000000000;
		15900: Delta = 44'sb00001000000000010000000000000000000000000000;
		4082: Delta = 44'sb11111000000000010000000000000000000000000000;
		13537: Delta = 44'sb00000111111111110000000000000000000000000000;
		1719: Delta = 44'sb11110111111111110000000000000000000000000000;
		4190: Delta = 44'sb00010000000000010000000000000000000000000000;
		15792: Delta = 44'sb11110000000000010000000000000000000000000000;
		1827: Delta = 44'sb00001111111111110000000000000000000000000000;
		13429: Delta = 44'sb11101111111111110000000000000000000000000000;
		16008: Delta = 44'sb00100000000000010000000000000000000000000000;
		3974: Delta = 44'sb11100000000000010000000000000000000000000000;
		13645: Delta = 44'sb00011111111111110000000000000000000000000000;
		1611: Delta = 44'sb11011111111111110000000000000000000000000000;
		4406: Delta = 44'sb01000000000000010000000000000000000000000000;
		15576: Delta = 44'sb11000000000000010000000000000000000000000000;
		2043: Delta = 44'sb00111111111111110000000000000000000000000000;
		13213: Delta = 44'sb10111111111111110000000000000000000000000000;
		7089: Delta = 44'sb00000000000001100000000000000000000000000000;
		10530: Delta = 44'sb11111111111110100000000000000000000000000000;
		11815: Delta = 44'sb00000000000010100000000000000000000000000000;
		5804: Delta = 44'sb11111111111101100000000000000000000000000000;
		3648: Delta = 44'sb00000000000100100000000000000000000000000000;
		1078: Delta = 44'sb11111111111100100000000000000000000000000000;
		16541: Delta = 44'sb00000000000011100000000000000000000000000000;
		13971: Delta = 44'sb11111111111011100000000000000000000000000000;
		4933: Delta = 44'sb00000000001000100000000000000000000000000000;
		17412: Delta = 44'sb11111111111000100000000000000000000000000000;
		207: Delta = 44'sb00000000000111100000000000000000000000000000;
		12686: Delta = 44'sb11111111110111100000000000000000000000000000;
		7503: Delta = 44'sb00000000010000100000000000000000000000000000;
		14842: Delta = 44'sb11111111110000100000000000000000000000000000;
		2777: Delta = 44'sb00000000001111100000000000000000000000000000;
		10116: Delta = 44'sb11111111101111100000000000000000000000000000;
		12643: Delta = 44'sb00000000100000100000000000000000000000000000;
		9702: Delta = 44'sb11111111100000100000000000000000000000000000;
		7917: Delta = 44'sb00000000011111100000000000000000000000000000;
		4976: Delta = 44'sb11111111011111100000000000000000000000000000;
		5304: Delta = 44'sb00000001000000100000000000000000000000000000;
		17041: Delta = 44'sb11111111000000100000000000000000000000000000;
		578: Delta = 44'sb00000000111111100000000000000000000000000000;
		12315: Delta = 44'sb11111110111111100000000000000000000000000000;
		8245: Delta = 44'sb00000010000000100000000000000000000000000000;
		14100: Delta = 44'sb11111110000000100000000000000000000000000000;
		3519: Delta = 44'sb00000001111111100000000000000000000000000000;
		9374: Delta = 44'sb11111101111111100000000000000000000000000000;
		14127: Delta = 44'sb00000100000000100000000000000000000000000000;
		8218: Delta = 44'sb11111100000000100000000000000000000000000000;
		9401: Delta = 44'sb00000011111111100000000000000000000000000000;
		3492: Delta = 44'sb11111011111111100000000000000000000000000000;
		8272: Delta = 44'sb00001000000000100000000000000000000000000000;
		14073: Delta = 44'sb11111000000000100000000000000000000000000000;
		3546: Delta = 44'sb00000111111111100000000000000000000000000000;
		9347: Delta = 44'sb11110111111111100000000000000000000000000000;
		14181: Delta = 44'sb00010000000000100000000000000000000000000000;
		8164: Delta = 44'sb11110000000000100000000000000000000000000000;
		9455: Delta = 44'sb00001111111111100000000000000000000000000000;
		3438: Delta = 44'sb11101111111111100000000000000000000000000000;
		8380: Delta = 44'sb00100000000000100000000000000000000000000000;
		13965: Delta = 44'sb11100000000000100000000000000000000000000000;
		3654: Delta = 44'sb00011111111111100000000000000000000000000000;
		9239: Delta = 44'sb11011111111111100000000000000000000000000000;
		14397: Delta = 44'sb01000000000000100000000000000000000000000000;
		7948: Delta = 44'sb11000000000000100000000000000000000000000000;
		9671: Delta = 44'sb00111111111111100000000000000000000000000000;
		3222: Delta = 44'sb10111111111111100000000000000000000000000000;
		14178: Delta = 44'sb00000000000011000000000000000000000000000000;
		3441: Delta = 44'sb11111111111101000000000000000000000000000000;
		6011: Delta = 44'sb00000000000101000000000000000000000000000000;
		11608: Delta = 44'sb11111111111011000000000000000000000000000000;
		7296: Delta = 44'sb00000000001001000000000000000000000000000000;
		2156: Delta = 44'sb11111111111001000000000000000000000000000000;
		15463: Delta = 44'sb00000000000111000000000000000000000000000000;
		10323: Delta = 44'sb11111111110111000000000000000000000000000000;
		9866: Delta = 44'sb00000000010001000000000000000000000000000000;
		17205: Delta = 44'sb11111111110001000000000000000000000000000000;
		414: Delta = 44'sb00000000001111000000000000000000000000000000;
		7753: Delta = 44'sb11111111101111000000000000000000000000000000;
		15006: Delta = 44'sb00000000100001000000000000000000000000000000;
		12065: Delta = 44'sb11111111100001000000000000000000000000000000;
		5554: Delta = 44'sb00000000011111000000000000000000000000000000;
		2613: Delta = 44'sb11111111011111000000000000000000000000000000;
		7667: Delta = 44'sb00000001000001000000000000000000000000000000;
		1785: Delta = 44'sb11111111000001000000000000000000000000000000;
		15834: Delta = 44'sb00000000111111000000000000000000000000000000;
		9952: Delta = 44'sb11111110111111000000000000000000000000000000;
		10608: Delta = 44'sb00000010000001000000000000000000000000000000;
		16463: Delta = 44'sb11111110000001000000000000000000000000000000;
		1156: Delta = 44'sb00000001111111000000000000000000000000000000;
		7011: Delta = 44'sb11111101111111000000000000000000000000000000;
		16490: Delta = 44'sb00000100000001000000000000000000000000000000;
		10581: Delta = 44'sb11111100000001000000000000000000000000000000;
		7038: Delta = 44'sb00000011111111000000000000000000000000000000;
		1129: Delta = 44'sb11111011111111000000000000000000000000000000;
		10635: Delta = 44'sb00001000000001000000000000000000000000000000;
		16436: Delta = 44'sb11111000000001000000000000000000000000000000;
		1183: Delta = 44'sb00000111111111000000000000000000000000000000;
		6984: Delta = 44'sb11110111111111000000000000000000000000000000;
		16544: Delta = 44'sb00010000000001000000000000000000000000000000;
		10527: Delta = 44'sb11110000000001000000000000000000000000000000;
		7092: Delta = 44'sb00001111111111000000000000000000000000000000;
		1075: Delta = 44'sb11101111111111000000000000000000000000000000;
		10743: Delta = 44'sb00100000000001000000000000000000000000000000;
		16328: Delta = 44'sb11100000000001000000000000000000000000000000;
		1291: Delta = 44'sb00011111111111000000000000000000000000000000;
		6876: Delta = 44'sb11011111111111000000000000000000000000000000;
		16760: Delta = 44'sb01000000000001000000000000000000000000000000;
		10311: Delta = 44'sb11000000000001000000000000000000000000000000;
		7308: Delta = 44'sb00111111111111000000000000000000000000000000;
		859: Delta = 44'sb10111111111111000000000000000000000000000000;
		10737: Delta = 44'sb00000000000110000000000000000000000000000000;
		6882: Delta = 44'sb11111111111010000000000000000000000000000000;
		12022: Delta = 44'sb00000000001010000000000000000000000000000000;
		5597: Delta = 44'sb11111111110110000000000000000000000000000000;
		14592: Delta = 44'sb00000000010010000000000000000000000000000000;
		4312: Delta = 44'sb11111111110010000000000000000000000000000000;
		13307: Delta = 44'sb00000000001110000000000000000000000000000000;
		3027: Delta = 44'sb11111111101110000000000000000000000000000000;
		2113: Delta = 44'sb00000000100010000000000000000000000000000000;
		16791: Delta = 44'sb11111111100010000000000000000000000000000000;
		828: Delta = 44'sb00000000011110000000000000000000000000000000;
		15506: Delta = 44'sb11111111011110000000000000000000000000000000;
		12393: Delta = 44'sb00000001000010000000000000000000000000000000;
		6511: Delta = 44'sb11111111000010000000000000000000000000000000;
		11108: Delta = 44'sb00000000111110000000000000000000000000000000;
		5226: Delta = 44'sb11111110111110000000000000000000000000000000;
		15334: Delta = 44'sb00000010000010000000000000000000000000000000;
		3570: Delta = 44'sb11111110000010000000000000000000000000000000;
		14049: Delta = 44'sb00000001111110000000000000000000000000000000;
		2285: Delta = 44'sb11111101111110000000000000000000000000000000;
		3597: Delta = 44'sb00000100000010000000000000000000000000000000;
		15307: Delta = 44'sb11111100000010000000000000000000000000000000;
		2312: Delta = 44'sb00000011111110000000000000000000000000000000;
		14022: Delta = 44'sb11111011111110000000000000000000000000000000;
		15361: Delta = 44'sb00001000000010000000000000000000000000000000;
		3543: Delta = 44'sb11111000000010000000000000000000000000000000;
		14076: Delta = 44'sb00000111111110000000000000000000000000000000;
		2258: Delta = 44'sb11110111111110000000000000000000000000000000;
		3651: Delta = 44'sb00010000000010000000000000000000000000000000;
		15253: Delta = 44'sb11110000000010000000000000000000000000000000;
		2366: Delta = 44'sb00001111111110000000000000000000000000000000;
		13968: Delta = 44'sb11101111111110000000000000000000000000000000;
		15469: Delta = 44'sb00100000000010000000000000000000000000000000;
		3435: Delta = 44'sb11100000000010000000000000000000000000000000;
		14184: Delta = 44'sb00011111111110000000000000000000000000000000;
		2150: Delta = 44'sb11011111111110000000000000000000000000000000;
		3867: Delta = 44'sb01000000000010000000000000000000000000000000;
		15037: Delta = 44'sb11000000000010000000000000000000000000000000;
		2582: Delta = 44'sb00111111111110000000000000000000000000000000;
		13752: Delta = 44'sb10111111111110000000000000000000000000000000;
		3855: Delta = 44'sb00000000001100000000000000000000000000000000;
		13764: Delta = 44'sb11111111110100000000000000000000000000000000;
		6425: Delta = 44'sb00000000010100000000000000000000000000000000;
		11194: Delta = 44'sb11111111101100000000000000000000000000000000;
		11565: Delta = 44'sb00000000100100000000000000000000000000000000;
		8624: Delta = 44'sb11111111100100000000000000000000000000000000;
		8995: Delta = 44'sb00000000011100000000000000000000000000000000;
		6054: Delta = 44'sb11111111011100000000000000000000000000000000;
		4226: Delta = 44'sb00000001000100000000000000000000000000000000;
		15963: Delta = 44'sb11111111000100000000000000000000000000000000;
		1656: Delta = 44'sb00000000111100000000000000000000000000000000;
		13393: Delta = 44'sb11111110111100000000000000000000000000000000;
		7167: Delta = 44'sb00000010000100000000000000000000000000000000;
		13022: Delta = 44'sb11111110000100000000000000000000000000000000;
		4597: Delta = 44'sb00000001111100000000000000000000000000000000;
		10452: Delta = 44'sb11111101111100000000000000000000000000000000;
		13049: Delta = 44'sb00000100000100000000000000000000000000000000;
		7140: Delta = 44'sb11111100000100000000000000000000000000000000;
		10479: Delta = 44'sb00000011111100000000000000000000000000000000;
		4570: Delta = 44'sb11111011111100000000000000000000000000000000;
		7194: Delta = 44'sb00001000000100000000000000000000000000000000;
		12995: Delta = 44'sb11111000000100000000000000000000000000000000;
		4624: Delta = 44'sb00000111111100000000000000000000000000000000;
		10425: Delta = 44'sb11110111111100000000000000000000000000000000;
		13103: Delta = 44'sb00010000000100000000000000000000000000000000;
		7086: Delta = 44'sb11110000000100000000000000000000000000000000;
		10533: Delta = 44'sb00001111111100000000000000000000000000000000;
		4516: Delta = 44'sb11101111111100000000000000000000000000000000;
		7302: Delta = 44'sb00100000000100000000000000000000000000000000;
		12887: Delta = 44'sb11100000000100000000000000000000000000000000;
		4732: Delta = 44'sb00011111111100000000000000000000000000000000;
		10317: Delta = 44'sb11011111111100000000000000000000000000000000;
		13319: Delta = 44'sb01000000000100000000000000000000000000000000;
		6870: Delta = 44'sb11000000000100000000000000000000000000000000;
		10749: Delta = 44'sb00111111111100000000000000000000000000000000;
		4300: Delta = 44'sb10111111111100000000000000000000000000000000;
		7710: Delta = 44'sb00000000011000000000000000000000000000000000;
		9909: Delta = 44'sb11111111101000000000000000000000000000000000;
		12850: Delta = 44'sb00000000101000000000000000000000000000000000;
		4769: Delta = 44'sb11111111011000000000000000000000000000000000;
		5511: Delta = 44'sb00000001001000000000000000000000000000000000;
		17248: Delta = 44'sb11111111001000000000000000000000000000000000;
		371: Delta = 44'sb00000000111000000000000000000000000000000000;
		12108: Delta = 44'sb11111110111000000000000000000000000000000000;
		8452: Delta = 44'sb00000010001000000000000000000000000000000000;
		14307: Delta = 44'sb11111110001000000000000000000000000000000000;
		3312: Delta = 44'sb00000001111000000000000000000000000000000000;
		9167: Delta = 44'sb11111101111000000000000000000000000000000000;
		14334: Delta = 44'sb00000100001000000000000000000000000000000000;
		8425: Delta = 44'sb11111100001000000000000000000000000000000000;
		9194: Delta = 44'sb00000011111000000000000000000000000000000000;
		3285: Delta = 44'sb11111011111000000000000000000000000000000000;
		8479: Delta = 44'sb00001000001000000000000000000000000000000000;
		14280: Delta = 44'sb11111000001000000000000000000000000000000000;
		3339: Delta = 44'sb00000111111000000000000000000000000000000000;
		9140: Delta = 44'sb11110111111000000000000000000000000000000000;
		14388: Delta = 44'sb00010000001000000000000000000000000000000000;
		8371: Delta = 44'sb11110000001000000000000000000000000000000000;
		9248: Delta = 44'sb00001111111000000000000000000000000000000000;
		3231: Delta = 44'sb11101111111000000000000000000000000000000000;
		8587: Delta = 44'sb00100000001000000000000000000000000000000000;
		14172: Delta = 44'sb11100000001000000000000000000000000000000000;
		3447: Delta = 44'sb00011111111000000000000000000000000000000000;
		9032: Delta = 44'sb11011111111000000000000000000000000000000000;
		14604: Delta = 44'sb01000000001000000000000000000000000000000000;
		8155: Delta = 44'sb11000000001000000000000000000000000000000000;
		9464: Delta = 44'sb00111111111000000000000000000000000000000000;
		3015: Delta = 44'sb10111111111000000000000000000000000000000000;
		15420: Delta = 44'sb00000000110000000000000000000000000000000000;
		2199: Delta = 44'sb11111111010000000000000000000000000000000000;
		8081: Delta = 44'sb00000001010000000000000000000000000000000000;
		9538: Delta = 44'sb11111110110000000000000000000000000000000000;
		11022: Delta = 44'sb00000010010000000000000000000000000000000000;
		16877: Delta = 44'sb11111110010000000000000000000000000000000000;
		742: Delta = 44'sb00000001110000000000000000000000000000000000;
		6597: Delta = 44'sb11111101110000000000000000000000000000000000;
		16904: Delta = 44'sb00000100010000000000000000000000000000000000;
		10995: Delta = 44'sb11111100010000000000000000000000000000000000;
		6624: Delta = 44'sb00000011110000000000000000000000000000000000;
		715: Delta = 44'sb11111011110000000000000000000000000000000000;
		11049: Delta = 44'sb00001000010000000000000000000000000000000000;
		16850: Delta = 44'sb11111000010000000000000000000000000000000000;
		769: Delta = 44'sb00000111110000000000000000000000000000000000;
		6570: Delta = 44'sb11110111110000000000000000000000000000000000;
		16958: Delta = 44'sb00010000010000000000000000000000000000000000;
		10941: Delta = 44'sb11110000010000000000000000000000000000000000;
		6678: Delta = 44'sb00001111110000000000000000000000000000000000;
		661: Delta = 44'sb11101111110000000000000000000000000000000000;
		11157: Delta = 44'sb00100000010000000000000000000000000000000000;
		16742: Delta = 44'sb11100000010000000000000000000000000000000000;
		877: Delta = 44'sb00011111110000000000000000000000000000000000;
		6462: Delta = 44'sb11011111110000000000000000000000000000000000;
		17174: Delta = 44'sb01000000010000000000000000000000000000000000;
		10725: Delta = 44'sb11000000010000000000000000000000000000000000;
		6894: Delta = 44'sb00111111110000000000000000000000000000000000;
		445: Delta = 44'sb10111111110000000000000000000000000000000000;
		13221: Delta = 44'sb00000001100000000000000000000000000000000000;
		4398: Delta = 44'sb11111110100000000000000000000000000000000000;
		16162: Delta = 44'sb00000010100000000000000000000000000000000000;
		1457: Delta = 44'sb11111101100000000000000000000000000000000000;
		4425: Delta = 44'sb00000100100000000000000000000000000000000000;
		16135: Delta = 44'sb11111100100000000000000000000000000000000000;
		1484: Delta = 44'sb00000011100000000000000000000000000000000000;
		13194: Delta = 44'sb11111011100000000000000000000000000000000000;
		16189: Delta = 44'sb00001000100000000000000000000000000000000000;
		4371: Delta = 44'sb11111000100000000000000000000000000000000000;
		13248: Delta = 44'sb00000111100000000000000000000000000000000000;
		1430: Delta = 44'sb11110111100000000000000000000000000000000000;
		4479: Delta = 44'sb00010000100000000000000000000000000000000000;
		16081: Delta = 44'sb11110000100000000000000000000000000000000000;
		1538: Delta = 44'sb00001111100000000000000000000000000000000000;
		13140: Delta = 44'sb11101111100000000000000000000000000000000000;
		16297: Delta = 44'sb00100000100000000000000000000000000000000000;
		4263: Delta = 44'sb11100000100000000000000000000000000000000000;
		13356: Delta = 44'sb00011111100000000000000000000000000000000000;
		1322: Delta = 44'sb11011111100000000000000000000000000000000000;
		4695: Delta = 44'sb01000000100000000000000000000000000000000000;
		15865: Delta = 44'sb11000000100000000000000000000000000000000000;
		1754: Delta = 44'sb00111111100000000000000000000000000000000000;
		12924: Delta = 44'sb10111111100000000000000000000000000000000000;
		8823: Delta = 44'sb00000011000000000000000000000000000000000000;
		8796: Delta = 44'sb11111101000000000000000000000000000000000000;
		14705: Delta = 44'sb00000101000000000000000000000000000000000000;
		2914: Delta = 44'sb11111011000000000000000000000000000000000000;
		8850: Delta = 44'sb00001001000000000000000000000000000000000000;
		14651: Delta = 44'sb11111001000000000000000000000000000000000000;
		2968: Delta = 44'sb00000111000000000000000000000000000000000000;
		8769: Delta = 44'sb11110111000000000000000000000000000000000000;
		14759: Delta = 44'sb00010001000000000000000000000000000000000000;
		8742: Delta = 44'sb11110001000000000000000000000000000000000000;
		8877: Delta = 44'sb00001111000000000000000000000000000000000000;
		2860: Delta = 44'sb11101111000000000000000000000000000000000000;
		8958: Delta = 44'sb00100001000000000000000000000000000000000000;
		14543: Delta = 44'sb11100001000000000000000000000000000000000000;
		3076: Delta = 44'sb00011111000000000000000000000000000000000000;
		8661: Delta = 44'sb11011111000000000000000000000000000000000000;
		14975: Delta = 44'sb01000001000000000000000000000000000000000000;
		8526: Delta = 44'sb11000001000000000000000000000000000000000000;
		9093: Delta = 44'sb00111111000000000000000000000000000000000000;
		2644: Delta = 44'sb10111111000000000000000000000000000000000000;
		27: Delta = 44'sb00000110000000000000000000000000000000000000;
		17592: Delta = 44'sb11111010000000000000000000000000000000000000;
		11791: Delta = 44'sb00001010000000000000000000000000000000000000;
		5828: Delta = 44'sb11110110000000000000000000000000000000000000;
		81: Delta = 44'sb00010010000000000000000000000000000000000000;
		11683: Delta = 44'sb11110010000000000000000000000000000000000000;
		5936: Delta = 44'sb00001110000000000000000000000000000000000000;
		17538: Delta = 44'sb11101110000000000000000000000000000000000000;
		11899: Delta = 44'sb00100010000000000000000000000000000000000000;
		17484: Delta = 44'sb11100010000000000000000000000000000000000000;
		135: Delta = 44'sb00011110000000000000000000000000000000000000;
		5720: Delta = 44'sb11011110000000000000000000000000000000000000;
		297: Delta = 44'sb01000010000000000000000000000000000000000000;
		11467: Delta = 44'sb11000010000000000000000000000000000000000000;
		6152: Delta = 44'sb00111110000000000000000000000000000000000000;
		17322: Delta = 44'sb10111110000000000000000000000000000000000000;
		54: Delta = 44'sb00001100000000000000000000000000000000000000;
		17565: Delta = 44'sb11110100000000000000000000000000000000000000;
		5963: Delta = 44'sb00010100000000000000000000000000000000000000;
		11656: Delta = 44'sb11101100000000000000000000000000000000000000;
		162: Delta = 44'sb00100100000000000000000000000000000000000000;
		5747: Delta = 44'sb11100100000000000000000000000000000000000000;
		11872: Delta = 44'sb00011100000000000000000000000000000000000000;
		17457: Delta = 44'sb11011100000000000000000000000000000000000000;
		6179: Delta = 44'sb01000100000000000000000000000000000000000000;
		17349: Delta = 44'sb11000100000000000000000000000000000000000000;
		270: Delta = 44'sb00111100000000000000000000000000000000000000;
		11440: Delta = 44'sb10111100000000000000000000000000000000000000;
		108: Delta = 44'sb00011000000000000000000000000000000000000000;
		17511: Delta = 44'sb11101000000000000000000000000000000000000000;
		11926: Delta = 44'sb00101000000000000000000000000000000000000000;
		5693: Delta = 44'sb11011000000000000000000000000000000000000000;
		324: Delta = 44'sb01001000000000000000000000000000000000000000;
		11494: Delta = 44'sb11001000000000000000000000000000000000000000;
		6125: Delta = 44'sb00111000000000000000000000000000000000000000;
		17295: Delta = 44'sb10111000000000000000000000000000000000000000;
		216: Delta = 44'sb00110000000000000000000000000000000000000000;
		17403: Delta = 44'sb11010000000000000000000000000000000000000000;
		6233: Delta = 44'sb01010000000000000000000000000000000000000000;
		11386: Delta = 44'sb10110000000000000000000000000000000000000000;
		432: Delta = 44'sb01100000000000000000000000000000000000000000;
		17187: Delta = 44'sb10100000000000000000000000000000000000000000;
		default: Delta =44'sb0;
	endcase
end

assign N = (W - Delta) / A;

endmodule

// Product (AN) Code SEC l-LUT
// SEC_lLUT24bits.v
// Received single error location l, output remainder r.
module SEC_lLUT24bits(l, r);
input	signed	[6:0]	l;
output	reg	[13:0]	r;
always@(*) begin
	case(l)
		1: r = 1;
		-1: r = 13836;
		2: r = 2;
		-2: r = 13835;
		3: r = 4;
		-3: r = 13833;
		4: r = 8;
		-4: r = 13829;
		5: r = 16;
		-5: r = 13821;
		6: r = 32;
		-6: r = 13805;
		7: r = 64;
		-7: r = 13773;
		8: r = 128;
		-8: r = 13709;
		9: r = 256;
		-9: r = 13581;
		10: r = 512;
		-10: r = 13325;
		11: r = 1024;
		-11: r = 12813;
		12: r = 2048;
		-12: r = 11789;
		13: r = 4096;
		-13: r = 9741;
		14: r = 8192;
		-14: r = 5645;
		15: r = 2547;
		-15: r = 11290;
		16: r = 5094;
		-16: r = 8743;
		17: r = 10188;
		-17: r = 3649;
		18: r = 6539;
		-18: r = 7298;
		19: r = 13078;
		-19: r = 759;
		20: r = 12319;
		-20: r = 1518;
		21: r = 10801;
		-21: r = 3036;
		22: r = 7765;
		-22: r = 6072;
		23: r = 1693;
		-23: r = 12144;
		24: r = 3386;
		-24: r = 10451;
		25: r = 6772;
		-25: r = 7065;
		26: r = 13544;
		-26: r = 293;
		27: r = 13251;
		-27: r = 586;
		28: r = 12665;
		-28: r = 1172;
		29: r = 11493;
		-29: r = 2344;
		30: r = 9149;
		-30: r = 4688;
		31: r = 4461;
		-31: r = 9376;
		32: r = 8922;
		-32: r = 4915;
		33: r = 4007;
		-33: r = 9830;
		34: r = 8014;
		-34: r = 5823;
		35: r = 2191;
		-35: r = 11646;
		36: r = 4382;
		-36: r = 9455;
		37: r = 8764;
		-37: r = 5073;
		38: r = 3691;
		-38: r = 10146;
		default: r = 0;
	endcase
end

endmodule

// Product (AN) Code DEC r-LUT
// DEC_rLUT12bits.v
// Used to do DEC, but corrected errors by locations, not AWE
// Received remainder r, output two error locations.
module DEC_rLUT12bits(r, l_1, l_2);
input 	[11:0]	r;
output	reg	signed	[5:0]	l_1;
output	reg	signed	[5:0]	l_2;
always@(*) begin
	case(r)
		1: begin l_1 = -1;
				 l_2 = +2; end
		3348: begin l_1 = +1;
				 l_2 = -2; end
		2: begin l_1 = +1;
				 l_2 = +1; end
		3347: begin l_1 = -1;
				 l_2 = -1; end
		4: begin l_1 = +2;
				 l_2 = +2; end
		3345: begin l_1 = -2;
				 l_2 = -2; end
		8: begin l_1 = +3;
				 l_2 = +3; end
		3341: begin l_1 = -3;
				 l_2 = -3; end
		16: begin l_1 = +4;
				 l_2 = +4; end
		3333: begin l_1 = -4;
				 l_2 = -4; end
		32: begin l_1 = +5;
				 l_2 = +5; end
		3317: begin l_1 = -5;
				 l_2 = -5; end
		64: begin l_1 = +6;
				 l_2 = +6; end
		3285: begin l_1 = -6;
				 l_2 = -6; end
		128: begin l_1 = +7;
				 l_2 = +7; end
		3221: begin l_1 = -7;
				 l_2 = -7; end
		256: begin l_1 = +8;
				 l_2 = +8; end
		3093: begin l_1 = -8;
				 l_2 = -8; end
		512: begin l_1 = +9;
				 l_2 = +9; end
		2837: begin l_1 = -9;
				 l_2 = -9; end
		1024: begin l_1 = +10;
				 l_2 = +10; end
		2325: begin l_1 = -10;
				 l_2 = -10; end
		2048: begin l_1 = +11;
				 l_2 = +11; end
		1301: begin l_1 = -11;
				 l_2 = -11; end
		747: begin l_1 = +12;
				 l_2 = +12; end
		2602: begin l_1 = -12;
				 l_2 = -12; end
		1494: begin l_1 = +13;
				 l_2 = +13; end
		1855: begin l_1 = -13;
				 l_2 = -13; end
		2988: begin l_1 = +14;
				 l_2 = +14; end
		361: begin l_1 = -14;
				 l_2 = -14; end
		2627: begin l_1 = +15;
				 l_2 = +15; end
		722: begin l_1 = -15;
				 l_2 = -15; end
		1905: begin l_1 = +16;
				 l_2 = +16; end
		1444: begin l_1 = -16;
				 l_2 = -16; end
		461: begin l_1 = +17;
				 l_2 = +17; end
		2888: begin l_1 = -17;
				 l_2 = -17; end
		922: begin l_1 = +18;
				 l_2 = +18; end
		2427: begin l_1 = -18;
				 l_2 = -18; end
		1844: begin l_1 = +19;
				 l_2 = +19; end
		1505: begin l_1 = -19;
				 l_2 = -19; end
		339: begin l_1 = +20;
				 l_2 = +20; end
		3010: begin l_1 = -20;
				 l_2 = -20; end
		678: begin l_1 = +21;
				 l_2 = +21; end
		2671: begin l_1 = -21;
				 l_2 = -21; end
		1356: begin l_1 = +22;
				 l_2 = +22; end
		1993: begin l_1 = -22;
				 l_2 = -22; end
		2712: begin l_1 = +23;
				 l_2 = +23; end
		637: begin l_1 = -23;
				 l_2 = -23; end
		3: begin l_1 = -1;
				 l_2 = +3; end
		3346: begin l_1 = -1;
				 l_2 = -2; end
		5: begin l_1 = +1;
				 l_2 = +3; end
		3344: begin l_1 = -1;
				 l_2 = -3; end
		9: begin l_1 = +1;
				 l_2 = +4; end
		3342: begin l_1 = +1;
				 l_2 = -4; end
		7: begin l_1 = -1;
				 l_2 = +4; end
		3340: begin l_1 = -1;
				 l_2 = -4; end
		17: begin l_1 = +1;
				 l_2 = +5; end
		3334: begin l_1 = +1;
				 l_2 = -5; end
		15: begin l_1 = -1;
				 l_2 = +5; end
		3332: begin l_1 = -1;
				 l_2 = -5; end
		33: begin l_1 = +1;
				 l_2 = +6; end
		3318: begin l_1 = +1;
				 l_2 = -6; end
		31: begin l_1 = -1;
				 l_2 = +6; end
		3316: begin l_1 = -1;
				 l_2 = -6; end
		65: begin l_1 = +1;
				 l_2 = +7; end
		3286: begin l_1 = +1;
				 l_2 = -7; end
		63: begin l_1 = -1;
				 l_2 = +7; end
		3284: begin l_1 = -1;
				 l_2 = -7; end
		129: begin l_1 = +1;
				 l_2 = +8; end
		3222: begin l_1 = +1;
				 l_2 = -8; end
		127: begin l_1 = -1;
				 l_2 = +8; end
		3220: begin l_1 = -1;
				 l_2 = -8; end
		257: begin l_1 = +1;
				 l_2 = +9; end
		3094: begin l_1 = +1;
				 l_2 = -9; end
		255: begin l_1 = -1;
				 l_2 = +9; end
		3092: begin l_1 = -1;
				 l_2 = -9; end
		513: begin l_1 = +1;
				 l_2 = +10; end
		2838: begin l_1 = +1;
				 l_2 = -10; end
		511: begin l_1 = -1;
				 l_2 = +10; end
		2836: begin l_1 = -1;
				 l_2 = -10; end
		1025: begin l_1 = +1;
				 l_2 = +11; end
		2326: begin l_1 = +1;
				 l_2 = -11; end
		1023: begin l_1 = -1;
				 l_2 = +11; end
		2324: begin l_1 = -1;
				 l_2 = -11; end
		2049: begin l_1 = +1;
				 l_2 = +12; end
		1302: begin l_1 = +1;
				 l_2 = -12; end
		2047: begin l_1 = -1;
				 l_2 = +12; end
		1300: begin l_1 = -1;
				 l_2 = -12; end
		748: begin l_1 = +1;
				 l_2 = +13; end
		2603: begin l_1 = +1;
				 l_2 = -13; end
		746: begin l_1 = -1;
				 l_2 = +13; end
		2601: begin l_1 = -1;
				 l_2 = -13; end
		1495: begin l_1 = +1;
				 l_2 = +14; end
		1856: begin l_1 = +1;
				 l_2 = -14; end
		1493: begin l_1 = -1;
				 l_2 = +14; end
		1854: begin l_1 = -1;
				 l_2 = -14; end
		2989: begin l_1 = +1;
				 l_2 = +15; end
		362: begin l_1 = +1;
				 l_2 = -15; end
		2987: begin l_1 = -1;
				 l_2 = +15; end
		360: begin l_1 = -1;
				 l_2 = -15; end
		2628: begin l_1 = +1;
				 l_2 = +16; end
		723: begin l_1 = +1;
				 l_2 = -16; end
		2626: begin l_1 = -1;
				 l_2 = +16; end
		721: begin l_1 = -1;
				 l_2 = -16; end
		1906: begin l_1 = +1;
				 l_2 = +17; end
		1445: begin l_1 = +1;
				 l_2 = -17; end
		1904: begin l_1 = -1;
				 l_2 = +17; end
		1443: begin l_1 = -1;
				 l_2 = -17; end
		462: begin l_1 = +1;
				 l_2 = +18; end
		2889: begin l_1 = +1;
				 l_2 = -18; end
		460: begin l_1 = -1;
				 l_2 = +18; end
		2887: begin l_1 = -1;
				 l_2 = -18; end
		923: begin l_1 = +1;
				 l_2 = +19; end
		2428: begin l_1 = +1;
				 l_2 = -19; end
		921: begin l_1 = -1;
				 l_2 = +19; end
		2426: begin l_1 = -1;
				 l_2 = -19; end
		1845: begin l_1 = +1;
				 l_2 = +20; end
		1506: begin l_1 = +1;
				 l_2 = -20; end
		1843: begin l_1 = -1;
				 l_2 = +20; end
		1504: begin l_1 = -1;
				 l_2 = -20; end
		340: begin l_1 = +1;
				 l_2 = +21; end
		3011: begin l_1 = +1;
				 l_2 = -21; end
		338: begin l_1 = -1;
				 l_2 = +21; end
		3009: begin l_1 = -1;
				 l_2 = -21; end
		679: begin l_1 = +1;
				 l_2 = +22; end
		2672: begin l_1 = +1;
				 l_2 = -22; end
		677: begin l_1 = -1;
				 l_2 = +22; end
		2670: begin l_1 = -1;
				 l_2 = -22; end
		1357: begin l_1 = +1;
				 l_2 = +23; end
		1994: begin l_1 = +1;
				 l_2 = -23; end
		1355: begin l_1 = -1;
				 l_2 = +23; end
		1992: begin l_1 = -1;
				 l_2 = -23; end
		2713: begin l_1 = +1;
				 l_2 = +24; end
		638: begin l_1 = +1;
				 l_2 = -24; end
		2711: begin l_1 = -1;
				 l_2 = +24; end
		636: begin l_1 = -1;
				 l_2 = -24; end
		6: begin l_1 = -2;
				 l_2 = +4; end
		3343: begin l_1 = -2;
				 l_2 = -3; end
		10: begin l_1 = +2;
				 l_2 = +4; end
		3339: begin l_1 = -2;
				 l_2 = -4; end
		18: begin l_1 = +2;
				 l_2 = +5; end
		3335: begin l_1 = +2;
				 l_2 = -5; end
		14: begin l_1 = -2;
				 l_2 = +5; end
		3331: begin l_1 = -2;
				 l_2 = -5; end
		34: begin l_1 = +2;
				 l_2 = +6; end
		3319: begin l_1 = +2;
				 l_2 = -6; end
		30: begin l_1 = -2;
				 l_2 = +6; end
		3315: begin l_1 = -2;
				 l_2 = -6; end
		66: begin l_1 = +2;
				 l_2 = +7; end
		3287: begin l_1 = +2;
				 l_2 = -7; end
		62: begin l_1 = -2;
				 l_2 = +7; end
		3283: begin l_1 = -2;
				 l_2 = -7; end
		130: begin l_1 = +2;
				 l_2 = +8; end
		3223: begin l_1 = +2;
				 l_2 = -8; end
		126: begin l_1 = -2;
				 l_2 = +8; end
		3219: begin l_1 = -2;
				 l_2 = -8; end
		258: begin l_1 = +2;
				 l_2 = +9; end
		3095: begin l_1 = +2;
				 l_2 = -9; end
		254: begin l_1 = -2;
				 l_2 = +9; end
		3091: begin l_1 = -2;
				 l_2 = -9; end
		514: begin l_1 = +2;
				 l_2 = +10; end
		2839: begin l_1 = +2;
				 l_2 = -10; end
		510: begin l_1 = -2;
				 l_2 = +10; end
		2835: begin l_1 = -2;
				 l_2 = -10; end
		1026: begin l_1 = +2;
				 l_2 = +11; end
		2327: begin l_1 = +2;
				 l_2 = -11; end
		1022: begin l_1 = -2;
				 l_2 = +11; end
		2323: begin l_1 = -2;
				 l_2 = -11; end
		2050: begin l_1 = +2;
				 l_2 = +12; end
		1303: begin l_1 = +2;
				 l_2 = -12; end
		2046: begin l_1 = -2;
				 l_2 = +12; end
		1299: begin l_1 = -2;
				 l_2 = -12; end
		749: begin l_1 = +2;
				 l_2 = +13; end
		2604: begin l_1 = +2;
				 l_2 = -13; end
		745: begin l_1 = -2;
				 l_2 = +13; end
		2600: begin l_1 = -2;
				 l_2 = -13; end
		1496: begin l_1 = +2;
				 l_2 = +14; end
		1857: begin l_1 = +2;
				 l_2 = -14; end
		1492: begin l_1 = -2;
				 l_2 = +14; end
		1853: begin l_1 = -2;
				 l_2 = -14; end
		2990: begin l_1 = +2;
				 l_2 = +15; end
		363: begin l_1 = +2;
				 l_2 = -15; end
		2986: begin l_1 = -2;
				 l_2 = +15; end
		359: begin l_1 = -2;
				 l_2 = -15; end
		2629: begin l_1 = +2;
				 l_2 = +16; end
		724: begin l_1 = +2;
				 l_2 = -16; end
		2625: begin l_1 = -2;
				 l_2 = +16; end
		720: begin l_1 = -2;
				 l_2 = -16; end
		1907: begin l_1 = +2;
				 l_2 = +17; end
		1446: begin l_1 = +2;
				 l_2 = -17; end
		1903: begin l_1 = -2;
				 l_2 = +17; end
		1442: begin l_1 = -2;
				 l_2 = -17; end
		463: begin l_1 = +2;
				 l_2 = +18; end
		2890: begin l_1 = +2;
				 l_2 = -18; end
		459: begin l_1 = -2;
				 l_2 = +18; end
		2886: begin l_1 = -2;
				 l_2 = -18; end
		924: begin l_1 = +2;
				 l_2 = +19; end
		2429: begin l_1 = +2;
				 l_2 = -19; end
		920: begin l_1 = -2;
				 l_2 = +19; end
		2425: begin l_1 = -2;
				 l_2 = -19; end
		1846: begin l_1 = +2;
				 l_2 = +20; end
		1507: begin l_1 = +2;
				 l_2 = -20; end
		1842: begin l_1 = -2;
				 l_2 = +20; end
		1503: begin l_1 = -2;
				 l_2 = -20; end
		341: begin l_1 = +2;
				 l_2 = +21; end
		3012: begin l_1 = +2;
				 l_2 = -21; end
		337: begin l_1 = -2;
				 l_2 = +21; end
		3008: begin l_1 = -2;
				 l_2 = -21; end
		680: begin l_1 = +2;
				 l_2 = +22; end
		2673: begin l_1 = +2;
				 l_2 = -22; end
		676: begin l_1 = -2;
				 l_2 = +22; end
		2669: begin l_1 = -2;
				 l_2 = -22; end
		1358: begin l_1 = +2;
				 l_2 = +23; end
		1995: begin l_1 = +2;
				 l_2 = -23; end
		1354: begin l_1 = -2;
				 l_2 = +23; end
		1991: begin l_1 = -2;
				 l_2 = -23; end
		2714: begin l_1 = +2;
				 l_2 = +24; end
		639: begin l_1 = +2;
				 l_2 = -24; end
		2710: begin l_1 = -2;
				 l_2 = +24; end
		635: begin l_1 = -2;
				 l_2 = -24; end
		12: begin l_1 = -3;
				 l_2 = +5; end
		3337: begin l_1 = -3;
				 l_2 = -4; end
		20: begin l_1 = +3;
				 l_2 = +5; end
		3329: begin l_1 = -3;
				 l_2 = -5; end
		36: begin l_1 = +3;
				 l_2 = +6; end
		3321: begin l_1 = +3;
				 l_2 = -6; end
		28: begin l_1 = -3;
				 l_2 = +6; end
		3313: begin l_1 = -3;
				 l_2 = -6; end
		68: begin l_1 = +3;
				 l_2 = +7; end
		3289: begin l_1 = +3;
				 l_2 = -7; end
		60: begin l_1 = -3;
				 l_2 = +7; end
		3281: begin l_1 = -3;
				 l_2 = -7; end
		132: begin l_1 = +3;
				 l_2 = +8; end
		3225: begin l_1 = +3;
				 l_2 = -8; end
		124: begin l_1 = -3;
				 l_2 = +8; end
		3217: begin l_1 = -3;
				 l_2 = -8; end
		260: begin l_1 = +3;
				 l_2 = +9; end
		3097: begin l_1 = +3;
				 l_2 = -9; end
		252: begin l_1 = -3;
				 l_2 = +9; end
		3089: begin l_1 = -3;
				 l_2 = -9; end
		516: begin l_1 = +3;
				 l_2 = +10; end
		2841: begin l_1 = +3;
				 l_2 = -10; end
		508: begin l_1 = -3;
				 l_2 = +10; end
		2833: begin l_1 = -3;
				 l_2 = -10; end
		1028: begin l_1 = +3;
				 l_2 = +11; end
		2329: begin l_1 = +3;
				 l_2 = -11; end
		1020: begin l_1 = -3;
				 l_2 = +11; end
		2321: begin l_1 = -3;
				 l_2 = -11; end
		2052: begin l_1 = +3;
				 l_2 = +12; end
		1305: begin l_1 = +3;
				 l_2 = -12; end
		2044: begin l_1 = -3;
				 l_2 = +12; end
		1297: begin l_1 = -3;
				 l_2 = -12; end
		751: begin l_1 = +3;
				 l_2 = +13; end
		2606: begin l_1 = +3;
				 l_2 = -13; end
		743: begin l_1 = -3;
				 l_2 = +13; end
		2598: begin l_1 = -3;
				 l_2 = -13; end
		1498: begin l_1 = +3;
				 l_2 = +14; end
		1859: begin l_1 = +3;
				 l_2 = -14; end
		1490: begin l_1 = -3;
				 l_2 = +14; end
		1851: begin l_1 = -3;
				 l_2 = -14; end
		2992: begin l_1 = +3;
				 l_2 = +15; end
		365: begin l_1 = +3;
				 l_2 = -15; end
		2984: begin l_1 = -3;
				 l_2 = +15; end
		357: begin l_1 = -3;
				 l_2 = -15; end
		2631: begin l_1 = +3;
				 l_2 = +16; end
		726: begin l_1 = +3;
				 l_2 = -16; end
		2623: begin l_1 = -3;
				 l_2 = +16; end
		718: begin l_1 = -3;
				 l_2 = -16; end
		1909: begin l_1 = +3;
				 l_2 = +17; end
		1448: begin l_1 = +3;
				 l_2 = -17; end
		1901: begin l_1 = -3;
				 l_2 = +17; end
		1440: begin l_1 = -3;
				 l_2 = -17; end
		465: begin l_1 = +3;
				 l_2 = +18; end
		2892: begin l_1 = +3;
				 l_2 = -18; end
		457: begin l_1 = -3;
				 l_2 = +18; end
		2884: begin l_1 = -3;
				 l_2 = -18; end
		926: begin l_1 = +3;
				 l_2 = +19; end
		2431: begin l_1 = +3;
				 l_2 = -19; end
		918: begin l_1 = -3;
				 l_2 = +19; end
		2423: begin l_1 = -3;
				 l_2 = -19; end
		1848: begin l_1 = +3;
				 l_2 = +20; end
		1509: begin l_1 = +3;
				 l_2 = -20; end
		1840: begin l_1 = -3;
				 l_2 = +20; end
		1501: begin l_1 = -3;
				 l_2 = -20; end
		343: begin l_1 = +3;
				 l_2 = +21; end
		3014: begin l_1 = +3;
				 l_2 = -21; end
		335: begin l_1 = -3;
				 l_2 = +21; end
		3006: begin l_1 = -3;
				 l_2 = -21; end
		682: begin l_1 = +3;
				 l_2 = +22; end
		2675: begin l_1 = +3;
				 l_2 = -22; end
		674: begin l_1 = -3;
				 l_2 = +22; end
		2667: begin l_1 = -3;
				 l_2 = -22; end
		1360: begin l_1 = +3;
				 l_2 = +23; end
		1997: begin l_1 = +3;
				 l_2 = -23; end
		1352: begin l_1 = -3;
				 l_2 = +23; end
		1989: begin l_1 = -3;
				 l_2 = -23; end
		2716: begin l_1 = +3;
				 l_2 = +24; end
		641: begin l_1 = +3;
				 l_2 = -24; end
		2708: begin l_1 = -3;
				 l_2 = +24; end
		633: begin l_1 = -3;
				 l_2 = -24; end
		24: begin l_1 = -4;
				 l_2 = +6; end
		3325: begin l_1 = -4;
				 l_2 = -5; end
		40: begin l_1 = +4;
				 l_2 = +6; end
		3309: begin l_1 = -4;
				 l_2 = -6; end
		72: begin l_1 = +4;
				 l_2 = +7; end
		3293: begin l_1 = +4;
				 l_2 = -7; end
		56: begin l_1 = -4;
				 l_2 = +7; end
		3277: begin l_1 = -4;
				 l_2 = -7; end
		136: begin l_1 = +4;
				 l_2 = +8; end
		3229: begin l_1 = +4;
				 l_2 = -8; end
		120: begin l_1 = -4;
				 l_2 = +8; end
		3213: begin l_1 = -4;
				 l_2 = -8; end
		264: begin l_1 = +4;
				 l_2 = +9; end
		3101: begin l_1 = +4;
				 l_2 = -9; end
		248: begin l_1 = -4;
				 l_2 = +9; end
		3085: begin l_1 = -4;
				 l_2 = -9; end
		520: begin l_1 = +4;
				 l_2 = +10; end
		2845: begin l_1 = +4;
				 l_2 = -10; end
		504: begin l_1 = -4;
				 l_2 = +10; end
		2829: begin l_1 = -4;
				 l_2 = -10; end
		1032: begin l_1 = +4;
				 l_2 = +11; end
		2333: begin l_1 = +4;
				 l_2 = -11; end
		1016: begin l_1 = -4;
				 l_2 = +11; end
		2317: begin l_1 = -4;
				 l_2 = -11; end
		2056: begin l_1 = +4;
				 l_2 = +12; end
		1309: begin l_1 = +4;
				 l_2 = -12; end
		2040: begin l_1 = -4;
				 l_2 = +12; end
		1293: begin l_1 = -4;
				 l_2 = -12; end
		755: begin l_1 = +4;
				 l_2 = +13; end
		2610: begin l_1 = +4;
				 l_2 = -13; end
		739: begin l_1 = -4;
				 l_2 = +13; end
		2594: begin l_1 = -4;
				 l_2 = -13; end
		1502: begin l_1 = +4;
				 l_2 = +14; end
		1863: begin l_1 = +4;
				 l_2 = -14; end
		1486: begin l_1 = -4;
				 l_2 = +14; end
		1847: begin l_1 = -4;
				 l_2 = -14; end
		2996: begin l_1 = +4;
				 l_2 = +15; end
		369: begin l_1 = +4;
				 l_2 = -15; end
		2980: begin l_1 = -4;
				 l_2 = +15; end
		353: begin l_1 = -4;
				 l_2 = -15; end
		2635: begin l_1 = +4;
				 l_2 = +16; end
		730: begin l_1 = +4;
				 l_2 = -16; end
		2619: begin l_1 = -4;
				 l_2 = +16; end
		714: begin l_1 = -4;
				 l_2 = -16; end
		1913: begin l_1 = +4;
				 l_2 = +17; end
		1452: begin l_1 = +4;
				 l_2 = -17; end
		1897: begin l_1 = -4;
				 l_2 = +17; end
		1436: begin l_1 = -4;
				 l_2 = -17; end
		469: begin l_1 = +4;
				 l_2 = +18; end
		2896: begin l_1 = +4;
				 l_2 = -18; end
		453: begin l_1 = -4;
				 l_2 = +18; end
		2880: begin l_1 = -4;
				 l_2 = -18; end
		930: begin l_1 = +4;
				 l_2 = +19; end
		2435: begin l_1 = +4;
				 l_2 = -19; end
		914: begin l_1 = -4;
				 l_2 = +19; end
		2419: begin l_1 = -4;
				 l_2 = -19; end
		1852: begin l_1 = +4;
				 l_2 = +20; end
		1513: begin l_1 = +4;
				 l_2 = -20; end
		1836: begin l_1 = -4;
				 l_2 = +20; end
		1497: begin l_1 = -4;
				 l_2 = -20; end
		347: begin l_1 = +4;
				 l_2 = +21; end
		3018: begin l_1 = +4;
				 l_2 = -21; end
		331: begin l_1 = -4;
				 l_2 = +21; end
		3002: begin l_1 = -4;
				 l_2 = -21; end
		686: begin l_1 = +4;
				 l_2 = +22; end
		2679: begin l_1 = +4;
				 l_2 = -22; end
		670: begin l_1 = -4;
				 l_2 = +22; end
		2663: begin l_1 = -4;
				 l_2 = -22; end
		1364: begin l_1 = +4;
				 l_2 = +23; end
		2001: begin l_1 = +4;
				 l_2 = -23; end
		1348: begin l_1 = -4;
				 l_2 = +23; end
		1985: begin l_1 = -4;
				 l_2 = -23; end
		2720: begin l_1 = +4;
				 l_2 = +24; end
		645: begin l_1 = +4;
				 l_2 = -24; end
		2704: begin l_1 = -4;
				 l_2 = +24; end
		629: begin l_1 = -4;
				 l_2 = -24; end
		48: begin l_1 = -5;
				 l_2 = +7; end
		3301: begin l_1 = -5;
				 l_2 = -6; end
		80: begin l_1 = +5;
				 l_2 = +7; end
		3269: begin l_1 = -5;
				 l_2 = -7; end
		144: begin l_1 = +5;
				 l_2 = +8; end
		3237: begin l_1 = +5;
				 l_2 = -8; end
		112: begin l_1 = -5;
				 l_2 = +8; end
		3205: begin l_1 = -5;
				 l_2 = -8; end
		272: begin l_1 = +5;
				 l_2 = +9; end
		3109: begin l_1 = +5;
				 l_2 = -9; end
		240: begin l_1 = -5;
				 l_2 = +9; end
		3077: begin l_1 = -5;
				 l_2 = -9; end
		528: begin l_1 = +5;
				 l_2 = +10; end
		2853: begin l_1 = +5;
				 l_2 = -10; end
		496: begin l_1 = -5;
				 l_2 = +10; end
		2821: begin l_1 = -5;
				 l_2 = -10; end
		1040: begin l_1 = +5;
				 l_2 = +11; end
		2341: begin l_1 = +5;
				 l_2 = -11; end
		1008: begin l_1 = -5;
				 l_2 = +11; end
		2309: begin l_1 = -5;
				 l_2 = -11; end
		2064: begin l_1 = +5;
				 l_2 = +12; end
		1317: begin l_1 = +5;
				 l_2 = -12; end
		2032: begin l_1 = -5;
				 l_2 = +12; end
		1285: begin l_1 = -5;
				 l_2 = -12; end
		763: begin l_1 = +5;
				 l_2 = +13; end
		2618: begin l_1 = +5;
				 l_2 = -13; end
		731: begin l_1 = -5;
				 l_2 = +13; end
		2586: begin l_1 = -5;
				 l_2 = -13; end
		1510: begin l_1 = +5;
				 l_2 = +14; end
		1871: begin l_1 = +5;
				 l_2 = -14; end
		1478: begin l_1 = -5;
				 l_2 = +14; end
		1839: begin l_1 = -5;
				 l_2 = -14; end
		3004: begin l_1 = +5;
				 l_2 = +15; end
		377: begin l_1 = +5;
				 l_2 = -15; end
		2972: begin l_1 = -5;
				 l_2 = +15; end
		345: begin l_1 = -5;
				 l_2 = -15; end
		2643: begin l_1 = +5;
				 l_2 = +16; end
		738: begin l_1 = +5;
				 l_2 = -16; end
		2611: begin l_1 = -5;
				 l_2 = +16; end
		706: begin l_1 = -5;
				 l_2 = -16; end
		1921: begin l_1 = +5;
				 l_2 = +17; end
		1460: begin l_1 = +5;
				 l_2 = -17; end
		1889: begin l_1 = -5;
				 l_2 = +17; end
		1428: begin l_1 = -5;
				 l_2 = -17; end
		477: begin l_1 = +5;
				 l_2 = +18; end
		2904: begin l_1 = +5;
				 l_2 = -18; end
		445: begin l_1 = -5;
				 l_2 = +18; end
		2872: begin l_1 = -5;
				 l_2 = -18; end
		938: begin l_1 = +5;
				 l_2 = +19; end
		2443: begin l_1 = +5;
				 l_2 = -19; end
		906: begin l_1 = -5;
				 l_2 = +19; end
		2411: begin l_1 = -5;
				 l_2 = -19; end
		1860: begin l_1 = +5;
				 l_2 = +20; end
		1521: begin l_1 = +5;
				 l_2 = -20; end
		1828: begin l_1 = -5;
				 l_2 = +20; end
		1489: begin l_1 = -5;
				 l_2 = -20; end
		355: begin l_1 = +5;
				 l_2 = +21; end
		3026: begin l_1 = +5;
				 l_2 = -21; end
		323: begin l_1 = -5;
				 l_2 = +21; end
		2994: begin l_1 = -5;
				 l_2 = -21; end
		694: begin l_1 = +5;
				 l_2 = +22; end
		2687: begin l_1 = +5;
				 l_2 = -22; end
		662: begin l_1 = -5;
				 l_2 = +22; end
		2655: begin l_1 = -5;
				 l_2 = -22; end
		1372: begin l_1 = +5;
				 l_2 = +23; end
		2009: begin l_1 = +5;
				 l_2 = -23; end
		1340: begin l_1 = -5;
				 l_2 = +23; end
		1977: begin l_1 = -5;
				 l_2 = -23; end
		2728: begin l_1 = +5;
				 l_2 = +24; end
		653: begin l_1 = +5;
				 l_2 = -24; end
		2696: begin l_1 = -5;
				 l_2 = +24; end
		621: begin l_1 = -5;
				 l_2 = -24; end
		96: begin l_1 = -6;
				 l_2 = +8; end
		3253: begin l_1 = -6;
				 l_2 = -7; end
		160: begin l_1 = +6;
				 l_2 = +8; end
		3189: begin l_1 = -6;
				 l_2 = -8; end
		288: begin l_1 = +6;
				 l_2 = +9; end
		3125: begin l_1 = +6;
				 l_2 = -9; end
		224: begin l_1 = -6;
				 l_2 = +9; end
		3061: begin l_1 = -6;
				 l_2 = -9; end
		544: begin l_1 = +6;
				 l_2 = +10; end
		2869: begin l_1 = +6;
				 l_2 = -10; end
		480: begin l_1 = -6;
				 l_2 = +10; end
		2805: begin l_1 = -6;
				 l_2 = -10; end
		1056: begin l_1 = +6;
				 l_2 = +11; end
		2357: begin l_1 = +6;
				 l_2 = -11; end
		992: begin l_1 = -6;
				 l_2 = +11; end
		2293: begin l_1 = -6;
				 l_2 = -11; end
		2080: begin l_1 = +6;
				 l_2 = +12; end
		1333: begin l_1 = +6;
				 l_2 = -12; end
		2016: begin l_1 = -6;
				 l_2 = +12; end
		1269: begin l_1 = -6;
				 l_2 = -12; end
		779: begin l_1 = +6;
				 l_2 = +13; end
		2634: begin l_1 = +6;
				 l_2 = -13; end
		715: begin l_1 = -6;
				 l_2 = +13; end
		2570: begin l_1 = -6;
				 l_2 = -13; end
		1526: begin l_1 = +6;
				 l_2 = +14; end
		1887: begin l_1 = +6;
				 l_2 = -14; end
		1462: begin l_1 = -6;
				 l_2 = +14; end
		1823: begin l_1 = -6;
				 l_2 = -14; end
		3020: begin l_1 = +6;
				 l_2 = +15; end
		393: begin l_1 = +6;
				 l_2 = -15; end
		2956: begin l_1 = -6;
				 l_2 = +15; end
		329: begin l_1 = -6;
				 l_2 = -15; end
		2659: begin l_1 = +6;
				 l_2 = +16; end
		754: begin l_1 = +6;
				 l_2 = -16; end
		2595: begin l_1 = -6;
				 l_2 = +16; end
		690: begin l_1 = -6;
				 l_2 = -16; end
		1937: begin l_1 = +6;
				 l_2 = +17; end
		1476: begin l_1 = +6;
				 l_2 = -17; end
		1873: begin l_1 = -6;
				 l_2 = +17; end
		1412: begin l_1 = -6;
				 l_2 = -17; end
		493: begin l_1 = +6;
				 l_2 = +18; end
		2920: begin l_1 = +6;
				 l_2 = -18; end
		429: begin l_1 = -6;
				 l_2 = +18; end
		2856: begin l_1 = -6;
				 l_2 = -18; end
		954: begin l_1 = +6;
				 l_2 = +19; end
		2459: begin l_1 = +6;
				 l_2 = -19; end
		890: begin l_1 = -6;
				 l_2 = +19; end
		2395: begin l_1 = -6;
				 l_2 = -19; end
		1876: begin l_1 = +6;
				 l_2 = +20; end
		1537: begin l_1 = +6;
				 l_2 = -20; end
		1812: begin l_1 = -6;
				 l_2 = +20; end
		1473: begin l_1 = -6;
				 l_2 = -20; end
		371: begin l_1 = +6;
				 l_2 = +21; end
		3042: begin l_1 = +6;
				 l_2 = -21; end
		307: begin l_1 = -6;
				 l_2 = +21; end
		2978: begin l_1 = -6;
				 l_2 = -21; end
		710: begin l_1 = +6;
				 l_2 = +22; end
		2703: begin l_1 = +6;
				 l_2 = -22; end
		646: begin l_1 = -6;
				 l_2 = +22; end
		2639: begin l_1 = -6;
				 l_2 = -22; end
		1388: begin l_1 = +6;
				 l_2 = +23; end
		2025: begin l_1 = +6;
				 l_2 = -23; end
		1324: begin l_1 = -6;
				 l_2 = +23; end
		1961: begin l_1 = -6;
				 l_2 = -23; end
		2744: begin l_1 = +6;
				 l_2 = +24; end
		669: begin l_1 = +6;
				 l_2 = -24; end
		2680: begin l_1 = -6;
				 l_2 = +24; end
		605: begin l_1 = -6;
				 l_2 = -24; end
		192: begin l_1 = -7;
				 l_2 = +9; end
		3157: begin l_1 = -7;
				 l_2 = -8; end
		320: begin l_1 = +7;
				 l_2 = +9; end
		3029: begin l_1 = -7;
				 l_2 = -9; end
		576: begin l_1 = +7;
				 l_2 = +10; end
		2901: begin l_1 = +7;
				 l_2 = -10; end
		448: begin l_1 = -7;
				 l_2 = +10; end
		2773: begin l_1 = -7;
				 l_2 = -10; end
		1088: begin l_1 = +7;
				 l_2 = +11; end
		2389: begin l_1 = +7;
				 l_2 = -11; end
		960: begin l_1 = -7;
				 l_2 = +11; end
		2261: begin l_1 = -7;
				 l_2 = -11; end
		2112: begin l_1 = +7;
				 l_2 = +12; end
		1365: begin l_1 = +7;
				 l_2 = -12; end
		1984: begin l_1 = -7;
				 l_2 = +12; end
		1237: begin l_1 = -7;
				 l_2 = -12; end
		811: begin l_1 = +7;
				 l_2 = +13; end
		2666: begin l_1 = +7;
				 l_2 = -13; end
		683: begin l_1 = -7;
				 l_2 = +13; end
		2538: begin l_1 = -7;
				 l_2 = -13; end
		1558: begin l_1 = +7;
				 l_2 = +14; end
		1919: begin l_1 = +7;
				 l_2 = -14; end
		1430: begin l_1 = -7;
				 l_2 = +14; end
		1791: begin l_1 = -7;
				 l_2 = -14; end
		3052: begin l_1 = +7;
				 l_2 = +15; end
		425: begin l_1 = +7;
				 l_2 = -15; end
		2924: begin l_1 = -7;
				 l_2 = +15; end
		297: begin l_1 = -7;
				 l_2 = -15; end
		2691: begin l_1 = +7;
				 l_2 = +16; end
		786: begin l_1 = +7;
				 l_2 = -16; end
		2563: begin l_1 = -7;
				 l_2 = +16; end
		658: begin l_1 = -7;
				 l_2 = -16; end
		1969: begin l_1 = +7;
				 l_2 = +17; end
		1508: begin l_1 = +7;
				 l_2 = -17; end
		1841: begin l_1 = -7;
				 l_2 = +17; end
		1380: begin l_1 = -7;
				 l_2 = -17; end
		525: begin l_1 = +7;
				 l_2 = +18; end
		2952: begin l_1 = +7;
				 l_2 = -18; end
		397: begin l_1 = -7;
				 l_2 = +18; end
		2824: begin l_1 = -7;
				 l_2 = -18; end
		986: begin l_1 = +7;
				 l_2 = +19; end
		2491: begin l_1 = +7;
				 l_2 = -19; end
		858: begin l_1 = -7;
				 l_2 = +19; end
		2363: begin l_1 = -7;
				 l_2 = -19; end
		1908: begin l_1 = +7;
				 l_2 = +20; end
		1569: begin l_1 = +7;
				 l_2 = -20; end
		1780: begin l_1 = -7;
				 l_2 = +20; end
		1441: begin l_1 = -7;
				 l_2 = -20; end
		403: begin l_1 = +7;
				 l_2 = +21; end
		3074: begin l_1 = +7;
				 l_2 = -21; end
		275: begin l_1 = -7;
				 l_2 = +21; end
		2946: begin l_1 = -7;
				 l_2 = -21; end
		742: begin l_1 = +7;
				 l_2 = +22; end
		2735: begin l_1 = +7;
				 l_2 = -22; end
		614: begin l_1 = -7;
				 l_2 = +22; end
		2607: begin l_1 = -7;
				 l_2 = -22; end
		1420: begin l_1 = +7;
				 l_2 = +23; end
		2057: begin l_1 = +7;
				 l_2 = -23; end
		1292: begin l_1 = -7;
				 l_2 = +23; end
		1929: begin l_1 = -7;
				 l_2 = -23; end
		2776: begin l_1 = +7;
				 l_2 = +24; end
		701: begin l_1 = +7;
				 l_2 = -24; end
		2648: begin l_1 = -7;
				 l_2 = +24; end
		573: begin l_1 = -7;
				 l_2 = -24; end
		384: begin l_1 = -8;
				 l_2 = +10; end
		2965: begin l_1 = -8;
				 l_2 = -9; end
		640: begin l_1 = +8;
				 l_2 = +10; end
		2709: begin l_1 = -8;
				 l_2 = -10; end
		1152: begin l_1 = +8;
				 l_2 = +11; end
		2453: begin l_1 = +8;
				 l_2 = -11; end
		896: begin l_1 = -8;
				 l_2 = +11; end
		2197: begin l_1 = -8;
				 l_2 = -11; end
		2176: begin l_1 = +8;
				 l_2 = +12; end
		1429: begin l_1 = +8;
				 l_2 = -12; end
		1920: begin l_1 = -8;
				 l_2 = +12; end
		1173: begin l_1 = -8;
				 l_2 = -12; end
		875: begin l_1 = +8;
				 l_2 = +13; end
		2730: begin l_1 = +8;
				 l_2 = -13; end
		619: begin l_1 = -8;
				 l_2 = +13; end
		2474: begin l_1 = -8;
				 l_2 = -13; end
		1622: begin l_1 = +8;
				 l_2 = +14; end
		1983: begin l_1 = +8;
				 l_2 = -14; end
		1366: begin l_1 = -8;
				 l_2 = +14; end
		1727: begin l_1 = -8;
				 l_2 = -14; end
		3116: begin l_1 = +8;
				 l_2 = +15; end
		489: begin l_1 = +8;
				 l_2 = -15; end
		2860: begin l_1 = -8;
				 l_2 = +15; end
		233: begin l_1 = -8;
				 l_2 = -15; end
		2755: begin l_1 = +8;
				 l_2 = +16; end
		850: begin l_1 = +8;
				 l_2 = -16; end
		2499: begin l_1 = -8;
				 l_2 = +16; end
		594: begin l_1 = -8;
				 l_2 = -16; end
		2033: begin l_1 = +8;
				 l_2 = +17; end
		1572: begin l_1 = +8;
				 l_2 = -17; end
		1777: begin l_1 = -8;
				 l_2 = +17; end
		1316: begin l_1 = -8;
				 l_2 = -17; end
		589: begin l_1 = +8;
				 l_2 = +18; end
		3016: begin l_1 = +8;
				 l_2 = -18; end
		333: begin l_1 = -8;
				 l_2 = +18; end
		2760: begin l_1 = -8;
				 l_2 = -18; end
		1050: begin l_1 = +8;
				 l_2 = +19; end
		2555: begin l_1 = +8;
				 l_2 = -19; end
		794: begin l_1 = -8;
				 l_2 = +19; end
		2299: begin l_1 = -8;
				 l_2 = -19; end
		1972: begin l_1 = +8;
				 l_2 = +20; end
		1633: begin l_1 = +8;
				 l_2 = -20; end
		1716: begin l_1 = -8;
				 l_2 = +20; end
		1377: begin l_1 = -8;
				 l_2 = -20; end
		467: begin l_1 = +8;
				 l_2 = +21; end
		3138: begin l_1 = +8;
				 l_2 = -21; end
		211: begin l_1 = -8;
				 l_2 = +21; end
		2882: begin l_1 = -8;
				 l_2 = -21; end
		806: begin l_1 = +8;
				 l_2 = +22; end
		2799: begin l_1 = +8;
				 l_2 = -22; end
		550: begin l_1 = -8;
				 l_2 = +22; end
		2543: begin l_1 = -8;
				 l_2 = -22; end
		1484: begin l_1 = +8;
				 l_2 = +23; end
		2121: begin l_1 = +8;
				 l_2 = -23; end
		1228: begin l_1 = -8;
				 l_2 = +23; end
		1865: begin l_1 = -8;
				 l_2 = -23; end
		2840: begin l_1 = +8;
				 l_2 = +24; end
		765: begin l_1 = +8;
				 l_2 = -24; end
		2584: begin l_1 = -8;
				 l_2 = +24; end
		509: begin l_1 = -8;
				 l_2 = -24; end
		768: begin l_1 = -9;
				 l_2 = +11; end
		2581: begin l_1 = -9;
				 l_2 = -10; end
		1280: begin l_1 = +9;
				 l_2 = +11; end
		2069: begin l_1 = -9;
				 l_2 = -11; end
		2304: begin l_1 = +9;
				 l_2 = +12; end
		1557: begin l_1 = +9;
				 l_2 = -12; end
		1792: begin l_1 = -9;
				 l_2 = +12; end
		1045: begin l_1 = -9;
				 l_2 = -12; end
		1003: begin l_1 = +9;
				 l_2 = +13; end
		2858: begin l_1 = +9;
				 l_2 = -13; end
		491: begin l_1 = -9;
				 l_2 = +13; end
		2346: begin l_1 = -9;
				 l_2 = -13; end
		1750: begin l_1 = +9;
				 l_2 = +14; end
		2111: begin l_1 = +9;
				 l_2 = -14; end
		1238: begin l_1 = -9;
				 l_2 = +14; end
		1599: begin l_1 = -9;
				 l_2 = -14; end
		3244: begin l_1 = +9;
				 l_2 = +15; end
		617: begin l_1 = +9;
				 l_2 = -15; end
		2732: begin l_1 = -9;
				 l_2 = +15; end
		105: begin l_1 = -9;
				 l_2 = -15; end
		2883: begin l_1 = +9;
				 l_2 = +16; end
		978: begin l_1 = +9;
				 l_2 = -16; end
		2371: begin l_1 = -9;
				 l_2 = +16; end
		466: begin l_1 = -9;
				 l_2 = -16; end
		2161: begin l_1 = +9;
				 l_2 = +17; end
		1700: begin l_1 = +9;
				 l_2 = -17; end
		1649: begin l_1 = -9;
				 l_2 = +17; end
		1188: begin l_1 = -9;
				 l_2 = -17; end
		717: begin l_1 = +9;
				 l_2 = +18; end
		3144: begin l_1 = +9;
				 l_2 = -18; end
		205: begin l_1 = -9;
				 l_2 = +18; end
		2632: begin l_1 = -9;
				 l_2 = -18; end
		1178: begin l_1 = +9;
				 l_2 = +19; end
		2683: begin l_1 = +9;
				 l_2 = -19; end
		666: begin l_1 = -9;
				 l_2 = +19; end
		2171: begin l_1 = -9;
				 l_2 = -19; end
		2100: begin l_1 = +9;
				 l_2 = +20; end
		1761: begin l_1 = +9;
				 l_2 = -20; end
		1588: begin l_1 = -9;
				 l_2 = +20; end
		1249: begin l_1 = -9;
				 l_2 = -20; end
		595: begin l_1 = +9;
				 l_2 = +21; end
		3266: begin l_1 = +9;
				 l_2 = -21; end
		83: begin l_1 = -9;
				 l_2 = +21; end
		2754: begin l_1 = -9;
				 l_2 = -21; end
		934: begin l_1 = +9;
				 l_2 = +22; end
		2927: begin l_1 = +9;
				 l_2 = -22; end
		422: begin l_1 = -9;
				 l_2 = +22; end
		2415: begin l_1 = -9;
				 l_2 = -22; end
		1612: begin l_1 = +9;
				 l_2 = +23; end
		2249: begin l_1 = +9;
				 l_2 = -23; end
		1100: begin l_1 = -9;
				 l_2 = +23; end
		1737: begin l_1 = -9;
				 l_2 = -23; end
		2968: begin l_1 = +9;
				 l_2 = +24; end
		893: begin l_1 = +9;
				 l_2 = -24; end
		2456: begin l_1 = -9;
				 l_2 = +24; end
		381: begin l_1 = -9;
				 l_2 = -24; end
		1536: begin l_1 = -10;
				 l_2 = +12; end
		1813: begin l_1 = -10;
				 l_2 = -11; end
		2560: begin l_1 = +10;
				 l_2 = +12; end
		789: begin l_1 = -10;
				 l_2 = -12; end
		1259: begin l_1 = +10;
				 l_2 = +13; end
		3114: begin l_1 = +10;
				 l_2 = -13; end
		235: begin l_1 = -10;
				 l_2 = +13; end
		2090: begin l_1 = -10;
				 l_2 = -13; end
		2006: begin l_1 = +10;
				 l_2 = +14; end
		2367: begin l_1 = +10;
				 l_2 = -14; end
		982: begin l_1 = -10;
				 l_2 = +14; end
		1343: begin l_1 = -10;
				 l_2 = -14; end
		151: begin l_1 = +10;
				 l_2 = +15; end
		873: begin l_1 = +10;
				 l_2 = -15; end
		2476: begin l_1 = -10;
				 l_2 = +15; end
		3198: begin l_1 = -10;
				 l_2 = -15; end
		3139: begin l_1 = +10;
				 l_2 = +16; end
		1234: begin l_1 = +10;
				 l_2 = -16; end
		2115: begin l_1 = -10;
				 l_2 = +16; end
		210: begin l_1 = -10;
				 l_2 = -16; end
		2417: begin l_1 = +10;
				 l_2 = +17; end
		1956: begin l_1 = +10;
				 l_2 = -17; end
		1393: begin l_1 = -10;
				 l_2 = +17; end
		932: begin l_1 = -10;
				 l_2 = -17; end
		973: begin l_1 = +10;
				 l_2 = +18; end
		51: begin l_1 = +10;
				 l_2 = -18; end
		3298: begin l_1 = -10;
				 l_2 = +18; end
		2376: begin l_1 = -10;
				 l_2 = -18; end
		1434: begin l_1 = +10;
				 l_2 = +19; end
		2939: begin l_1 = +10;
				 l_2 = -19; end
		410: begin l_1 = -10;
				 l_2 = +19; end
		1915: begin l_1 = -10;
				 l_2 = -19; end
		2356: begin l_1 = +10;
				 l_2 = +20; end
		2017: begin l_1 = +10;
				 l_2 = -20; end
		1332: begin l_1 = -10;
				 l_2 = +20; end
		993: begin l_1 = -10;
				 l_2 = -20; end
		851: begin l_1 = +10;
				 l_2 = +21; end
		173: begin l_1 = +10;
				 l_2 = -21; end
		3176: begin l_1 = -10;
				 l_2 = +21; end
		2498: begin l_1 = -10;
				 l_2 = -21; end
		1190: begin l_1 = +10;
				 l_2 = +22; end
		3183: begin l_1 = +10;
				 l_2 = -22; end
		166: begin l_1 = -10;
				 l_2 = +22; end
		2159: begin l_1 = -10;
				 l_2 = -22; end
		1868: begin l_1 = +10;
				 l_2 = +23; end
		2505: begin l_1 = +10;
				 l_2 = -23; end
		844: begin l_1 = -10;
				 l_2 = +23; end
		1481: begin l_1 = -10;
				 l_2 = -23; end
		3224: begin l_1 = +10;
				 l_2 = +24; end
		1149: begin l_1 = +10;
				 l_2 = -24; end
		2200: begin l_1 = -10;
				 l_2 = +24; end
		125: begin l_1 = -10;
				 l_2 = -24; end
		3072: begin l_1 = -11;
				 l_2 = +13; end
		277: begin l_1 = -11;
				 l_2 = -12; end
		1771: begin l_1 = +11;
				 l_2 = +13; end
		1578: begin l_1 = -11;
				 l_2 = -13; end
		2518: begin l_1 = +11;
				 l_2 = +14; end
		2879: begin l_1 = +11;
				 l_2 = -14; end
		470: begin l_1 = -11;
				 l_2 = +14; end
		831: begin l_1 = -11;
				 l_2 = -14; end
		663: begin l_1 = +11;
				 l_2 = +15; end
		1385: begin l_1 = +11;
				 l_2 = -15; end
		1964: begin l_1 = -11;
				 l_2 = +15; end
		2686: begin l_1 = -11;
				 l_2 = -15; end
		302: begin l_1 = +11;
				 l_2 = +16; end
		1746: begin l_1 = +11;
				 l_2 = -16; end
		1603: begin l_1 = -11;
				 l_2 = +16; end
		3047: begin l_1 = -11;
				 l_2 = -16; end
		2929: begin l_1 = +11;
				 l_2 = +17; end
		2468: begin l_1 = +11;
				 l_2 = -17; end
		881: begin l_1 = -11;
				 l_2 = +17; end
		420: begin l_1 = -11;
				 l_2 = -17; end
		1485: begin l_1 = +11;
				 l_2 = +18; end
		563: begin l_1 = +11;
				 l_2 = -18; end
		2786: begin l_1 = -11;
				 l_2 = +18; end
		1864: begin l_1 = -11;
				 l_2 = -18; end
		1946: begin l_1 = +11;
				 l_2 = +19; end
		102: begin l_1 = +11;
				 l_2 = -19; end
		3247: begin l_1 = -11;
				 l_2 = +19; end
		1403: begin l_1 = -11;
				 l_2 = -19; end
		2868: begin l_1 = +11;
				 l_2 = +20; end
		2529: begin l_1 = +11;
				 l_2 = -20; end
		820: begin l_1 = -11;
				 l_2 = +20; end
		481: begin l_1 = -11;
				 l_2 = -20; end
		1363: begin l_1 = +11;
				 l_2 = +21; end
		685: begin l_1 = +11;
				 l_2 = -21; end
		2664: begin l_1 = -11;
				 l_2 = +21; end
		1986: begin l_1 = -11;
				 l_2 = -21; end
		1702: begin l_1 = +11;
				 l_2 = +22; end
		346: begin l_1 = +11;
				 l_2 = -22; end
		3003: begin l_1 = -11;
				 l_2 = +22; end
		1647: begin l_1 = -11;
				 l_2 = -22; end
		2380: begin l_1 = +11;
				 l_2 = +23; end
		3017: begin l_1 = +11;
				 l_2 = -23; end
		332: begin l_1 = -11;
				 l_2 = +23; end
		969: begin l_1 = -11;
				 l_2 = -23; end
		387: begin l_1 = +11;
				 l_2 = +24; end
		1661: begin l_1 = +11;
				 l_2 = -24; end
		1688: begin l_1 = -11;
				 l_2 = +24; end
		2962: begin l_1 = -11;
				 l_2 = -24; end
		2795: begin l_1 = -12;
				 l_2 = +14; end
		554: begin l_1 = -12;
				 l_2 = -13; end
		193: begin l_1 = +12;
				 l_2 = +14; end
		3156: begin l_1 = -12;
				 l_2 = -14; end
		1687: begin l_1 = +12;
				 l_2 = +15; end
		2409: begin l_1 = +12;
				 l_2 = -15; end
		940: begin l_1 = -12;
				 l_2 = +15; end
		1662: begin l_1 = -12;
				 l_2 = -15; end
		1326: begin l_1 = +12;
				 l_2 = +16; end
		2770: begin l_1 = +12;
				 l_2 = -16; end
		579: begin l_1 = -12;
				 l_2 = +16; end
		2023: begin l_1 = -12;
				 l_2 = -16; end
		604: begin l_1 = +12;
				 l_2 = +17; end
		143: begin l_1 = +12;
				 l_2 = -17; end
		3206: begin l_1 = -12;
				 l_2 = +17; end
		2745: begin l_1 = -12;
				 l_2 = -17; end
		2509: begin l_1 = +12;
				 l_2 = +18; end
		1587: begin l_1 = +12;
				 l_2 = -18; end
		1762: begin l_1 = -12;
				 l_2 = +18; end
		840: begin l_1 = -12;
				 l_2 = -18; end
		2970: begin l_1 = +12;
				 l_2 = +19; end
		1126: begin l_1 = +12;
				 l_2 = -19; end
		2223: begin l_1 = -12;
				 l_2 = +19; end
		379: begin l_1 = -12;
				 l_2 = -19; end
		543: begin l_1 = +12;
				 l_2 = +20; end
		204: begin l_1 = +12;
				 l_2 = -20; end
		3145: begin l_1 = -12;
				 l_2 = +20; end
		2806: begin l_1 = -12;
				 l_2 = -20; end
		2387: begin l_1 = +12;
				 l_2 = +21; end
		1709: begin l_1 = +12;
				 l_2 = -21; end
		1640: begin l_1 = -12;
				 l_2 = +21; end
		962: begin l_1 = -12;
				 l_2 = -21; end
		2726: begin l_1 = +12;
				 l_2 = +22; end
		1370: begin l_1 = +12;
				 l_2 = -22; end
		1979: begin l_1 = -12;
				 l_2 = +22; end
		623: begin l_1 = -12;
				 l_2 = -22; end
		55: begin l_1 = +12;
				 l_2 = +23; end
		692: begin l_1 = +12;
				 l_2 = -23; end
		2657: begin l_1 = -12;
				 l_2 = +23; end
		3294: begin l_1 = -12;
				 l_2 = -23; end
		1411: begin l_1 = +12;
				 l_2 = +24; end
		2685: begin l_1 = +12;
				 l_2 = -24; end
		664: begin l_1 = -12;
				 l_2 = +24; end
		1938: begin l_1 = -12;
				 l_2 = -24; end
		2241: begin l_1 = -13;
				 l_2 = +15; end
		1108: begin l_1 = -13;
				 l_2 = -14; end
		386: begin l_1 = +13;
				 l_2 = +15; end
		2963: begin l_1 = -13;
				 l_2 = -15; end
		25: begin l_1 = +13;
				 l_2 = +16; end
		1469: begin l_1 = +13;
				 l_2 = -16; end
		1880: begin l_1 = -13;
				 l_2 = +16; end
		3324: begin l_1 = -13;
				 l_2 = -16; end
		2652: begin l_1 = +13;
				 l_2 = +17; end
		2191: begin l_1 = +13;
				 l_2 = -17; end
		1158: begin l_1 = -13;
				 l_2 = +17; end
		697: begin l_1 = -13;
				 l_2 = -17; end
		1208: begin l_1 = +13;
				 l_2 = +18; end
		286: begin l_1 = +13;
				 l_2 = -18; end
		3063: begin l_1 = -13;
				 l_2 = +18; end
		2141: begin l_1 = -13;
				 l_2 = -18; end
		1669: begin l_1 = +13;
				 l_2 = +19; end
		3174: begin l_1 = +13;
				 l_2 = -19; end
		175: begin l_1 = -13;
				 l_2 = +19; end
		1680: begin l_1 = -13;
				 l_2 = -19; end
		2591: begin l_1 = +13;
				 l_2 = +20; end
		2252: begin l_1 = +13;
				 l_2 = -20; end
		1097: begin l_1 = -13;
				 l_2 = +20; end
		758: begin l_1 = -13;
				 l_2 = -20; end
		1086: begin l_1 = +13;
				 l_2 = +21; end
		408: begin l_1 = +13;
				 l_2 = -21; end
		2941: begin l_1 = -13;
				 l_2 = +21; end
		2263: begin l_1 = -13;
				 l_2 = -21; end
		1425: begin l_1 = +13;
				 l_2 = +22; end
		69: begin l_1 = +13;
				 l_2 = -22; end
		3280: begin l_1 = -13;
				 l_2 = +22; end
		1924: begin l_1 = -13;
				 l_2 = -22; end
		2103: begin l_1 = +13;
				 l_2 = +23; end
		2740: begin l_1 = +13;
				 l_2 = -23; end
		609: begin l_1 = -13;
				 l_2 = +23; end
		1246: begin l_1 = -13;
				 l_2 = -23; end
		110: begin l_1 = +13;
				 l_2 = +24; end
		1384: begin l_1 = +13;
				 l_2 = -24; end
		1965: begin l_1 = -13;
				 l_2 = +24; end
		3239: begin l_1 = -13;
				 l_2 = -24; end
		1133: begin l_1 = -14;
				 l_2 = +16; end
		2216: begin l_1 = -14;
				 l_2 = -15; end
		772: begin l_1 = +14;
				 l_2 = +16; end
		2577: begin l_1 = -14;
				 l_2 = -16; end
		50: begin l_1 = +14;
				 l_2 = +17; end
		2938: begin l_1 = +14;
				 l_2 = -17; end
		411: begin l_1 = -14;
				 l_2 = +17; end
		3299: begin l_1 = -14;
				 l_2 = -17; end
		1955: begin l_1 = +14;
				 l_2 = +18; end
		1033: begin l_1 = +14;
				 l_2 = -18; end
		2316: begin l_1 = -14;
				 l_2 = +18; end
		1394: begin l_1 = -14;
				 l_2 = -18; end
		2416: begin l_1 = +14;
				 l_2 = +19; end
		572: begin l_1 = +14;
				 l_2 = -19; end
		2777: begin l_1 = -14;
				 l_2 = +19; end
		933: begin l_1 = -14;
				 l_2 = -19; end
		3338: begin l_1 = +14;
				 l_2 = +20; end
		2999: begin l_1 = +14;
				 l_2 = -20; end
		350: begin l_1 = -14;
				 l_2 = +20; end
		11: begin l_1 = -14;
				 l_2 = -20; end
		1833: begin l_1 = +14;
				 l_2 = +21; end
		1155: begin l_1 = +14;
				 l_2 = -21; end
		2194: begin l_1 = -14;
				 l_2 = +21; end
		1516: begin l_1 = -14;
				 l_2 = -21; end
		2172: begin l_1 = +14;
				 l_2 = +22; end
		816: begin l_1 = +14;
				 l_2 = -22; end
		2533: begin l_1 = -14;
				 l_2 = +22; end
		1177: begin l_1 = -14;
				 l_2 = -22; end
		2850: begin l_1 = +14;
				 l_2 = +23; end
		138: begin l_1 = +14;
				 l_2 = -23; end
		3211: begin l_1 = -14;
				 l_2 = +23; end
		499: begin l_1 = -14;
				 l_2 = -23; end
		857: begin l_1 = +14;
				 l_2 = +24; end
		2131: begin l_1 = +14;
				 l_2 = -24; end
		1218: begin l_1 = -14;
				 l_2 = +24; end
		2492: begin l_1 = -14;
				 l_2 = -24; end
		2266: begin l_1 = -15;
				 l_2 = +17; end
		1083: begin l_1 = -15;
				 l_2 = -16; end
		1544: begin l_1 = +15;
				 l_2 = +17; end
		1805: begin l_1 = -15;
				 l_2 = -17; end
		100: begin l_1 = +15;
				 l_2 = +18; end
		2527: begin l_1 = +15;
				 l_2 = -18; end
		822: begin l_1 = -15;
				 l_2 = +18; end
		3249: begin l_1 = -15;
				 l_2 = -18; end
		561: begin l_1 = +15;
				 l_2 = +19; end
		2066: begin l_1 = +15;
				 l_2 = -19; end
		1283: begin l_1 = -15;
				 l_2 = +19; end
		2788: begin l_1 = -15;
				 l_2 = -19; end
		1483: begin l_1 = +15;
				 l_2 = +20; end
		1144: begin l_1 = +15;
				 l_2 = -20; end
		2205: begin l_1 = -15;
				 l_2 = +20; end
		1866: begin l_1 = -15;
				 l_2 = -20; end
		3327: begin l_1 = +15;
				 l_2 = +21; end
		2649: begin l_1 = +15;
				 l_2 = -21; end
		700: begin l_1 = -15;
				 l_2 = +21; end
		22: begin l_1 = -15;
				 l_2 = -21; end
		317: begin l_1 = +15;
				 l_2 = +22; end
		2310: begin l_1 = +15;
				 l_2 = -22; end
		1039: begin l_1 = -15;
				 l_2 = +22; end
		3032: begin l_1 = -15;
				 l_2 = -22; end
		995: begin l_1 = +15;
				 l_2 = +23; end
		1632: begin l_1 = +15;
				 l_2 = -23; end
		1717: begin l_1 = -15;
				 l_2 = +23; end
		2354: begin l_1 = -15;
				 l_2 = -23; end
		2351: begin l_1 = +15;
				 l_2 = +24; end
		276: begin l_1 = +15;
				 l_2 = -24; end
		3073: begin l_1 = -15;
				 l_2 = +24; end
		998: begin l_1 = -15;
				 l_2 = -24; end
		1183: begin l_1 = -16;
				 l_2 = +18; end
		2166: begin l_1 = -16;
				 l_2 = -17; end
		3088: begin l_1 = +16;
				 l_2 = +18; end
		261: begin l_1 = -16;
				 l_2 = -18; end
		200: begin l_1 = +16;
				 l_2 = +19; end
		1705: begin l_1 = +16;
				 l_2 = -19; end
		1644: begin l_1 = -16;
				 l_2 = +19; end
		3149: begin l_1 = -16;
				 l_2 = -19; end
		1122: begin l_1 = +16;
				 l_2 = +20; end
		783: begin l_1 = +16;
				 l_2 = -20; end
		2566: begin l_1 = -16;
				 l_2 = +20; end
		2227: begin l_1 = -16;
				 l_2 = -20; end
		2966: begin l_1 = +16;
				 l_2 = +21; end
		2288: begin l_1 = +16;
				 l_2 = -21; end
		1061: begin l_1 = -16;
				 l_2 = +21; end
		383: begin l_1 = -16;
				 l_2 = -21; end
		3305: begin l_1 = +16;
				 l_2 = +22; end
		1949: begin l_1 = +16;
				 l_2 = -22; end
		1400: begin l_1 = -16;
				 l_2 = +22; end
		44: begin l_1 = -16;
				 l_2 = -22; end
		634: begin l_1 = +16;
				 l_2 = +23; end
		1271: begin l_1 = +16;
				 l_2 = -23; end
		2078: begin l_1 = -16;
				 l_2 = +23; end
		2715: begin l_1 = -16;
				 l_2 = -23; end
		1990: begin l_1 = +16;
				 l_2 = +24; end
		3264: begin l_1 = +16;
				 l_2 = -24; end
		85: begin l_1 = -16;
				 l_2 = +24; end
		1359: begin l_1 = -16;
				 l_2 = -24; end
		2366: begin l_1 = -17;
				 l_2 = +19; end
		983: begin l_1 = -17;
				 l_2 = -18; end
		2827: begin l_1 = +17;
				 l_2 = +19; end
		522: begin l_1 = -17;
				 l_2 = -19; end
		400: begin l_1 = +17;
				 l_2 = +20; end
		61: begin l_1 = +17;
				 l_2 = -20; end
		3288: begin l_1 = -17;
				 l_2 = +20; end
		2949: begin l_1 = -17;
				 l_2 = -20; end
		2244: begin l_1 = +17;
				 l_2 = +21; end
		1566: begin l_1 = +17;
				 l_2 = -21; end
		1783: begin l_1 = -17;
				 l_2 = +21; end
		1105: begin l_1 = -17;
				 l_2 = -21; end
		2583: begin l_1 = +17;
				 l_2 = +22; end
		1227: begin l_1 = +17;
				 l_2 = -22; end
		2122: begin l_1 = -17;
				 l_2 = +22; end
		766: begin l_1 = -17;
				 l_2 = -22; end
		3261: begin l_1 = +17;
				 l_2 = +23; end
		549: begin l_1 = +17;
				 l_2 = -23; end
		2800: begin l_1 = -17;
				 l_2 = +23; end
		88: begin l_1 = -17;
				 l_2 = -23; end
		1268: begin l_1 = +17;
				 l_2 = +24; end
		2542: begin l_1 = +17;
				 l_2 = -24; end
		807: begin l_1 = -17;
				 l_2 = +24; end
		2081: begin l_1 = -17;
				 l_2 = -24; end
		1383: begin l_1 = -18;
				 l_2 = +20; end
		1966: begin l_1 = -18;
				 l_2 = -19; end
		2305: begin l_1 = +18;
				 l_2 = +20; end
		1044: begin l_1 = -18;
				 l_2 = -20; end
		800: begin l_1 = +18;
				 l_2 = +21; end
		122: begin l_1 = +18;
				 l_2 = -21; end
		3227: begin l_1 = -18;
				 l_2 = +21; end
		2549: begin l_1 = -18;
				 l_2 = -21; end
		1139: begin l_1 = +18;
				 l_2 = +22; end
		3132: begin l_1 = +18;
				 l_2 = -22; end
		217: begin l_1 = -18;
				 l_2 = +22; end
		2210: begin l_1 = -18;
				 l_2 = -22; end
		1817: begin l_1 = +18;
				 l_2 = +23; end
		2454: begin l_1 = +18;
				 l_2 = -23; end
		895: begin l_1 = -18;
				 l_2 = +23; end
		1532: begin l_1 = -18;
				 l_2 = -23; end
		3173: begin l_1 = +18;
				 l_2 = +24; end
		1098: begin l_1 = +18;
				 l_2 = -24; end
		2251: begin l_1 = -18;
				 l_2 = +24; end
		176: begin l_1 = -18;
				 l_2 = -24; end
		2766: begin l_1 = -19;
				 l_2 = +21; end
		583: begin l_1 = -19;
				 l_2 = -20; end
		1261: begin l_1 = +19;
				 l_2 = +21; end
		2088: begin l_1 = -19;
				 l_2 = -21; end
		1600: begin l_1 = +19;
				 l_2 = +22; end
		244: begin l_1 = +19;
				 l_2 = -22; end
		3105: begin l_1 = -19;
				 l_2 = +22; end
		1749: begin l_1 = -19;
				 l_2 = -22; end
		2278: begin l_1 = +19;
				 l_2 = +23; end
		2915: begin l_1 = +19;
				 l_2 = -23; end
		434: begin l_1 = -19;
				 l_2 = +23; end
		1071: begin l_1 = -19;
				 l_2 = -23; end
		285: begin l_1 = +19;
				 l_2 = +24; end
		1559: begin l_1 = +19;
				 l_2 = -24; end
		1790: begin l_1 = -19;
				 l_2 = +24; end
		3064: begin l_1 = -19;
				 l_2 = -24; end
		2183: begin l_1 = -20;
				 l_2 = +22; end
		1166: begin l_1 = -20;
				 l_2 = -21; end
		2522: begin l_1 = +20;
				 l_2 = +22; end
		827: begin l_1 = -20;
				 l_2 = -22; end
		3200: begin l_1 = +20;
				 l_2 = +23; end
		488: begin l_1 = +20;
				 l_2 = -23; end
		2861: begin l_1 = -20;
				 l_2 = +23; end
		149: begin l_1 = -20;
				 l_2 = -23; end
		1207: begin l_1 = +20;
				 l_2 = +24; end
		2481: begin l_1 = +20;
				 l_2 = -24; end
		868: begin l_1 = -20;
				 l_2 = +24; end
		2142: begin l_1 = -20;
				 l_2 = -24; end
		1017: begin l_1 = -21;
				 l_2 = +23; end
		2332: begin l_1 = -21;
				 l_2 = -22; end
		1695: begin l_1 = +21;
				 l_2 = +23; end
		1654: begin l_1 = -21;
				 l_2 = -23; end
		3051: begin l_1 = +21;
				 l_2 = +24; end
		976: begin l_1 = +21;
				 l_2 = -24; end
		2373: begin l_1 = -21;
				 l_2 = +24; end
		298: begin l_1 = -21;
				 l_2 = -24; end
		2034: begin l_1 = -22;
				 l_2 = +24; end
		1315: begin l_1 = -22;
				 l_2 = -23; end
		41: begin l_1 = +22;
				 l_2 = +24; end
		3308: begin l_1 = -22;
				 l_2 = -24; end
		719: begin l_1 = +23;
				 l_2 = +24; end
		2630: begin l_1 = -23;
				 l_2 = -24; end
		default: begin l_1 = 0;
					   l_2 = 0; end
	endcase
end

endmodule

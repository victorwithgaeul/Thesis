// Product (AN) Code SEC l-LUT
// SEC_lLUT28bits.v
// Received single error location l, output remainder r.
module SEC_lLUT28bits(l, r);
input	signed	[6:0]	l;
output	reg	[14:0]	r;
always@(*) begin
	case(l)
		1: r = 1;
		-1: r = 17618;
		2: r = 2;
		-2: r = 17617;
		3: r = 4;
		-3: r = 17615;
		4: r = 8;
		-4: r = 17611;
		5: r = 16;
		-5: r = 17603;
		6: r = 32;
		-6: r = 17587;
		7: r = 64;
		-7: r = 17555;
		8: r = 128;
		-8: r = 17491;
		9: r = 256;
		-9: r = 17363;
		10: r = 512;
		-10: r = 17107;
		11: r = 1024;
		-11: r = 16595;
		12: r = 2048;
		-12: r = 15571;
		13: r = 4096;
		-13: r = 13523;
		14: r = 8192;
		-14: r = 9427;
		15: r = 16384;
		-15: r = 1235;
		16: r = 15149;
		-16: r = 2470;
		17: r = 12679;
		-17: r = 4940;
		18: r = 7739;
		-18: r = 9880;
		19: r = 15478;
		-19: r = 2141;
		20: r = 13337;
		-20: r = 4282;
		21: r = 9055;
		-21: r = 8564;
		22: r = 491;
		-22: r = 17128;
		23: r = 982;
		-23: r = 16637;
		24: r = 1964;
		-24: r = 15655;
		25: r = 3928;
		-25: r = 13691;
		26: r = 7856;
		-26: r = 9763;
		27: r = 15712;
		-27: r = 1907;
		28: r = 13805;
		-28: r = 3814;
		29: r = 9991;
		-29: r = 7628;
		30: r = 2363;
		-30: r = 15256;
		31: r = 4726;
		-31: r = 12893;
		32: r = 9452;
		-32: r = 8167;
		33: r = 1285;
		-33: r = 16334;
		34: r = 2570;
		-34: r = 15049;
		35: r = 5140;
		-35: r = 12479;
		36: r = 10280;
		-36: r = 7339;
		37: r = 2941;
		-37: r = 14678;
		38: r = 5882;
		-38: r = 11737;
		39: r = 11764;
		-39: r = 5855;
		40: r = 5909;
		-40: r = 11710;
		41: r = 11818;
		-41: r = 5801;
		42: r = 6017;
		-42: r = 11602;
		43: r = 12034;
		-43: r = 5585;
		default: r = 0;
	endcase
end

endmodule

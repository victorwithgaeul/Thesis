// Product (AN) Code SEC_LUT_Decoder
// SEC_LUT_Decoder24bits.v
// Received codeword W = AN + e, e is single arithmetic weight error (AWE), +2^i or -2^i.
module SEC_LUT_Decoder24bits(W, N);
input 	[37:0]	W;
output	[23:0]	N;
parameter A = 13837;

wire 	[23:0]	Q;
wire 	[13:0]	R;
assign Q = W / A;
assign R = W - (A * Q);

reg	signed	[38:0]	Delta;
always@(*) begin
	case(R)
		1: Delta = 39'sb000000000000000000000000000000000000001;
		13836: Delta = 39'sb111111111111111111111111111111111111111;
		2: Delta = 39'sb000000000000000000000000000000000000010;
		13835: Delta = 39'sb111111111111111111111111111111111111110;
		4: Delta = 39'sb000000000000000000000000000000000000100;
		13833: Delta = 39'sb111111111111111111111111111111111111100;
		8: Delta = 39'sb000000000000000000000000000000000001000;
		13829: Delta = 39'sb111111111111111111111111111111111111000;
		16: Delta = 39'sb000000000000000000000000000000000010000;
		13821: Delta = 39'sb111111111111111111111111111111111110000;
		32: Delta = 39'sb000000000000000000000000000000000100000;
		13805: Delta = 39'sb111111111111111111111111111111111100000;
		64: Delta = 39'sb000000000000000000000000000000001000000;
		13773: Delta = 39'sb111111111111111111111111111111111000000;
		128: Delta = 39'sb000000000000000000000000000000010000000;
		13709: Delta = 39'sb111111111111111111111111111111110000000;
		256: Delta = 39'sb000000000000000000000000000000100000000;
		13581: Delta = 39'sb111111111111111111111111111111100000000;
		512: Delta = 39'sb000000000000000000000000000001000000000;
		13325: Delta = 39'sb111111111111111111111111111111000000000;
		1024: Delta = 39'sb000000000000000000000000000010000000000;
		12813: Delta = 39'sb111111111111111111111111111110000000000;
		2048: Delta = 39'sb000000000000000000000000000100000000000;
		11789: Delta = 39'sb111111111111111111111111111100000000000;
		4096: Delta = 39'sb000000000000000000000000001000000000000;
		9741: Delta = 39'sb111111111111111111111111111000000000000;
		8192: Delta = 39'sb000000000000000000000000010000000000000;
		5645: Delta = 39'sb111111111111111111111111110000000000000;
		2547: Delta = 39'sb000000000000000000000000100000000000000;
		11290: Delta = 39'sb111111111111111111111111100000000000000;
		5094: Delta = 39'sb000000000000000000000001000000000000000;
		8743: Delta = 39'sb111111111111111111111111000000000000000;
		10188: Delta = 39'sb000000000000000000000010000000000000000;
		3649: Delta = 39'sb111111111111111111111110000000000000000;
		6539: Delta = 39'sb000000000000000000000100000000000000000;
		7298: Delta = 39'sb111111111111111111111100000000000000000;
		13078: Delta = 39'sb000000000000000000001000000000000000000;
		759: Delta = 39'sb111111111111111111111000000000000000000;
		12319: Delta = 39'sb000000000000000000010000000000000000000;
		1518: Delta = 39'sb111111111111111111110000000000000000000;
		10801: Delta = 39'sb000000000000000000100000000000000000000;
		3036: Delta = 39'sb111111111111111111100000000000000000000;
		7765: Delta = 39'sb000000000000000001000000000000000000000;
		6072: Delta = 39'sb111111111111111111000000000000000000000;
		1693: Delta = 39'sb000000000000000010000000000000000000000;
		12144: Delta = 39'sb111111111111111110000000000000000000000;
		3386: Delta = 39'sb000000000000000100000000000000000000000;
		10451: Delta = 39'sb111111111111111100000000000000000000000;
		6772: Delta = 39'sb000000000000001000000000000000000000000;
		7065: Delta = 39'sb111111111111111000000000000000000000000;
		13544: Delta = 39'sb000000000000010000000000000000000000000;
		293: Delta = 39'sb111111111111110000000000000000000000000;
		13251: Delta = 39'sb000000000000100000000000000000000000000;
		586: Delta = 39'sb111111111111100000000000000000000000000;
		12665: Delta = 39'sb000000000001000000000000000000000000000;
		1172: Delta = 39'sb111111111111000000000000000000000000000;
		11493: Delta = 39'sb000000000010000000000000000000000000000;
		2344: Delta = 39'sb111111111110000000000000000000000000000;
		9149: Delta = 39'sb000000000100000000000000000000000000000;
		4688: Delta = 39'sb111111111100000000000000000000000000000;
		4461: Delta = 39'sb000000001000000000000000000000000000000;
		9376: Delta = 39'sb111111111000000000000000000000000000000;
		8922: Delta = 39'sb000000010000000000000000000000000000000;
		4915: Delta = 39'sb111111110000000000000000000000000000000;
		4007: Delta = 39'sb000000100000000000000000000000000000000;
		9830: Delta = 39'sb111111100000000000000000000000000000000;
		8014: Delta = 39'sb000001000000000000000000000000000000000;
		5823: Delta = 39'sb111111000000000000000000000000000000000;
		2191: Delta = 39'sb000010000000000000000000000000000000000;
		11646: Delta = 39'sb111110000000000000000000000000000000000;
		4382: Delta = 39'sb000100000000000000000000000000000000000;
		9455: Delta = 39'sb111100000000000000000000000000000000000;
		8764: Delta = 39'sb001000000000000000000000000000000000000;
		5073: Delta = 39'sb111000000000000000000000000000000000000;
		3691: Delta = 39'sb010000000000000000000000000000000000000;
		10146: Delta = 39'sb110000000000000000000000000000000000000;
		default: Delta =39'sb0;
	endcase
end

assign N = (W - Delta) / A;

endmodule

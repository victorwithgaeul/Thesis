// Product (AN) Code DEC_LUT_Decoder
// DEC_LUT_Decoder24bits.v
// Received codeword W = AN + E, E is double AWE (E = e1 + e2), +2^i or -2^i.
module DEC_LUT_Decoder24bits(W, N);
input 	[37:0]	W;
output	[23:0]	N;
parameter A = 13837;

wire 	[23:0]	Q;
wire 	[13:0]	R;
assign Q = W / A;
assign R = W - (A * Q);

reg	signed	[38:0]	Delta;
always@(*) begin
	case(R)
		1: Delta = 39'sb000000000000000000000000000000000000001;
		13836: Delta = 39'sb111111111111111111111111111111111111111;
		2: Delta = 39'sb000000000000000000000000000000000000010;
		13835: Delta = 39'sb111111111111111111111111111111111111110;
		4: Delta = 39'sb000000000000000000000000000000000000100;
		13833: Delta = 39'sb111111111111111111111111111111111111100;
		8: Delta = 39'sb000000000000000000000000000000000001000;
		13829: Delta = 39'sb111111111111111111111111111111111111000;
		16: Delta = 39'sb000000000000000000000000000000000010000;
		13821: Delta = 39'sb111111111111111111111111111111111110000;
		32: Delta = 39'sb000000000000000000000000000000000100000;
		13805: Delta = 39'sb111111111111111111111111111111111100000;
		64: Delta = 39'sb000000000000000000000000000000001000000;
		13773: Delta = 39'sb111111111111111111111111111111111000000;
		128: Delta = 39'sb000000000000000000000000000000010000000;
		13709: Delta = 39'sb111111111111111111111111111111110000000;
		256: Delta = 39'sb000000000000000000000000000000100000000;
		13581: Delta = 39'sb111111111111111111111111111111100000000;
		512: Delta = 39'sb000000000000000000000000000001000000000;
		13325: Delta = 39'sb111111111111111111111111111111000000000;
		1024: Delta = 39'sb000000000000000000000000000010000000000;
		12813: Delta = 39'sb111111111111111111111111111110000000000;
		2048: Delta = 39'sb000000000000000000000000000100000000000;
		11789: Delta = 39'sb111111111111111111111111111100000000000;
		4096: Delta = 39'sb000000000000000000000000001000000000000;
		9741: Delta = 39'sb111111111111111111111111111000000000000;
		8192: Delta = 39'sb000000000000000000000000010000000000000;
		5645: Delta = 39'sb111111111111111111111111110000000000000;
		2547: Delta = 39'sb000000000000000000000000100000000000000;
		11290: Delta = 39'sb111111111111111111111111100000000000000;
		5094: Delta = 39'sb000000000000000000000001000000000000000;
		8743: Delta = 39'sb111111111111111111111111000000000000000;
		10188: Delta = 39'sb000000000000000000000010000000000000000;
		3649: Delta = 39'sb111111111111111111111110000000000000000;
		6539: Delta = 39'sb000000000000000000000100000000000000000;
		7298: Delta = 39'sb111111111111111111111100000000000000000;
		13078: Delta = 39'sb000000000000000000001000000000000000000;
		759: Delta = 39'sb111111111111111111111000000000000000000;
		12319: Delta = 39'sb000000000000000000010000000000000000000;
		1518: Delta = 39'sb111111111111111111110000000000000000000;
		10801: Delta = 39'sb000000000000000000100000000000000000000;
		3036: Delta = 39'sb111111111111111111100000000000000000000;
		7765: Delta = 39'sb000000000000000001000000000000000000000;
		6072: Delta = 39'sb111111111111111111000000000000000000000;
		1693: Delta = 39'sb000000000000000010000000000000000000000;
		12144: Delta = 39'sb111111111111111110000000000000000000000;
		3386: Delta = 39'sb000000000000000100000000000000000000000;
		10451: Delta = 39'sb111111111111111100000000000000000000000;
		6772: Delta = 39'sb000000000000001000000000000000000000000;
		7065: Delta = 39'sb111111111111111000000000000000000000000;
		13544: Delta = 39'sb000000000000010000000000000000000000000;
		293: Delta = 39'sb111111111111110000000000000000000000000;
		13251: Delta = 39'sb000000000000100000000000000000000000000;
		586: Delta = 39'sb111111111111100000000000000000000000000;
		12665: Delta = 39'sb000000000001000000000000000000000000000;
		1172: Delta = 39'sb111111111111000000000000000000000000000;
		11493: Delta = 39'sb000000000010000000000000000000000000000;
		2344: Delta = 39'sb111111111110000000000000000000000000000;
		9149: Delta = 39'sb000000000100000000000000000000000000000;
		4688: Delta = 39'sb111111111100000000000000000000000000000;
		4461: Delta = 39'sb000000001000000000000000000000000000000;
		9376: Delta = 39'sb111111111000000000000000000000000000000;
		8922: Delta = 39'sb000000010000000000000000000000000000000;
		4915: Delta = 39'sb111111110000000000000000000000000000000;
		4007: Delta = 39'sb000000100000000000000000000000000000000;
		9830: Delta = 39'sb111111100000000000000000000000000000000;
		8014: Delta = 39'sb000001000000000000000000000000000000000;
		5823: Delta = 39'sb111111000000000000000000000000000000000;
		2191: Delta = 39'sb000010000000000000000000000000000000000;
		11646: Delta = 39'sb111110000000000000000000000000000000000;
		4382: Delta = 39'sb000100000000000000000000000000000000000;
		9455: Delta = 39'sb111100000000000000000000000000000000000;
		8764: Delta = 39'sb001000000000000000000000000000000000000;
		5073: Delta = 39'sb111000000000000000000000000000000000000;
		3691: Delta = 39'sb010000000000000000000000000000000000000;
		10146: Delta = 39'sb110000000000000000000000000000000000000;
		3: Delta = 39'sb000000000000000000000000000000000000011;
		13834: Delta = 39'sb111111111111111111111111111111111111101;
		5: Delta = 39'sb000000000000000000000000000000000000101;
		13832: Delta = 39'sb111111111111111111111111111111111111011;
		9: Delta = 39'sb000000000000000000000000000000000001001;
		13830: Delta = 39'sb111111111111111111111111111111111111001;
		7: Delta = 39'sb000000000000000000000000000000000000111;
		13828: Delta = 39'sb111111111111111111111111111111111110111;
		17: Delta = 39'sb000000000000000000000000000000000010001;
		13822: Delta = 39'sb111111111111111111111111111111111110001;
		15: Delta = 39'sb000000000000000000000000000000000001111;
		13820: Delta = 39'sb111111111111111111111111111111111101111;
		33: Delta = 39'sb000000000000000000000000000000000100001;
		13806: Delta = 39'sb111111111111111111111111111111111100001;
		31: Delta = 39'sb000000000000000000000000000000000011111;
		13804: Delta = 39'sb111111111111111111111111111111111011111;
		65: Delta = 39'sb000000000000000000000000000000001000001;
		13774: Delta = 39'sb111111111111111111111111111111111000001;
		63: Delta = 39'sb000000000000000000000000000000000111111;
		13772: Delta = 39'sb111111111111111111111111111111110111111;
		129: Delta = 39'sb000000000000000000000000000000010000001;
		13710: Delta = 39'sb111111111111111111111111111111110000001;
		127: Delta = 39'sb000000000000000000000000000000001111111;
		13708: Delta = 39'sb111111111111111111111111111111101111111;
		257: Delta = 39'sb000000000000000000000000000000100000001;
		13582: Delta = 39'sb111111111111111111111111111111100000001;
		255: Delta = 39'sb000000000000000000000000000000011111111;
		13580: Delta = 39'sb111111111111111111111111111111011111111;
		513: Delta = 39'sb000000000000000000000000000001000000001;
		13326: Delta = 39'sb111111111111111111111111111111000000001;
		511: Delta = 39'sb000000000000000000000000000000111111111;
		13324: Delta = 39'sb111111111111111111111111111110111111111;
		1025: Delta = 39'sb000000000000000000000000000010000000001;
		12814: Delta = 39'sb111111111111111111111111111110000000001;
		1023: Delta = 39'sb000000000000000000000000000001111111111;
		12812: Delta = 39'sb111111111111111111111111111101111111111;
		2049: Delta = 39'sb000000000000000000000000000100000000001;
		11790: Delta = 39'sb111111111111111111111111111100000000001;
		2047: Delta = 39'sb000000000000000000000000000011111111111;
		11788: Delta = 39'sb111111111111111111111111111011111111111;
		4097: Delta = 39'sb000000000000000000000000001000000000001;
		9742: Delta = 39'sb111111111111111111111111111000000000001;
		4095: Delta = 39'sb000000000000000000000000000111111111111;
		9740: Delta = 39'sb111111111111111111111111110111111111111;
		8193: Delta = 39'sb000000000000000000000000010000000000001;
		5646: Delta = 39'sb111111111111111111111111110000000000001;
		8191: Delta = 39'sb000000000000000000000000001111111111111;
		5644: Delta = 39'sb111111111111111111111111101111111111111;
		2548: Delta = 39'sb000000000000000000000000100000000000001;
		11291: Delta = 39'sb111111111111111111111111100000000000001;
		2546: Delta = 39'sb000000000000000000000000011111111111111;
		11289: Delta = 39'sb111111111111111111111111011111111111111;
		5095: Delta = 39'sb000000000000000000000001000000000000001;
		8744: Delta = 39'sb111111111111111111111111000000000000001;
		5093: Delta = 39'sb000000000000000000000000111111111111111;
		8742: Delta = 39'sb111111111111111111111110111111111111111;
		10189: Delta = 39'sb000000000000000000000010000000000000001;
		3650: Delta = 39'sb111111111111111111111110000000000000001;
		10187: Delta = 39'sb000000000000000000000001111111111111111;
		3648: Delta = 39'sb111111111111111111111101111111111111111;
		6540: Delta = 39'sb000000000000000000000100000000000000001;
		7299: Delta = 39'sb111111111111111111111100000000000000001;
		6538: Delta = 39'sb000000000000000000000011111111111111111;
		7297: Delta = 39'sb111111111111111111111011111111111111111;
		13079: Delta = 39'sb000000000000000000001000000000000000001;
		760: Delta = 39'sb111111111111111111111000000000000000001;
		13077: Delta = 39'sb000000000000000000000111111111111111111;
		758: Delta = 39'sb111111111111111111110111111111111111111;
		12320: Delta = 39'sb000000000000000000010000000000000000001;
		1519: Delta = 39'sb111111111111111111110000000000000000001;
		12318: Delta = 39'sb000000000000000000001111111111111111111;
		1517: Delta = 39'sb111111111111111111101111111111111111111;
		10802: Delta = 39'sb000000000000000000100000000000000000001;
		3037: Delta = 39'sb111111111111111111100000000000000000001;
		10800: Delta = 39'sb000000000000000000011111111111111111111;
		3035: Delta = 39'sb111111111111111111011111111111111111111;
		7766: Delta = 39'sb000000000000000001000000000000000000001;
		6073: Delta = 39'sb111111111111111111000000000000000000001;
		7764: Delta = 39'sb000000000000000000111111111111111111111;
		6071: Delta = 39'sb111111111111111110111111111111111111111;
		1694: Delta = 39'sb000000000000000010000000000000000000001;
		12145: Delta = 39'sb111111111111111110000000000000000000001;
		1692: Delta = 39'sb000000000000000001111111111111111111111;
		12143: Delta = 39'sb111111111111111101111111111111111111111;
		3387: Delta = 39'sb000000000000000100000000000000000000001;
		10452: Delta = 39'sb111111111111111100000000000000000000001;
		3385: Delta = 39'sb000000000000000011111111111111111111111;
		10450: Delta = 39'sb111111111111111011111111111111111111111;
		6773: Delta = 39'sb000000000000001000000000000000000000001;
		7066: Delta = 39'sb111111111111111000000000000000000000001;
		6771: Delta = 39'sb000000000000000111111111111111111111111;
		7064: Delta = 39'sb111111111111110111111111111111111111111;
		13545: Delta = 39'sb000000000000010000000000000000000000001;
		294: Delta = 39'sb111111111111110000000000000000000000001;
		13543: Delta = 39'sb000000000000001111111111111111111111111;
		292: Delta = 39'sb111111111111101111111111111111111111111;
		13252: Delta = 39'sb000000000000100000000000000000000000001;
		587: Delta = 39'sb111111111111100000000000000000000000001;
		13250: Delta = 39'sb000000000000011111111111111111111111111;
		585: Delta = 39'sb111111111111011111111111111111111111111;
		12666: Delta = 39'sb000000000001000000000000000000000000001;
		1173: Delta = 39'sb111111111111000000000000000000000000001;
		12664: Delta = 39'sb000000000000111111111111111111111111111;
		1171: Delta = 39'sb111111111110111111111111111111111111111;
		11494: Delta = 39'sb000000000010000000000000000000000000001;
		2345: Delta = 39'sb111111111110000000000000000000000000001;
		11492: Delta = 39'sb000000000001111111111111111111111111111;
		2343: Delta = 39'sb111111111101111111111111111111111111111;
		9150: Delta = 39'sb000000000100000000000000000000000000001;
		4689: Delta = 39'sb111111111100000000000000000000000000001;
		9148: Delta = 39'sb000000000011111111111111111111111111111;
		4687: Delta = 39'sb111111111011111111111111111111111111111;
		4462: Delta = 39'sb000000001000000000000000000000000000001;
		9377: Delta = 39'sb111111111000000000000000000000000000001;
		4460: Delta = 39'sb000000000111111111111111111111111111111;
		9375: Delta = 39'sb111111110111111111111111111111111111111;
		8923: Delta = 39'sb000000010000000000000000000000000000001;
		4916: Delta = 39'sb111111110000000000000000000000000000001;
		8921: Delta = 39'sb000000001111111111111111111111111111111;
		4914: Delta = 39'sb111111101111111111111111111111111111111;
		4008: Delta = 39'sb000000100000000000000000000000000000001;
		9831: Delta = 39'sb111111100000000000000000000000000000001;
		4006: Delta = 39'sb000000011111111111111111111111111111111;
		9829: Delta = 39'sb111111011111111111111111111111111111111;
		8015: Delta = 39'sb000001000000000000000000000000000000001;
		5824: Delta = 39'sb111111000000000000000000000000000000001;
		8013: Delta = 39'sb000000111111111111111111111111111111111;
		5822: Delta = 39'sb111110111111111111111111111111111111111;
		2192: Delta = 39'sb000010000000000000000000000000000000001;
		11647: Delta = 39'sb111110000000000000000000000000000000001;
		2190: Delta = 39'sb000001111111111111111111111111111111111;
		11645: Delta = 39'sb111101111111111111111111111111111111111;
		4383: Delta = 39'sb000100000000000000000000000000000000001;
		9456: Delta = 39'sb111100000000000000000000000000000000001;
		4381: Delta = 39'sb000011111111111111111111111111111111111;
		9454: Delta = 39'sb111011111111111111111111111111111111111;
		8765: Delta = 39'sb001000000000000000000000000000000000001;
		5074: Delta = 39'sb111000000000000000000000000000000000001;
		8763: Delta = 39'sb000111111111111111111111111111111111111;
		5072: Delta = 39'sb110111111111111111111111111111111111111;
		3692: Delta = 39'sb010000000000000000000000000000000000001;
		10147: Delta = 39'sb110000000000000000000000000000000000001;
		3690: Delta = 39'sb001111111111111111111111111111111111111;
		10145: Delta = 39'sb101111111111111111111111111111111111111;
		6: Delta = 39'sb000000000000000000000000000000000000110;
		13831: Delta = 39'sb111111111111111111111111111111111111010;
		10: Delta = 39'sb000000000000000000000000000000000001010;
		13827: Delta = 39'sb111111111111111111111111111111111110110;
		18: Delta = 39'sb000000000000000000000000000000000010010;
		13823: Delta = 39'sb111111111111111111111111111111111110010;
		14: Delta = 39'sb000000000000000000000000000000000001110;
		13819: Delta = 39'sb111111111111111111111111111111111101110;
		34: Delta = 39'sb000000000000000000000000000000000100010;
		13807: Delta = 39'sb111111111111111111111111111111111100010;
		30: Delta = 39'sb000000000000000000000000000000000011110;
		13803: Delta = 39'sb111111111111111111111111111111111011110;
		66: Delta = 39'sb000000000000000000000000000000001000010;
		13775: Delta = 39'sb111111111111111111111111111111111000010;
		62: Delta = 39'sb000000000000000000000000000000000111110;
		13771: Delta = 39'sb111111111111111111111111111111110111110;
		130: Delta = 39'sb000000000000000000000000000000010000010;
		13711: Delta = 39'sb111111111111111111111111111111110000010;
		126: Delta = 39'sb000000000000000000000000000000001111110;
		13707: Delta = 39'sb111111111111111111111111111111101111110;
		258: Delta = 39'sb000000000000000000000000000000100000010;
		13583: Delta = 39'sb111111111111111111111111111111100000010;
		254: Delta = 39'sb000000000000000000000000000000011111110;
		13579: Delta = 39'sb111111111111111111111111111111011111110;
		514: Delta = 39'sb000000000000000000000000000001000000010;
		13327: Delta = 39'sb111111111111111111111111111111000000010;
		510: Delta = 39'sb000000000000000000000000000000111111110;
		13323: Delta = 39'sb111111111111111111111111111110111111110;
		1026: Delta = 39'sb000000000000000000000000000010000000010;
		12815: Delta = 39'sb111111111111111111111111111110000000010;
		1022: Delta = 39'sb000000000000000000000000000001111111110;
		12811: Delta = 39'sb111111111111111111111111111101111111110;
		2050: Delta = 39'sb000000000000000000000000000100000000010;
		11791: Delta = 39'sb111111111111111111111111111100000000010;
		2046: Delta = 39'sb000000000000000000000000000011111111110;
		11787: Delta = 39'sb111111111111111111111111111011111111110;
		4098: Delta = 39'sb000000000000000000000000001000000000010;
		9743: Delta = 39'sb111111111111111111111111111000000000010;
		4094: Delta = 39'sb000000000000000000000000000111111111110;
		9739: Delta = 39'sb111111111111111111111111110111111111110;
		8194: Delta = 39'sb000000000000000000000000010000000000010;
		5647: Delta = 39'sb111111111111111111111111110000000000010;
		8190: Delta = 39'sb000000000000000000000000001111111111110;
		5643: Delta = 39'sb111111111111111111111111101111111111110;
		2549: Delta = 39'sb000000000000000000000000100000000000010;
		11292: Delta = 39'sb111111111111111111111111100000000000010;
		2545: Delta = 39'sb000000000000000000000000011111111111110;
		11288: Delta = 39'sb111111111111111111111111011111111111110;
		5096: Delta = 39'sb000000000000000000000001000000000000010;
		8745: Delta = 39'sb111111111111111111111111000000000000010;
		5092: Delta = 39'sb000000000000000000000000111111111111110;
		8741: Delta = 39'sb111111111111111111111110111111111111110;
		10190: Delta = 39'sb000000000000000000000010000000000000010;
		3651: Delta = 39'sb111111111111111111111110000000000000010;
		10186: Delta = 39'sb000000000000000000000001111111111111110;
		3647: Delta = 39'sb111111111111111111111101111111111111110;
		6541: Delta = 39'sb000000000000000000000100000000000000010;
		7300: Delta = 39'sb111111111111111111111100000000000000010;
		6537: Delta = 39'sb000000000000000000000011111111111111110;
		7296: Delta = 39'sb111111111111111111111011111111111111110;
		13080: Delta = 39'sb000000000000000000001000000000000000010;
		761: Delta = 39'sb111111111111111111111000000000000000010;
		13076: Delta = 39'sb000000000000000000000111111111111111110;
		757: Delta = 39'sb111111111111111111110111111111111111110;
		12321: Delta = 39'sb000000000000000000010000000000000000010;
		1520: Delta = 39'sb111111111111111111110000000000000000010;
		12317: Delta = 39'sb000000000000000000001111111111111111110;
		1516: Delta = 39'sb111111111111111111101111111111111111110;
		10803: Delta = 39'sb000000000000000000100000000000000000010;
		3038: Delta = 39'sb111111111111111111100000000000000000010;
		10799: Delta = 39'sb000000000000000000011111111111111111110;
		3034: Delta = 39'sb111111111111111111011111111111111111110;
		7767: Delta = 39'sb000000000000000001000000000000000000010;
		6074: Delta = 39'sb111111111111111111000000000000000000010;
		7763: Delta = 39'sb000000000000000000111111111111111111110;
		6070: Delta = 39'sb111111111111111110111111111111111111110;
		1695: Delta = 39'sb000000000000000010000000000000000000010;
		12146: Delta = 39'sb111111111111111110000000000000000000010;
		1691: Delta = 39'sb000000000000000001111111111111111111110;
		12142: Delta = 39'sb111111111111111101111111111111111111110;
		3388: Delta = 39'sb000000000000000100000000000000000000010;
		10453: Delta = 39'sb111111111111111100000000000000000000010;
		3384: Delta = 39'sb000000000000000011111111111111111111110;
		10449: Delta = 39'sb111111111111111011111111111111111111110;
		6774: Delta = 39'sb000000000000001000000000000000000000010;
		7067: Delta = 39'sb111111111111111000000000000000000000010;
		6770: Delta = 39'sb000000000000000111111111111111111111110;
		7063: Delta = 39'sb111111111111110111111111111111111111110;
		13546: Delta = 39'sb000000000000010000000000000000000000010;
		295: Delta = 39'sb111111111111110000000000000000000000010;
		13542: Delta = 39'sb000000000000001111111111111111111111110;
		291: Delta = 39'sb111111111111101111111111111111111111110;
		13253: Delta = 39'sb000000000000100000000000000000000000010;
		588: Delta = 39'sb111111111111100000000000000000000000010;
		13249: Delta = 39'sb000000000000011111111111111111111111110;
		584: Delta = 39'sb111111111111011111111111111111111111110;
		12667: Delta = 39'sb000000000001000000000000000000000000010;
		1174: Delta = 39'sb111111111111000000000000000000000000010;
		12663: Delta = 39'sb000000000000111111111111111111111111110;
		1170: Delta = 39'sb111111111110111111111111111111111111110;
		11495: Delta = 39'sb000000000010000000000000000000000000010;
		2346: Delta = 39'sb111111111110000000000000000000000000010;
		11491: Delta = 39'sb000000000001111111111111111111111111110;
		2342: Delta = 39'sb111111111101111111111111111111111111110;
		9151: Delta = 39'sb000000000100000000000000000000000000010;
		4690: Delta = 39'sb111111111100000000000000000000000000010;
		9147: Delta = 39'sb000000000011111111111111111111111111110;
		4686: Delta = 39'sb111111111011111111111111111111111111110;
		4463: Delta = 39'sb000000001000000000000000000000000000010;
		9378: Delta = 39'sb111111111000000000000000000000000000010;
		4459: Delta = 39'sb000000000111111111111111111111111111110;
		9374: Delta = 39'sb111111110111111111111111111111111111110;
		8924: Delta = 39'sb000000010000000000000000000000000000010;
		4917: Delta = 39'sb111111110000000000000000000000000000010;
		8920: Delta = 39'sb000000001111111111111111111111111111110;
		4913: Delta = 39'sb111111101111111111111111111111111111110;
		4009: Delta = 39'sb000000100000000000000000000000000000010;
		9832: Delta = 39'sb111111100000000000000000000000000000010;
		4005: Delta = 39'sb000000011111111111111111111111111111110;
		9828: Delta = 39'sb111111011111111111111111111111111111110;
		8016: Delta = 39'sb000001000000000000000000000000000000010;
		5825: Delta = 39'sb111111000000000000000000000000000000010;
		8012: Delta = 39'sb000000111111111111111111111111111111110;
		5821: Delta = 39'sb111110111111111111111111111111111111110;
		2193: Delta = 39'sb000010000000000000000000000000000000010;
		11648: Delta = 39'sb111110000000000000000000000000000000010;
		2189: Delta = 39'sb000001111111111111111111111111111111110;
		11644: Delta = 39'sb111101111111111111111111111111111111110;
		4384: Delta = 39'sb000100000000000000000000000000000000010;
		9457: Delta = 39'sb111100000000000000000000000000000000010;
		4380: Delta = 39'sb000011111111111111111111111111111111110;
		9453: Delta = 39'sb111011111111111111111111111111111111110;
		8766: Delta = 39'sb001000000000000000000000000000000000010;
		5075: Delta = 39'sb111000000000000000000000000000000000010;
		8762: Delta = 39'sb000111111111111111111111111111111111110;
		5071: Delta = 39'sb110111111111111111111111111111111111110;
		3693: Delta = 39'sb010000000000000000000000000000000000010;
		10148: Delta = 39'sb110000000000000000000000000000000000010;
		3689: Delta = 39'sb001111111111111111111111111111111111110;
		10144: Delta = 39'sb101111111111111111111111111111111111110;
		12: Delta = 39'sb000000000000000000000000000000000001100;
		13825: Delta = 39'sb111111111111111111111111111111111110100;
		20: Delta = 39'sb000000000000000000000000000000000010100;
		13817: Delta = 39'sb111111111111111111111111111111111101100;
		36: Delta = 39'sb000000000000000000000000000000000100100;
		13809: Delta = 39'sb111111111111111111111111111111111100100;
		28: Delta = 39'sb000000000000000000000000000000000011100;
		13801: Delta = 39'sb111111111111111111111111111111111011100;
		68: Delta = 39'sb000000000000000000000000000000001000100;
		13777: Delta = 39'sb111111111111111111111111111111111000100;
		60: Delta = 39'sb000000000000000000000000000000000111100;
		13769: Delta = 39'sb111111111111111111111111111111110111100;
		132: Delta = 39'sb000000000000000000000000000000010000100;
		13713: Delta = 39'sb111111111111111111111111111111110000100;
		124: Delta = 39'sb000000000000000000000000000000001111100;
		13705: Delta = 39'sb111111111111111111111111111111101111100;
		260: Delta = 39'sb000000000000000000000000000000100000100;
		13585: Delta = 39'sb111111111111111111111111111111100000100;
		252: Delta = 39'sb000000000000000000000000000000011111100;
		13577: Delta = 39'sb111111111111111111111111111111011111100;
		516: Delta = 39'sb000000000000000000000000000001000000100;
		13329: Delta = 39'sb111111111111111111111111111111000000100;
		508: Delta = 39'sb000000000000000000000000000000111111100;
		13321: Delta = 39'sb111111111111111111111111111110111111100;
		1028: Delta = 39'sb000000000000000000000000000010000000100;
		12817: Delta = 39'sb111111111111111111111111111110000000100;
		1020: Delta = 39'sb000000000000000000000000000001111111100;
		12809: Delta = 39'sb111111111111111111111111111101111111100;
		2052: Delta = 39'sb000000000000000000000000000100000000100;
		11793: Delta = 39'sb111111111111111111111111111100000000100;
		2044: Delta = 39'sb000000000000000000000000000011111111100;
		11785: Delta = 39'sb111111111111111111111111111011111111100;
		4100: Delta = 39'sb000000000000000000000000001000000000100;
		9745: Delta = 39'sb111111111111111111111111111000000000100;
		4092: Delta = 39'sb000000000000000000000000000111111111100;
		9737: Delta = 39'sb111111111111111111111111110111111111100;
		8196: Delta = 39'sb000000000000000000000000010000000000100;
		5649: Delta = 39'sb111111111111111111111111110000000000100;
		8188: Delta = 39'sb000000000000000000000000001111111111100;
		5641: Delta = 39'sb111111111111111111111111101111111111100;
		2551: Delta = 39'sb000000000000000000000000100000000000100;
		11294: Delta = 39'sb111111111111111111111111100000000000100;
		2543: Delta = 39'sb000000000000000000000000011111111111100;
		11286: Delta = 39'sb111111111111111111111111011111111111100;
		5098: Delta = 39'sb000000000000000000000001000000000000100;
		8747: Delta = 39'sb111111111111111111111111000000000000100;
		5090: Delta = 39'sb000000000000000000000000111111111111100;
		8739: Delta = 39'sb111111111111111111111110111111111111100;
		10192: Delta = 39'sb000000000000000000000010000000000000100;
		3653: Delta = 39'sb111111111111111111111110000000000000100;
		10184: Delta = 39'sb000000000000000000000001111111111111100;
		3645: Delta = 39'sb111111111111111111111101111111111111100;
		6543: Delta = 39'sb000000000000000000000100000000000000100;
		7302: Delta = 39'sb111111111111111111111100000000000000100;
		6535: Delta = 39'sb000000000000000000000011111111111111100;
		7294: Delta = 39'sb111111111111111111111011111111111111100;
		13082: Delta = 39'sb000000000000000000001000000000000000100;
		763: Delta = 39'sb111111111111111111111000000000000000100;
		13074: Delta = 39'sb000000000000000000000111111111111111100;
		755: Delta = 39'sb111111111111111111110111111111111111100;
		12323: Delta = 39'sb000000000000000000010000000000000000100;
		1522: Delta = 39'sb111111111111111111110000000000000000100;
		12315: Delta = 39'sb000000000000000000001111111111111111100;
		1514: Delta = 39'sb111111111111111111101111111111111111100;
		10805: Delta = 39'sb000000000000000000100000000000000000100;
		3040: Delta = 39'sb111111111111111111100000000000000000100;
		10797: Delta = 39'sb000000000000000000011111111111111111100;
		3032: Delta = 39'sb111111111111111111011111111111111111100;
		7769: Delta = 39'sb000000000000000001000000000000000000100;
		6076: Delta = 39'sb111111111111111111000000000000000000100;
		7761: Delta = 39'sb000000000000000000111111111111111111100;
		6068: Delta = 39'sb111111111111111110111111111111111111100;
		1697: Delta = 39'sb000000000000000010000000000000000000100;
		12148: Delta = 39'sb111111111111111110000000000000000000100;
		1689: Delta = 39'sb000000000000000001111111111111111111100;
		12140: Delta = 39'sb111111111111111101111111111111111111100;
		3390: Delta = 39'sb000000000000000100000000000000000000100;
		10455: Delta = 39'sb111111111111111100000000000000000000100;
		3382: Delta = 39'sb000000000000000011111111111111111111100;
		10447: Delta = 39'sb111111111111111011111111111111111111100;
		6776: Delta = 39'sb000000000000001000000000000000000000100;
		7069: Delta = 39'sb111111111111111000000000000000000000100;
		6768: Delta = 39'sb000000000000000111111111111111111111100;
		7061: Delta = 39'sb111111111111110111111111111111111111100;
		13548: Delta = 39'sb000000000000010000000000000000000000100;
		297: Delta = 39'sb111111111111110000000000000000000000100;
		13540: Delta = 39'sb000000000000001111111111111111111111100;
		289: Delta = 39'sb111111111111101111111111111111111111100;
		13255: Delta = 39'sb000000000000100000000000000000000000100;
		590: Delta = 39'sb111111111111100000000000000000000000100;
		13247: Delta = 39'sb000000000000011111111111111111111111100;
		582: Delta = 39'sb111111111111011111111111111111111111100;
		12669: Delta = 39'sb000000000001000000000000000000000000100;
		1176: Delta = 39'sb111111111111000000000000000000000000100;
		12661: Delta = 39'sb000000000000111111111111111111111111100;
		1168: Delta = 39'sb111111111110111111111111111111111111100;
		11497: Delta = 39'sb000000000010000000000000000000000000100;
		2348: Delta = 39'sb111111111110000000000000000000000000100;
		11489: Delta = 39'sb000000000001111111111111111111111111100;
		2340: Delta = 39'sb111111111101111111111111111111111111100;
		9153: Delta = 39'sb000000000100000000000000000000000000100;
		4692: Delta = 39'sb111111111100000000000000000000000000100;
		9145: Delta = 39'sb000000000011111111111111111111111111100;
		4684: Delta = 39'sb111111111011111111111111111111111111100;
		4465: Delta = 39'sb000000001000000000000000000000000000100;
		9380: Delta = 39'sb111111111000000000000000000000000000100;
		4457: Delta = 39'sb000000000111111111111111111111111111100;
		9372: Delta = 39'sb111111110111111111111111111111111111100;
		8926: Delta = 39'sb000000010000000000000000000000000000100;
		4919: Delta = 39'sb111111110000000000000000000000000000100;
		8918: Delta = 39'sb000000001111111111111111111111111111100;
		4911: Delta = 39'sb111111101111111111111111111111111111100;
		4011: Delta = 39'sb000000100000000000000000000000000000100;
		9834: Delta = 39'sb111111100000000000000000000000000000100;
		4003: Delta = 39'sb000000011111111111111111111111111111100;
		9826: Delta = 39'sb111111011111111111111111111111111111100;
		8018: Delta = 39'sb000001000000000000000000000000000000100;
		5827: Delta = 39'sb111111000000000000000000000000000000100;
		8010: Delta = 39'sb000000111111111111111111111111111111100;
		5819: Delta = 39'sb111110111111111111111111111111111111100;
		2195: Delta = 39'sb000010000000000000000000000000000000100;
		11650: Delta = 39'sb111110000000000000000000000000000000100;
		2187: Delta = 39'sb000001111111111111111111111111111111100;
		11642: Delta = 39'sb111101111111111111111111111111111111100;
		4386: Delta = 39'sb000100000000000000000000000000000000100;
		9459: Delta = 39'sb111100000000000000000000000000000000100;
		4378: Delta = 39'sb000011111111111111111111111111111111100;
		9451: Delta = 39'sb111011111111111111111111111111111111100;
		8768: Delta = 39'sb001000000000000000000000000000000000100;
		5077: Delta = 39'sb111000000000000000000000000000000000100;
		8760: Delta = 39'sb000111111111111111111111111111111111100;
		5069: Delta = 39'sb110111111111111111111111111111111111100;
		3695: Delta = 39'sb010000000000000000000000000000000000100;
		10150: Delta = 39'sb110000000000000000000000000000000000100;
		3687: Delta = 39'sb001111111111111111111111111111111111100;
		10142: Delta = 39'sb101111111111111111111111111111111111100;
		24: Delta = 39'sb000000000000000000000000000000000011000;
		13813: Delta = 39'sb111111111111111111111111111111111101000;
		40: Delta = 39'sb000000000000000000000000000000000101000;
		13797: Delta = 39'sb111111111111111111111111111111111011000;
		72: Delta = 39'sb000000000000000000000000000000001001000;
		13781: Delta = 39'sb111111111111111111111111111111111001000;
		56: Delta = 39'sb000000000000000000000000000000000111000;
		13765: Delta = 39'sb111111111111111111111111111111110111000;
		136: Delta = 39'sb000000000000000000000000000000010001000;
		13717: Delta = 39'sb111111111111111111111111111111110001000;
		120: Delta = 39'sb000000000000000000000000000000001111000;
		13701: Delta = 39'sb111111111111111111111111111111101111000;
		264: Delta = 39'sb000000000000000000000000000000100001000;
		13589: Delta = 39'sb111111111111111111111111111111100001000;
		248: Delta = 39'sb000000000000000000000000000000011111000;
		13573: Delta = 39'sb111111111111111111111111111111011111000;
		520: Delta = 39'sb000000000000000000000000000001000001000;
		13333: Delta = 39'sb111111111111111111111111111111000001000;
		504: Delta = 39'sb000000000000000000000000000000111111000;
		13317: Delta = 39'sb111111111111111111111111111110111111000;
		1032: Delta = 39'sb000000000000000000000000000010000001000;
		12821: Delta = 39'sb111111111111111111111111111110000001000;
		1016: Delta = 39'sb000000000000000000000000000001111111000;
		12805: Delta = 39'sb111111111111111111111111111101111111000;
		2056: Delta = 39'sb000000000000000000000000000100000001000;
		11797: Delta = 39'sb111111111111111111111111111100000001000;
		2040: Delta = 39'sb000000000000000000000000000011111111000;
		11781: Delta = 39'sb111111111111111111111111111011111111000;
		4104: Delta = 39'sb000000000000000000000000001000000001000;
		9749: Delta = 39'sb111111111111111111111111111000000001000;
		4088: Delta = 39'sb000000000000000000000000000111111111000;
		9733: Delta = 39'sb111111111111111111111111110111111111000;
		8200: Delta = 39'sb000000000000000000000000010000000001000;
		5653: Delta = 39'sb111111111111111111111111110000000001000;
		8184: Delta = 39'sb000000000000000000000000001111111111000;
		5637: Delta = 39'sb111111111111111111111111101111111111000;
		2555: Delta = 39'sb000000000000000000000000100000000001000;
		11298: Delta = 39'sb111111111111111111111111100000000001000;
		2539: Delta = 39'sb000000000000000000000000011111111111000;
		11282: Delta = 39'sb111111111111111111111111011111111111000;
		5102: Delta = 39'sb000000000000000000000001000000000001000;
		8751: Delta = 39'sb111111111111111111111111000000000001000;
		5086: Delta = 39'sb000000000000000000000000111111111111000;
		8735: Delta = 39'sb111111111111111111111110111111111111000;
		10196: Delta = 39'sb000000000000000000000010000000000001000;
		3657: Delta = 39'sb111111111111111111111110000000000001000;
		10180: Delta = 39'sb000000000000000000000001111111111111000;
		3641: Delta = 39'sb111111111111111111111101111111111111000;
		6547: Delta = 39'sb000000000000000000000100000000000001000;
		7306: Delta = 39'sb111111111111111111111100000000000001000;
		6531: Delta = 39'sb000000000000000000000011111111111111000;
		7290: Delta = 39'sb111111111111111111111011111111111111000;
		13086: Delta = 39'sb000000000000000000001000000000000001000;
		767: Delta = 39'sb111111111111111111111000000000000001000;
		13070: Delta = 39'sb000000000000000000000111111111111111000;
		751: Delta = 39'sb111111111111111111110111111111111111000;
		12327: Delta = 39'sb000000000000000000010000000000000001000;
		1526: Delta = 39'sb111111111111111111110000000000000001000;
		12311: Delta = 39'sb000000000000000000001111111111111111000;
		1510: Delta = 39'sb111111111111111111101111111111111111000;
		10809: Delta = 39'sb000000000000000000100000000000000001000;
		3044: Delta = 39'sb111111111111111111100000000000000001000;
		10793: Delta = 39'sb000000000000000000011111111111111111000;
		3028: Delta = 39'sb111111111111111111011111111111111111000;
		7773: Delta = 39'sb000000000000000001000000000000000001000;
		6080: Delta = 39'sb111111111111111111000000000000000001000;
		7757: Delta = 39'sb000000000000000000111111111111111111000;
		6064: Delta = 39'sb111111111111111110111111111111111111000;
		1701: Delta = 39'sb000000000000000010000000000000000001000;
		12152: Delta = 39'sb111111111111111110000000000000000001000;
		1685: Delta = 39'sb000000000000000001111111111111111111000;
		12136: Delta = 39'sb111111111111111101111111111111111111000;
		3394: Delta = 39'sb000000000000000100000000000000000001000;
		10459: Delta = 39'sb111111111111111100000000000000000001000;
		3378: Delta = 39'sb000000000000000011111111111111111111000;
		10443: Delta = 39'sb111111111111111011111111111111111111000;
		6780: Delta = 39'sb000000000000001000000000000000000001000;
		7073: Delta = 39'sb111111111111111000000000000000000001000;
		6764: Delta = 39'sb000000000000000111111111111111111111000;
		7057: Delta = 39'sb111111111111110111111111111111111111000;
		13552: Delta = 39'sb000000000000010000000000000000000001000;
		301: Delta = 39'sb111111111111110000000000000000000001000;
		13536: Delta = 39'sb000000000000001111111111111111111111000;
		285: Delta = 39'sb111111111111101111111111111111111111000;
		13259: Delta = 39'sb000000000000100000000000000000000001000;
		594: Delta = 39'sb111111111111100000000000000000000001000;
		13243: Delta = 39'sb000000000000011111111111111111111111000;
		578: Delta = 39'sb111111111111011111111111111111111111000;
		12673: Delta = 39'sb000000000001000000000000000000000001000;
		1180: Delta = 39'sb111111111111000000000000000000000001000;
		12657: Delta = 39'sb000000000000111111111111111111111111000;
		1164: Delta = 39'sb111111111110111111111111111111111111000;
		11501: Delta = 39'sb000000000010000000000000000000000001000;
		2352: Delta = 39'sb111111111110000000000000000000000001000;
		11485: Delta = 39'sb000000000001111111111111111111111111000;
		2336: Delta = 39'sb111111111101111111111111111111111111000;
		9157: Delta = 39'sb000000000100000000000000000000000001000;
		4696: Delta = 39'sb111111111100000000000000000000000001000;
		9141: Delta = 39'sb000000000011111111111111111111111111000;
		4680: Delta = 39'sb111111111011111111111111111111111111000;
		4469: Delta = 39'sb000000001000000000000000000000000001000;
		9384: Delta = 39'sb111111111000000000000000000000000001000;
		4453: Delta = 39'sb000000000111111111111111111111111111000;
		9368: Delta = 39'sb111111110111111111111111111111111111000;
		8930: Delta = 39'sb000000010000000000000000000000000001000;
		4923: Delta = 39'sb111111110000000000000000000000000001000;
		8914: Delta = 39'sb000000001111111111111111111111111111000;
		4907: Delta = 39'sb111111101111111111111111111111111111000;
		4015: Delta = 39'sb000000100000000000000000000000000001000;
		9838: Delta = 39'sb111111100000000000000000000000000001000;
		3999: Delta = 39'sb000000011111111111111111111111111111000;
		9822: Delta = 39'sb111111011111111111111111111111111111000;
		8022: Delta = 39'sb000001000000000000000000000000000001000;
		5831: Delta = 39'sb111111000000000000000000000000000001000;
		8006: Delta = 39'sb000000111111111111111111111111111111000;
		5815: Delta = 39'sb111110111111111111111111111111111111000;
		2199: Delta = 39'sb000010000000000000000000000000000001000;
		11654: Delta = 39'sb111110000000000000000000000000000001000;
		2183: Delta = 39'sb000001111111111111111111111111111111000;
		11638: Delta = 39'sb111101111111111111111111111111111111000;
		4390: Delta = 39'sb000100000000000000000000000000000001000;
		9463: Delta = 39'sb111100000000000000000000000000000001000;
		4374: Delta = 39'sb000011111111111111111111111111111111000;
		9447: Delta = 39'sb111011111111111111111111111111111111000;
		8772: Delta = 39'sb001000000000000000000000000000000001000;
		5081: Delta = 39'sb111000000000000000000000000000000001000;
		8756: Delta = 39'sb000111111111111111111111111111111111000;
		5065: Delta = 39'sb110111111111111111111111111111111111000;
		3699: Delta = 39'sb010000000000000000000000000000000001000;
		10154: Delta = 39'sb110000000000000000000000000000000001000;
		3683: Delta = 39'sb001111111111111111111111111111111111000;
		10138: Delta = 39'sb101111111111111111111111111111111111000;
		48: Delta = 39'sb000000000000000000000000000000000110000;
		13789: Delta = 39'sb111111111111111111111111111111111010000;
		80: Delta = 39'sb000000000000000000000000000000001010000;
		13757: Delta = 39'sb111111111111111111111111111111110110000;
		144: Delta = 39'sb000000000000000000000000000000010010000;
		13725: Delta = 39'sb111111111111111111111111111111110010000;
		112: Delta = 39'sb000000000000000000000000000000001110000;
		13693: Delta = 39'sb111111111111111111111111111111101110000;
		272: Delta = 39'sb000000000000000000000000000000100010000;
		13597: Delta = 39'sb111111111111111111111111111111100010000;
		240: Delta = 39'sb000000000000000000000000000000011110000;
		13565: Delta = 39'sb111111111111111111111111111111011110000;
		528: Delta = 39'sb000000000000000000000000000001000010000;
		13341: Delta = 39'sb111111111111111111111111111111000010000;
		496: Delta = 39'sb000000000000000000000000000000111110000;
		13309: Delta = 39'sb111111111111111111111111111110111110000;
		1040: Delta = 39'sb000000000000000000000000000010000010000;
		12829: Delta = 39'sb111111111111111111111111111110000010000;
		1008: Delta = 39'sb000000000000000000000000000001111110000;
		12797: Delta = 39'sb111111111111111111111111111101111110000;
		2064: Delta = 39'sb000000000000000000000000000100000010000;
		11805: Delta = 39'sb111111111111111111111111111100000010000;
		2032: Delta = 39'sb000000000000000000000000000011111110000;
		11773: Delta = 39'sb111111111111111111111111111011111110000;
		4112: Delta = 39'sb000000000000000000000000001000000010000;
		9757: Delta = 39'sb111111111111111111111111111000000010000;
		4080: Delta = 39'sb000000000000000000000000000111111110000;
		9725: Delta = 39'sb111111111111111111111111110111111110000;
		8208: Delta = 39'sb000000000000000000000000010000000010000;
		5661: Delta = 39'sb111111111111111111111111110000000010000;
		8176: Delta = 39'sb000000000000000000000000001111111110000;
		5629: Delta = 39'sb111111111111111111111111101111111110000;
		2563: Delta = 39'sb000000000000000000000000100000000010000;
		11306: Delta = 39'sb111111111111111111111111100000000010000;
		2531: Delta = 39'sb000000000000000000000000011111111110000;
		11274: Delta = 39'sb111111111111111111111111011111111110000;
		5110: Delta = 39'sb000000000000000000000001000000000010000;
		8759: Delta = 39'sb111111111111111111111111000000000010000;
		5078: Delta = 39'sb000000000000000000000000111111111110000;
		8727: Delta = 39'sb111111111111111111111110111111111110000;
		10204: Delta = 39'sb000000000000000000000010000000000010000;
		3665: Delta = 39'sb111111111111111111111110000000000010000;
		10172: Delta = 39'sb000000000000000000000001111111111110000;
		3633: Delta = 39'sb111111111111111111111101111111111110000;
		6555: Delta = 39'sb000000000000000000000100000000000010000;
		7314: Delta = 39'sb111111111111111111111100000000000010000;
		6523: Delta = 39'sb000000000000000000000011111111111110000;
		7282: Delta = 39'sb111111111111111111111011111111111110000;
		13094: Delta = 39'sb000000000000000000001000000000000010000;
		775: Delta = 39'sb111111111111111111111000000000000010000;
		13062: Delta = 39'sb000000000000000000000111111111111110000;
		743: Delta = 39'sb111111111111111111110111111111111110000;
		12335: Delta = 39'sb000000000000000000010000000000000010000;
		1534: Delta = 39'sb111111111111111111110000000000000010000;
		12303: Delta = 39'sb000000000000000000001111111111111110000;
		1502: Delta = 39'sb111111111111111111101111111111111110000;
		10817: Delta = 39'sb000000000000000000100000000000000010000;
		3052: Delta = 39'sb111111111111111111100000000000000010000;
		10785: Delta = 39'sb000000000000000000011111111111111110000;
		3020: Delta = 39'sb111111111111111111011111111111111110000;
		7781: Delta = 39'sb000000000000000001000000000000000010000;
		6088: Delta = 39'sb111111111111111111000000000000000010000;
		7749: Delta = 39'sb000000000000000000111111111111111110000;
		6056: Delta = 39'sb111111111111111110111111111111111110000;
		1709: Delta = 39'sb000000000000000010000000000000000010000;
		12160: Delta = 39'sb111111111111111110000000000000000010000;
		1677: Delta = 39'sb000000000000000001111111111111111110000;
		12128: Delta = 39'sb111111111111111101111111111111111110000;
		3402: Delta = 39'sb000000000000000100000000000000000010000;
		10467: Delta = 39'sb111111111111111100000000000000000010000;
		3370: Delta = 39'sb000000000000000011111111111111111110000;
		10435: Delta = 39'sb111111111111111011111111111111111110000;
		6788: Delta = 39'sb000000000000001000000000000000000010000;
		7081: Delta = 39'sb111111111111111000000000000000000010000;
		6756: Delta = 39'sb000000000000000111111111111111111110000;
		7049: Delta = 39'sb111111111111110111111111111111111110000;
		13560: Delta = 39'sb000000000000010000000000000000000010000;
		309: Delta = 39'sb111111111111110000000000000000000010000;
		13528: Delta = 39'sb000000000000001111111111111111111110000;
		277: Delta = 39'sb111111111111101111111111111111111110000;
		13267: Delta = 39'sb000000000000100000000000000000000010000;
		602: Delta = 39'sb111111111111100000000000000000000010000;
		13235: Delta = 39'sb000000000000011111111111111111111110000;
		570: Delta = 39'sb111111111111011111111111111111111110000;
		12681: Delta = 39'sb000000000001000000000000000000000010000;
		1188: Delta = 39'sb111111111111000000000000000000000010000;
		12649: Delta = 39'sb000000000000111111111111111111111110000;
		1156: Delta = 39'sb111111111110111111111111111111111110000;
		11509: Delta = 39'sb000000000010000000000000000000000010000;
		2360: Delta = 39'sb111111111110000000000000000000000010000;
		11477: Delta = 39'sb000000000001111111111111111111111110000;
		2328: Delta = 39'sb111111111101111111111111111111111110000;
		9165: Delta = 39'sb000000000100000000000000000000000010000;
		4704: Delta = 39'sb111111111100000000000000000000000010000;
		9133: Delta = 39'sb000000000011111111111111111111111110000;
		4672: Delta = 39'sb111111111011111111111111111111111110000;
		4477: Delta = 39'sb000000001000000000000000000000000010000;
		9392: Delta = 39'sb111111111000000000000000000000000010000;
		4445: Delta = 39'sb000000000111111111111111111111111110000;
		9360: Delta = 39'sb111111110111111111111111111111111110000;
		8938: Delta = 39'sb000000010000000000000000000000000010000;
		4931: Delta = 39'sb111111110000000000000000000000000010000;
		8906: Delta = 39'sb000000001111111111111111111111111110000;
		4899: Delta = 39'sb111111101111111111111111111111111110000;
		4023: Delta = 39'sb000000100000000000000000000000000010000;
		9846: Delta = 39'sb111111100000000000000000000000000010000;
		3991: Delta = 39'sb000000011111111111111111111111111110000;
		9814: Delta = 39'sb111111011111111111111111111111111110000;
		8030: Delta = 39'sb000001000000000000000000000000000010000;
		5839: Delta = 39'sb111111000000000000000000000000000010000;
		7998: Delta = 39'sb000000111111111111111111111111111110000;
		5807: Delta = 39'sb111110111111111111111111111111111110000;
		2207: Delta = 39'sb000010000000000000000000000000000010000;
		11662: Delta = 39'sb111110000000000000000000000000000010000;
		2175: Delta = 39'sb000001111111111111111111111111111110000;
		11630: Delta = 39'sb111101111111111111111111111111111110000;
		4398: Delta = 39'sb000100000000000000000000000000000010000;
		9471: Delta = 39'sb111100000000000000000000000000000010000;
		4366: Delta = 39'sb000011111111111111111111111111111110000;
		9439: Delta = 39'sb111011111111111111111111111111111110000;
		8780: Delta = 39'sb001000000000000000000000000000000010000;
		5089: Delta = 39'sb111000000000000000000000000000000010000;
		8748: Delta = 39'sb000111111111111111111111111111111110000;
		5057: Delta = 39'sb110111111111111111111111111111111110000;
		3707: Delta = 39'sb010000000000000000000000000000000010000;
		10162: Delta = 39'sb110000000000000000000000000000000010000;
		3675: Delta = 39'sb001111111111111111111111111111111110000;
		10130: Delta = 39'sb101111111111111111111111111111111110000;
		96: Delta = 39'sb000000000000000000000000000000001100000;
		13741: Delta = 39'sb111111111111111111111111111111110100000;
		160: Delta = 39'sb000000000000000000000000000000010100000;
		13677: Delta = 39'sb111111111111111111111111111111101100000;
		288: Delta = 39'sb000000000000000000000000000000100100000;
		13613: Delta = 39'sb111111111111111111111111111111100100000;
		224: Delta = 39'sb000000000000000000000000000000011100000;
		13549: Delta = 39'sb111111111111111111111111111111011100000;
		544: Delta = 39'sb000000000000000000000000000001000100000;
		13357: Delta = 39'sb111111111111111111111111111111000100000;
		480: Delta = 39'sb000000000000000000000000000000111100000;
		13293: Delta = 39'sb111111111111111111111111111110111100000;
		1056: Delta = 39'sb000000000000000000000000000010000100000;
		12845: Delta = 39'sb111111111111111111111111111110000100000;
		992: Delta = 39'sb000000000000000000000000000001111100000;
		12781: Delta = 39'sb111111111111111111111111111101111100000;
		2080: Delta = 39'sb000000000000000000000000000100000100000;
		11821: Delta = 39'sb111111111111111111111111111100000100000;
		2016: Delta = 39'sb000000000000000000000000000011111100000;
		11757: Delta = 39'sb111111111111111111111111111011111100000;
		4128: Delta = 39'sb000000000000000000000000001000000100000;
		9773: Delta = 39'sb111111111111111111111111111000000100000;
		4064: Delta = 39'sb000000000000000000000000000111111100000;
		9709: Delta = 39'sb111111111111111111111111110111111100000;
		8224: Delta = 39'sb000000000000000000000000010000000100000;
		5677: Delta = 39'sb111111111111111111111111110000000100000;
		8160: Delta = 39'sb000000000000000000000000001111111100000;
		5613: Delta = 39'sb111111111111111111111111101111111100000;
		2579: Delta = 39'sb000000000000000000000000100000000100000;
		11322: Delta = 39'sb111111111111111111111111100000000100000;
		2515: Delta = 39'sb000000000000000000000000011111111100000;
		11258: Delta = 39'sb111111111111111111111111011111111100000;
		5126: Delta = 39'sb000000000000000000000001000000000100000;
		8775: Delta = 39'sb111111111111111111111111000000000100000;
		5062: Delta = 39'sb000000000000000000000000111111111100000;
		8711: Delta = 39'sb111111111111111111111110111111111100000;
		10220: Delta = 39'sb000000000000000000000010000000000100000;
		3681: Delta = 39'sb111111111111111111111110000000000100000;
		10156: Delta = 39'sb000000000000000000000001111111111100000;
		3617: Delta = 39'sb111111111111111111111101111111111100000;
		6571: Delta = 39'sb000000000000000000000100000000000100000;
		7330: Delta = 39'sb111111111111111111111100000000000100000;
		6507: Delta = 39'sb000000000000000000000011111111111100000;
		7266: Delta = 39'sb111111111111111111111011111111111100000;
		13110: Delta = 39'sb000000000000000000001000000000000100000;
		791: Delta = 39'sb111111111111111111111000000000000100000;
		13046: Delta = 39'sb000000000000000000000111111111111100000;
		727: Delta = 39'sb111111111111111111110111111111111100000;
		12351: Delta = 39'sb000000000000000000010000000000000100000;
		1550: Delta = 39'sb111111111111111111110000000000000100000;
		12287: Delta = 39'sb000000000000000000001111111111111100000;
		1486: Delta = 39'sb111111111111111111101111111111111100000;
		10833: Delta = 39'sb000000000000000000100000000000000100000;
		3068: Delta = 39'sb111111111111111111100000000000000100000;
		10769: Delta = 39'sb000000000000000000011111111111111100000;
		3004: Delta = 39'sb111111111111111111011111111111111100000;
		7797: Delta = 39'sb000000000000000001000000000000000100000;
		6104: Delta = 39'sb111111111111111111000000000000000100000;
		7733: Delta = 39'sb000000000000000000111111111111111100000;
		6040: Delta = 39'sb111111111111111110111111111111111100000;
		1725: Delta = 39'sb000000000000000010000000000000000100000;
		12176: Delta = 39'sb111111111111111110000000000000000100000;
		1661: Delta = 39'sb000000000000000001111111111111111100000;
		12112: Delta = 39'sb111111111111111101111111111111111100000;
		3418: Delta = 39'sb000000000000000100000000000000000100000;
		10483: Delta = 39'sb111111111111111100000000000000000100000;
		3354: Delta = 39'sb000000000000000011111111111111111100000;
		10419: Delta = 39'sb111111111111111011111111111111111100000;
		6804: Delta = 39'sb000000000000001000000000000000000100000;
		7097: Delta = 39'sb111111111111111000000000000000000100000;
		6740: Delta = 39'sb000000000000000111111111111111111100000;
		7033: Delta = 39'sb111111111111110111111111111111111100000;
		13576: Delta = 39'sb000000000000010000000000000000000100000;
		325: Delta = 39'sb111111111111110000000000000000000100000;
		13512: Delta = 39'sb000000000000001111111111111111111100000;
		261: Delta = 39'sb111111111111101111111111111111111100000;
		13283: Delta = 39'sb000000000000100000000000000000000100000;
		618: Delta = 39'sb111111111111100000000000000000000100000;
		13219: Delta = 39'sb000000000000011111111111111111111100000;
		554: Delta = 39'sb111111111111011111111111111111111100000;
		12697: Delta = 39'sb000000000001000000000000000000000100000;
		1204: Delta = 39'sb111111111111000000000000000000000100000;
		12633: Delta = 39'sb000000000000111111111111111111111100000;
		1140: Delta = 39'sb111111111110111111111111111111111100000;
		11525: Delta = 39'sb000000000010000000000000000000000100000;
		2376: Delta = 39'sb111111111110000000000000000000000100000;
		11461: Delta = 39'sb000000000001111111111111111111111100000;
		2312: Delta = 39'sb111111111101111111111111111111111100000;
		9181: Delta = 39'sb000000000100000000000000000000000100000;
		4720: Delta = 39'sb111111111100000000000000000000000100000;
		9117: Delta = 39'sb000000000011111111111111111111111100000;
		4656: Delta = 39'sb111111111011111111111111111111111100000;
		4493: Delta = 39'sb000000001000000000000000000000000100000;
		9408: Delta = 39'sb111111111000000000000000000000000100000;
		4429: Delta = 39'sb000000000111111111111111111111111100000;
		9344: Delta = 39'sb111111110111111111111111111111111100000;
		8954: Delta = 39'sb000000010000000000000000000000000100000;
		4947: Delta = 39'sb111111110000000000000000000000000100000;
		8890: Delta = 39'sb000000001111111111111111111111111100000;
		4883: Delta = 39'sb111111101111111111111111111111111100000;
		4039: Delta = 39'sb000000100000000000000000000000000100000;
		9862: Delta = 39'sb111111100000000000000000000000000100000;
		3975: Delta = 39'sb000000011111111111111111111111111100000;
		9798: Delta = 39'sb111111011111111111111111111111111100000;
		8046: Delta = 39'sb000001000000000000000000000000000100000;
		5855: Delta = 39'sb111111000000000000000000000000000100000;
		7982: Delta = 39'sb000000111111111111111111111111111100000;
		5791: Delta = 39'sb111110111111111111111111111111111100000;
		2223: Delta = 39'sb000010000000000000000000000000000100000;
		11678: Delta = 39'sb111110000000000000000000000000000100000;
		2159: Delta = 39'sb000001111111111111111111111111111100000;
		11614: Delta = 39'sb111101111111111111111111111111111100000;
		4414: Delta = 39'sb000100000000000000000000000000000100000;
		9487: Delta = 39'sb111100000000000000000000000000000100000;
		4350: Delta = 39'sb000011111111111111111111111111111100000;
		9423: Delta = 39'sb111011111111111111111111111111111100000;
		8796: Delta = 39'sb001000000000000000000000000000000100000;
		5105: Delta = 39'sb111000000000000000000000000000000100000;
		8732: Delta = 39'sb000111111111111111111111111111111100000;
		5041: Delta = 39'sb110111111111111111111111111111111100000;
		3723: Delta = 39'sb010000000000000000000000000000000100000;
		10178: Delta = 39'sb110000000000000000000000000000000100000;
		3659: Delta = 39'sb001111111111111111111111111111111100000;
		10114: Delta = 39'sb101111111111111111111111111111111100000;
		192: Delta = 39'sb000000000000000000000000000000011000000;
		13645: Delta = 39'sb111111111111111111111111111111101000000;
		320: Delta = 39'sb000000000000000000000000000000101000000;
		13517: Delta = 39'sb111111111111111111111111111111011000000;
		576: Delta = 39'sb000000000000000000000000000001001000000;
		13389: Delta = 39'sb111111111111111111111111111111001000000;
		448: Delta = 39'sb000000000000000000000000000000111000000;
		13261: Delta = 39'sb111111111111111111111111111110111000000;
		1088: Delta = 39'sb000000000000000000000000000010001000000;
		12877: Delta = 39'sb111111111111111111111111111110001000000;
		960: Delta = 39'sb000000000000000000000000000001111000000;
		12749: Delta = 39'sb111111111111111111111111111101111000000;
		2112: Delta = 39'sb000000000000000000000000000100001000000;
		11853: Delta = 39'sb111111111111111111111111111100001000000;
		1984: Delta = 39'sb000000000000000000000000000011111000000;
		11725: Delta = 39'sb111111111111111111111111111011111000000;
		4160: Delta = 39'sb000000000000000000000000001000001000000;
		9805: Delta = 39'sb111111111111111111111111111000001000000;
		4032: Delta = 39'sb000000000000000000000000000111111000000;
		9677: Delta = 39'sb111111111111111111111111110111111000000;
		8256: Delta = 39'sb000000000000000000000000010000001000000;
		5709: Delta = 39'sb111111111111111111111111110000001000000;
		8128: Delta = 39'sb000000000000000000000000001111111000000;
		5581: Delta = 39'sb111111111111111111111111101111111000000;
		2611: Delta = 39'sb000000000000000000000000100000001000000;
		11354: Delta = 39'sb111111111111111111111111100000001000000;
		2483: Delta = 39'sb000000000000000000000000011111111000000;
		11226: Delta = 39'sb111111111111111111111111011111111000000;
		5158: Delta = 39'sb000000000000000000000001000000001000000;
		8807: Delta = 39'sb111111111111111111111111000000001000000;
		5030: Delta = 39'sb000000000000000000000000111111111000000;
		8679: Delta = 39'sb111111111111111111111110111111111000000;
		10252: Delta = 39'sb000000000000000000000010000000001000000;
		3713: Delta = 39'sb111111111111111111111110000000001000000;
		10124: Delta = 39'sb000000000000000000000001111111111000000;
		3585: Delta = 39'sb111111111111111111111101111111111000000;
		6603: Delta = 39'sb000000000000000000000100000000001000000;
		7362: Delta = 39'sb111111111111111111111100000000001000000;
		6475: Delta = 39'sb000000000000000000000011111111111000000;
		7234: Delta = 39'sb111111111111111111111011111111111000000;
		13142: Delta = 39'sb000000000000000000001000000000001000000;
		823: Delta = 39'sb111111111111111111111000000000001000000;
		13014: Delta = 39'sb000000000000000000000111111111111000000;
		695: Delta = 39'sb111111111111111111110111111111111000000;
		12383: Delta = 39'sb000000000000000000010000000000001000000;
		1582: Delta = 39'sb111111111111111111110000000000001000000;
		12255: Delta = 39'sb000000000000000000001111111111111000000;
		1454: Delta = 39'sb111111111111111111101111111111111000000;
		10865: Delta = 39'sb000000000000000000100000000000001000000;
		3100: Delta = 39'sb111111111111111111100000000000001000000;
		10737: Delta = 39'sb000000000000000000011111111111111000000;
		2972: Delta = 39'sb111111111111111111011111111111111000000;
		7829: Delta = 39'sb000000000000000001000000000000001000000;
		6136: Delta = 39'sb111111111111111111000000000000001000000;
		7701: Delta = 39'sb000000000000000000111111111111111000000;
		6008: Delta = 39'sb111111111111111110111111111111111000000;
		1757: Delta = 39'sb000000000000000010000000000000001000000;
		12208: Delta = 39'sb111111111111111110000000000000001000000;
		1629: Delta = 39'sb000000000000000001111111111111111000000;
		12080: Delta = 39'sb111111111111111101111111111111111000000;
		3450: Delta = 39'sb000000000000000100000000000000001000000;
		10515: Delta = 39'sb111111111111111100000000000000001000000;
		3322: Delta = 39'sb000000000000000011111111111111111000000;
		10387: Delta = 39'sb111111111111111011111111111111111000000;
		6836: Delta = 39'sb000000000000001000000000000000001000000;
		7129: Delta = 39'sb111111111111111000000000000000001000000;
		6708: Delta = 39'sb000000000000000111111111111111111000000;
		7001: Delta = 39'sb111111111111110111111111111111111000000;
		13608: Delta = 39'sb000000000000010000000000000000001000000;
		357: Delta = 39'sb111111111111110000000000000000001000000;
		13480: Delta = 39'sb000000000000001111111111111111111000000;
		229: Delta = 39'sb111111111111101111111111111111111000000;
		13315: Delta = 39'sb000000000000100000000000000000001000000;
		650: Delta = 39'sb111111111111100000000000000000001000000;
		13187: Delta = 39'sb000000000000011111111111111111111000000;
		522: Delta = 39'sb111111111111011111111111111111111000000;
		12729: Delta = 39'sb000000000001000000000000000000001000000;
		1236: Delta = 39'sb111111111111000000000000000000001000000;
		12601: Delta = 39'sb000000000000111111111111111111111000000;
		1108: Delta = 39'sb111111111110111111111111111111111000000;
		11557: Delta = 39'sb000000000010000000000000000000001000000;
		2408: Delta = 39'sb111111111110000000000000000000001000000;
		11429: Delta = 39'sb000000000001111111111111111111111000000;
		2280: Delta = 39'sb111111111101111111111111111111111000000;
		9213: Delta = 39'sb000000000100000000000000000000001000000;
		4752: Delta = 39'sb111111111100000000000000000000001000000;
		9085: Delta = 39'sb000000000011111111111111111111111000000;
		4624: Delta = 39'sb111111111011111111111111111111111000000;
		4525: Delta = 39'sb000000001000000000000000000000001000000;
		9440: Delta = 39'sb111111111000000000000000000000001000000;
		4397: Delta = 39'sb000000000111111111111111111111111000000;
		9312: Delta = 39'sb111111110111111111111111111111111000000;
		8986: Delta = 39'sb000000010000000000000000000000001000000;
		4979: Delta = 39'sb111111110000000000000000000000001000000;
		8858: Delta = 39'sb000000001111111111111111111111111000000;
		4851: Delta = 39'sb111111101111111111111111111111111000000;
		4071: Delta = 39'sb000000100000000000000000000000001000000;
		9894: Delta = 39'sb111111100000000000000000000000001000000;
		3943: Delta = 39'sb000000011111111111111111111111111000000;
		9766: Delta = 39'sb111111011111111111111111111111111000000;
		8078: Delta = 39'sb000001000000000000000000000000001000000;
		5887: Delta = 39'sb111111000000000000000000000000001000000;
		7950: Delta = 39'sb000000111111111111111111111111111000000;
		5759: Delta = 39'sb111110111111111111111111111111111000000;
		2255: Delta = 39'sb000010000000000000000000000000001000000;
		11710: Delta = 39'sb111110000000000000000000000000001000000;
		2127: Delta = 39'sb000001111111111111111111111111111000000;
		11582: Delta = 39'sb111101111111111111111111111111111000000;
		4446: Delta = 39'sb000100000000000000000000000000001000000;
		9519: Delta = 39'sb111100000000000000000000000000001000000;
		4318: Delta = 39'sb000011111111111111111111111111111000000;
		9391: Delta = 39'sb111011111111111111111111111111111000000;
		8828: Delta = 39'sb001000000000000000000000000000001000000;
		5137: Delta = 39'sb111000000000000000000000000000001000000;
		8700: Delta = 39'sb000111111111111111111111111111111000000;
		5009: Delta = 39'sb110111111111111111111111111111111000000;
		3755: Delta = 39'sb010000000000000000000000000000001000000;
		10210: Delta = 39'sb110000000000000000000000000000001000000;
		3627: Delta = 39'sb001111111111111111111111111111111000000;
		10082: Delta = 39'sb101111111111111111111111111111111000000;
		384: Delta = 39'sb000000000000000000000000000000110000000;
		13453: Delta = 39'sb111111111111111111111111111111010000000;
		640: Delta = 39'sb000000000000000000000000000001010000000;
		13197: Delta = 39'sb111111111111111111111111111110110000000;
		1152: Delta = 39'sb000000000000000000000000000010010000000;
		12941: Delta = 39'sb111111111111111111111111111110010000000;
		896: Delta = 39'sb000000000000000000000000000001110000000;
		12685: Delta = 39'sb111111111111111111111111111101110000000;
		2176: Delta = 39'sb000000000000000000000000000100010000000;
		11917: Delta = 39'sb111111111111111111111111111100010000000;
		1920: Delta = 39'sb000000000000000000000000000011110000000;
		11661: Delta = 39'sb111111111111111111111111111011110000000;
		4224: Delta = 39'sb000000000000000000000000001000010000000;
		9869: Delta = 39'sb111111111111111111111111111000010000000;
		3968: Delta = 39'sb000000000000000000000000000111110000000;
		9613: Delta = 39'sb111111111111111111111111110111110000000;
		8320: Delta = 39'sb000000000000000000000000010000010000000;
		5773: Delta = 39'sb111111111111111111111111110000010000000;
		8064: Delta = 39'sb000000000000000000000000001111110000000;
		5517: Delta = 39'sb111111111111111111111111101111110000000;
		2675: Delta = 39'sb000000000000000000000000100000010000000;
		11418: Delta = 39'sb111111111111111111111111100000010000000;
		2419: Delta = 39'sb000000000000000000000000011111110000000;
		11162: Delta = 39'sb111111111111111111111111011111110000000;
		5222: Delta = 39'sb000000000000000000000001000000010000000;
		8871: Delta = 39'sb111111111111111111111111000000010000000;
		4966: Delta = 39'sb000000000000000000000000111111110000000;
		8615: Delta = 39'sb111111111111111111111110111111110000000;
		10316: Delta = 39'sb000000000000000000000010000000010000000;
		3777: Delta = 39'sb111111111111111111111110000000010000000;
		10060: Delta = 39'sb000000000000000000000001111111110000000;
		3521: Delta = 39'sb111111111111111111111101111111110000000;
		6667: Delta = 39'sb000000000000000000000100000000010000000;
		7426: Delta = 39'sb111111111111111111111100000000010000000;
		6411: Delta = 39'sb000000000000000000000011111111110000000;
		7170: Delta = 39'sb111111111111111111111011111111110000000;
		13206: Delta = 39'sb000000000000000000001000000000010000000;
		887: Delta = 39'sb111111111111111111111000000000010000000;
		12950: Delta = 39'sb000000000000000000000111111111110000000;
		631: Delta = 39'sb111111111111111111110111111111110000000;
		12447: Delta = 39'sb000000000000000000010000000000010000000;
		1646: Delta = 39'sb111111111111111111110000000000010000000;
		12191: Delta = 39'sb000000000000000000001111111111110000000;
		1390: Delta = 39'sb111111111111111111101111111111110000000;
		10929: Delta = 39'sb000000000000000000100000000000010000000;
		3164: Delta = 39'sb111111111111111111100000000000010000000;
		10673: Delta = 39'sb000000000000000000011111111111110000000;
		2908: Delta = 39'sb111111111111111111011111111111110000000;
		7893: Delta = 39'sb000000000000000001000000000000010000000;
		6200: Delta = 39'sb111111111111111111000000000000010000000;
		7637: Delta = 39'sb000000000000000000111111111111110000000;
		5944: Delta = 39'sb111111111111111110111111111111110000000;
		1821: Delta = 39'sb000000000000000010000000000000010000000;
		12272: Delta = 39'sb111111111111111110000000000000010000000;
		1565: Delta = 39'sb000000000000000001111111111111110000000;
		12016: Delta = 39'sb111111111111111101111111111111110000000;
		3514: Delta = 39'sb000000000000000100000000000000010000000;
		10579: Delta = 39'sb111111111111111100000000000000010000000;
		3258: Delta = 39'sb000000000000000011111111111111110000000;
		10323: Delta = 39'sb111111111111111011111111111111110000000;
		6900: Delta = 39'sb000000000000001000000000000000010000000;
		7193: Delta = 39'sb111111111111111000000000000000010000000;
		6644: Delta = 39'sb000000000000000111111111111111110000000;
		6937: Delta = 39'sb111111111111110111111111111111110000000;
		13672: Delta = 39'sb000000000000010000000000000000010000000;
		421: Delta = 39'sb111111111111110000000000000000010000000;
		13416: Delta = 39'sb000000000000001111111111111111110000000;
		165: Delta = 39'sb111111111111101111111111111111110000000;
		13379: Delta = 39'sb000000000000100000000000000000010000000;
		714: Delta = 39'sb111111111111100000000000000000010000000;
		13123: Delta = 39'sb000000000000011111111111111111110000000;
		458: Delta = 39'sb111111111111011111111111111111110000000;
		12793: Delta = 39'sb000000000001000000000000000000010000000;
		1300: Delta = 39'sb111111111111000000000000000000010000000;
		12537: Delta = 39'sb000000000000111111111111111111110000000;
		1044: Delta = 39'sb111111111110111111111111111111110000000;
		11621: Delta = 39'sb000000000010000000000000000000010000000;
		2472: Delta = 39'sb111111111110000000000000000000010000000;
		11365: Delta = 39'sb000000000001111111111111111111110000000;
		2216: Delta = 39'sb111111111101111111111111111111110000000;
		9277: Delta = 39'sb000000000100000000000000000000010000000;
		4816: Delta = 39'sb111111111100000000000000000000010000000;
		9021: Delta = 39'sb000000000011111111111111111111110000000;
		4560: Delta = 39'sb111111111011111111111111111111110000000;
		4589: Delta = 39'sb000000001000000000000000000000010000000;
		9504: Delta = 39'sb111111111000000000000000000000010000000;
		4333: Delta = 39'sb000000000111111111111111111111110000000;
		9248: Delta = 39'sb111111110111111111111111111111110000000;
		9050: Delta = 39'sb000000010000000000000000000000010000000;
		5043: Delta = 39'sb111111110000000000000000000000010000000;
		8794: Delta = 39'sb000000001111111111111111111111110000000;
		4787: Delta = 39'sb111111101111111111111111111111110000000;
		4135: Delta = 39'sb000000100000000000000000000000010000000;
		9958: Delta = 39'sb111111100000000000000000000000010000000;
		3879: Delta = 39'sb000000011111111111111111111111110000000;
		9702: Delta = 39'sb111111011111111111111111111111110000000;
		8142: Delta = 39'sb000001000000000000000000000000010000000;
		5951: Delta = 39'sb111111000000000000000000000000010000000;
		7886: Delta = 39'sb000000111111111111111111111111110000000;
		5695: Delta = 39'sb111110111111111111111111111111110000000;
		2319: Delta = 39'sb000010000000000000000000000000010000000;
		11774: Delta = 39'sb111110000000000000000000000000010000000;
		2063: Delta = 39'sb000001111111111111111111111111110000000;
		11518: Delta = 39'sb111101111111111111111111111111110000000;
		4510: Delta = 39'sb000100000000000000000000000000010000000;
		9583: Delta = 39'sb111100000000000000000000000000010000000;
		4254: Delta = 39'sb000011111111111111111111111111110000000;
		9327: Delta = 39'sb111011111111111111111111111111110000000;
		8892: Delta = 39'sb001000000000000000000000000000010000000;
		5201: Delta = 39'sb111000000000000000000000000000010000000;
		8636: Delta = 39'sb000111111111111111111111111111110000000;
		4945: Delta = 39'sb110111111111111111111111111111110000000;
		3819: Delta = 39'sb010000000000000000000000000000010000000;
		10274: Delta = 39'sb110000000000000000000000000000010000000;
		3563: Delta = 39'sb001111111111111111111111111111110000000;
		10018: Delta = 39'sb101111111111111111111111111111110000000;
		768: Delta = 39'sb000000000000000000000000000001100000000;
		13069: Delta = 39'sb111111111111111111111111111110100000000;
		1280: Delta = 39'sb000000000000000000000000000010100000000;
		12557: Delta = 39'sb111111111111111111111111111101100000000;
		2304: Delta = 39'sb000000000000000000000000000100100000000;
		12045: Delta = 39'sb111111111111111111111111111100100000000;
		1792: Delta = 39'sb000000000000000000000000000011100000000;
		11533: Delta = 39'sb111111111111111111111111111011100000000;
		4352: Delta = 39'sb000000000000000000000000001000100000000;
		9997: Delta = 39'sb111111111111111111111111111000100000000;
		3840: Delta = 39'sb000000000000000000000000000111100000000;
		9485: Delta = 39'sb111111111111111111111111110111100000000;
		8448: Delta = 39'sb000000000000000000000000010000100000000;
		5901: Delta = 39'sb111111111111111111111111110000100000000;
		7936: Delta = 39'sb000000000000000000000000001111100000000;
		5389: Delta = 39'sb111111111111111111111111101111100000000;
		2803: Delta = 39'sb000000000000000000000000100000100000000;
		11546: Delta = 39'sb111111111111111111111111100000100000000;
		2291: Delta = 39'sb000000000000000000000000011111100000000;
		11034: Delta = 39'sb111111111111111111111111011111100000000;
		5350: Delta = 39'sb000000000000000000000001000000100000000;
		8999: Delta = 39'sb111111111111111111111111000000100000000;
		4838: Delta = 39'sb000000000000000000000000111111100000000;
		8487: Delta = 39'sb111111111111111111111110111111100000000;
		10444: Delta = 39'sb000000000000000000000010000000100000000;
		3905: Delta = 39'sb111111111111111111111110000000100000000;
		9932: Delta = 39'sb000000000000000000000001111111100000000;
		3393: Delta = 39'sb111111111111111111111101111111100000000;
		6795: Delta = 39'sb000000000000000000000100000000100000000;
		7554: Delta = 39'sb111111111111111111111100000000100000000;
		6283: Delta = 39'sb000000000000000000000011111111100000000;
		7042: Delta = 39'sb111111111111111111111011111111100000000;
		13334: Delta = 39'sb000000000000000000001000000000100000000;
		1015: Delta = 39'sb111111111111111111111000000000100000000;
		12822: Delta = 39'sb000000000000000000000111111111100000000;
		503: Delta = 39'sb111111111111111111110111111111100000000;
		12575: Delta = 39'sb000000000000000000010000000000100000000;
		1774: Delta = 39'sb111111111111111111110000000000100000000;
		12063: Delta = 39'sb000000000000000000001111111111100000000;
		1262: Delta = 39'sb111111111111111111101111111111100000000;
		11057: Delta = 39'sb000000000000000000100000000000100000000;
		3292: Delta = 39'sb111111111111111111100000000000100000000;
		10545: Delta = 39'sb000000000000000000011111111111100000000;
		2780: Delta = 39'sb111111111111111111011111111111100000000;
		8021: Delta = 39'sb000000000000000001000000000000100000000;
		6328: Delta = 39'sb111111111111111111000000000000100000000;
		7509: Delta = 39'sb000000000000000000111111111111100000000;
		5816: Delta = 39'sb111111111111111110111111111111100000000;
		1949: Delta = 39'sb000000000000000010000000000000100000000;
		12400: Delta = 39'sb111111111111111110000000000000100000000;
		1437: Delta = 39'sb000000000000000001111111111111100000000;
		11888: Delta = 39'sb111111111111111101111111111111100000000;
		3642: Delta = 39'sb000000000000000100000000000000100000000;
		10707: Delta = 39'sb111111111111111100000000000000100000000;
		3130: Delta = 39'sb000000000000000011111111111111100000000;
		10195: Delta = 39'sb111111111111111011111111111111100000000;
		7028: Delta = 39'sb000000000000001000000000000000100000000;
		7321: Delta = 39'sb111111111111111000000000000000100000000;
		6516: Delta = 39'sb000000000000000111111111111111100000000;
		6809: Delta = 39'sb111111111111110111111111111111100000000;
		13800: Delta = 39'sb000000000000010000000000000000100000000;
		549: Delta = 39'sb111111111111110000000000000000100000000;
		13288: Delta = 39'sb000000000000001111111111111111100000000;
		37: Delta = 39'sb111111111111101111111111111111100000000;
		13507: Delta = 39'sb000000000000100000000000000000100000000;
		842: Delta = 39'sb111111111111100000000000000000100000000;
		12995: Delta = 39'sb000000000000011111111111111111100000000;
		330: Delta = 39'sb111111111111011111111111111111100000000;
		12921: Delta = 39'sb000000000001000000000000000000100000000;
		1428: Delta = 39'sb111111111111000000000000000000100000000;
		12409: Delta = 39'sb000000000000111111111111111111100000000;
		916: Delta = 39'sb111111111110111111111111111111100000000;
		11749: Delta = 39'sb000000000010000000000000000000100000000;
		2600: Delta = 39'sb111111111110000000000000000000100000000;
		11237: Delta = 39'sb000000000001111111111111111111100000000;
		2088: Delta = 39'sb111111111101111111111111111111100000000;
		9405: Delta = 39'sb000000000100000000000000000000100000000;
		4944: Delta = 39'sb111111111100000000000000000000100000000;
		8893: Delta = 39'sb000000000011111111111111111111100000000;
		4432: Delta = 39'sb111111111011111111111111111111100000000;
		4717: Delta = 39'sb000000001000000000000000000000100000000;
		9632: Delta = 39'sb111111111000000000000000000000100000000;
		4205: Delta = 39'sb000000000111111111111111111111100000000;
		9120: Delta = 39'sb111111110111111111111111111111100000000;
		9178: Delta = 39'sb000000010000000000000000000000100000000;
		5171: Delta = 39'sb111111110000000000000000000000100000000;
		8666: Delta = 39'sb000000001111111111111111111111100000000;
		4659: Delta = 39'sb111111101111111111111111111111100000000;
		4263: Delta = 39'sb000000100000000000000000000000100000000;
		10086: Delta = 39'sb111111100000000000000000000000100000000;
		3751: Delta = 39'sb000000011111111111111111111111100000000;
		9574: Delta = 39'sb111111011111111111111111111111100000000;
		8270: Delta = 39'sb000001000000000000000000000000100000000;
		6079: Delta = 39'sb111111000000000000000000000000100000000;
		7758: Delta = 39'sb000000111111111111111111111111100000000;
		5567: Delta = 39'sb111110111111111111111111111111100000000;
		2447: Delta = 39'sb000010000000000000000000000000100000000;
		11902: Delta = 39'sb111110000000000000000000000000100000000;
		1935: Delta = 39'sb000001111111111111111111111111100000000;
		11390: Delta = 39'sb111101111111111111111111111111100000000;
		4638: Delta = 39'sb000100000000000000000000000000100000000;
		9711: Delta = 39'sb111100000000000000000000000000100000000;
		4126: Delta = 39'sb000011111111111111111111111111100000000;
		9199: Delta = 39'sb111011111111111111111111111111100000000;
		9020: Delta = 39'sb001000000000000000000000000000100000000;
		5329: Delta = 39'sb111000000000000000000000000000100000000;
		8508: Delta = 39'sb000111111111111111111111111111100000000;
		4817: Delta = 39'sb110111111111111111111111111111100000000;
		3947: Delta = 39'sb010000000000000000000000000000100000000;
		10402: Delta = 39'sb110000000000000000000000000000100000000;
		3435: Delta = 39'sb001111111111111111111111111111100000000;
		9890: Delta = 39'sb101111111111111111111111111111100000000;
		1536: Delta = 39'sb000000000000000000000000000011000000000;
		12301: Delta = 39'sb111111111111111111111111111101000000000;
		2560: Delta = 39'sb000000000000000000000000000101000000000;
		11277: Delta = 39'sb111111111111111111111111111011000000000;
		4608: Delta = 39'sb000000000000000000000000001001000000000;
		10253: Delta = 39'sb111111111111111111111111111001000000000;
		3584: Delta = 39'sb000000000000000000000000000111000000000;
		9229: Delta = 39'sb111111111111111111111111110111000000000;
		8704: Delta = 39'sb000000000000000000000000010001000000000;
		6157: Delta = 39'sb111111111111111111111111110001000000000;
		7680: Delta = 39'sb000000000000000000000000001111000000000;
		5133: Delta = 39'sb111111111111111111111111101111000000000;
		3059: Delta = 39'sb000000000000000000000000100001000000000;
		11802: Delta = 39'sb111111111111111111111111100001000000000;
		2035: Delta = 39'sb000000000000000000000000011111000000000;
		10778: Delta = 39'sb111111111111111111111111011111000000000;
		5606: Delta = 39'sb000000000000000000000001000001000000000;
		9255: Delta = 39'sb111111111111111111111111000001000000000;
		4582: Delta = 39'sb000000000000000000000000111111000000000;
		8231: Delta = 39'sb111111111111111111111110111111000000000;
		10700: Delta = 39'sb000000000000000000000010000001000000000;
		4161: Delta = 39'sb111111111111111111111110000001000000000;
		9676: Delta = 39'sb000000000000000000000001111111000000000;
		3137: Delta = 39'sb111111111111111111111101111111000000000;
		7051: Delta = 39'sb000000000000000000000100000001000000000;
		7810: Delta = 39'sb111111111111111111111100000001000000000;
		6027: Delta = 39'sb000000000000000000000011111111000000000;
		6786: Delta = 39'sb111111111111111111111011111111000000000;
		13590: Delta = 39'sb000000000000000000001000000001000000000;
		1271: Delta = 39'sb111111111111111111111000000001000000000;
		12566: Delta = 39'sb000000000000000000000111111111000000000;
		247: Delta = 39'sb111111111111111111110111111111000000000;
		12831: Delta = 39'sb000000000000000000010000000001000000000;
		2030: Delta = 39'sb111111111111111111110000000001000000000;
		11807: Delta = 39'sb000000000000000000001111111111000000000;
		1006: Delta = 39'sb111111111111111111101111111111000000000;
		11313: Delta = 39'sb000000000000000000100000000001000000000;
		3548: Delta = 39'sb111111111111111111100000000001000000000;
		10289: Delta = 39'sb000000000000000000011111111111000000000;
		2524: Delta = 39'sb111111111111111111011111111111000000000;
		8277: Delta = 39'sb000000000000000001000000000001000000000;
		6584: Delta = 39'sb111111111111111111000000000001000000000;
		7253: Delta = 39'sb000000000000000000111111111111000000000;
		5560: Delta = 39'sb111111111111111110111111111111000000000;
		2205: Delta = 39'sb000000000000000010000000000001000000000;
		12656: Delta = 39'sb111111111111111110000000000001000000000;
		1181: Delta = 39'sb000000000000000001111111111111000000000;
		11632: Delta = 39'sb111111111111111101111111111111000000000;
		3898: Delta = 39'sb000000000000000100000000000001000000000;
		10963: Delta = 39'sb111111111111111100000000000001000000000;
		2874: Delta = 39'sb000000000000000011111111111111000000000;
		9939: Delta = 39'sb111111111111111011111111111111000000000;
		7284: Delta = 39'sb000000000000001000000000000001000000000;
		7577: Delta = 39'sb111111111111111000000000000001000000000;
		6260: Delta = 39'sb000000000000000111111111111111000000000;
		6553: Delta = 39'sb111111111111110111111111111111000000000;
		219: Delta = 39'sb000000000000010000000000000001000000000;
		805: Delta = 39'sb111111111111110000000000000001000000000;
		13032: Delta = 39'sb000000000000001111111111111111000000000;
		13618: Delta = 39'sb111111111111101111111111111111000000000;
		13763: Delta = 39'sb000000000000100000000000000001000000000;
		1098: Delta = 39'sb111111111111100000000000000001000000000;
		12739: Delta = 39'sb000000000000011111111111111111000000000;
		74: Delta = 39'sb111111111111011111111111111111000000000;
		13177: Delta = 39'sb000000000001000000000000000001000000000;
		1684: Delta = 39'sb111111111111000000000000000001000000000;
		12153: Delta = 39'sb000000000000111111111111111111000000000;
		660: Delta = 39'sb111111111110111111111111111111000000000;
		12005: Delta = 39'sb000000000010000000000000000001000000000;
		2856: Delta = 39'sb111111111110000000000000000001000000000;
		10981: Delta = 39'sb000000000001111111111111111111000000000;
		1832: Delta = 39'sb111111111101111111111111111111000000000;
		9661: Delta = 39'sb000000000100000000000000000001000000000;
		5200: Delta = 39'sb111111111100000000000000000001000000000;
		8637: Delta = 39'sb000000000011111111111111111111000000000;
		4176: Delta = 39'sb111111111011111111111111111111000000000;
		4973: Delta = 39'sb000000001000000000000000000001000000000;
		9888: Delta = 39'sb111111111000000000000000000001000000000;
		3949: Delta = 39'sb000000000111111111111111111111000000000;
		8864: Delta = 39'sb111111110111111111111111111111000000000;
		9434: Delta = 39'sb000000010000000000000000000001000000000;
		5427: Delta = 39'sb111111110000000000000000000001000000000;
		8410: Delta = 39'sb000000001111111111111111111111000000000;
		4403: Delta = 39'sb111111101111111111111111111111000000000;
		4519: Delta = 39'sb000000100000000000000000000001000000000;
		10342: Delta = 39'sb111111100000000000000000000001000000000;
		3495: Delta = 39'sb000000011111111111111111111111000000000;
		9318: Delta = 39'sb111111011111111111111111111111000000000;
		8526: Delta = 39'sb000001000000000000000000000001000000000;
		6335: Delta = 39'sb111111000000000000000000000001000000000;
		7502: Delta = 39'sb000000111111111111111111111111000000000;
		5311: Delta = 39'sb111110111111111111111111111111000000000;
		2703: Delta = 39'sb000010000000000000000000000001000000000;
		12158: Delta = 39'sb111110000000000000000000000001000000000;
		1679: Delta = 39'sb000001111111111111111111111111000000000;
		11134: Delta = 39'sb111101111111111111111111111111000000000;
		4894: Delta = 39'sb000100000000000000000000000001000000000;
		9967: Delta = 39'sb111100000000000000000000000001000000000;
		3870: Delta = 39'sb000011111111111111111111111111000000000;
		8943: Delta = 39'sb111011111111111111111111111111000000000;
		9276: Delta = 39'sb001000000000000000000000000001000000000;
		5585: Delta = 39'sb111000000000000000000000000001000000000;
		8252: Delta = 39'sb000111111111111111111111111111000000000;
		4561: Delta = 39'sb110111111111111111111111111111000000000;
		4203: Delta = 39'sb010000000000000000000000000001000000000;
		10658: Delta = 39'sb110000000000000000000000000001000000000;
		3179: Delta = 39'sb001111111111111111111111111111000000000;
		9634: Delta = 39'sb101111111111111111111111111111000000000;
		3072: Delta = 39'sb000000000000000000000000000110000000000;
		10765: Delta = 39'sb111111111111111111111111111010000000000;
		5120: Delta = 39'sb000000000000000000000000001010000000000;
		8717: Delta = 39'sb111111111111111111111111110110000000000;
		9216: Delta = 39'sb000000000000000000000000010010000000000;
		6669: Delta = 39'sb111111111111111111111111110010000000000;
		7168: Delta = 39'sb000000000000000000000000001110000000000;
		4621: Delta = 39'sb111111111111111111111111101110000000000;
		3571: Delta = 39'sb000000000000000000000000100010000000000;
		12314: Delta = 39'sb111111111111111111111111100010000000000;
		1523: Delta = 39'sb000000000000000000000000011110000000000;
		10266: Delta = 39'sb111111111111111111111111011110000000000;
		6118: Delta = 39'sb000000000000000000000001000010000000000;
		9767: Delta = 39'sb111111111111111111111111000010000000000;
		4070: Delta = 39'sb000000000000000000000000111110000000000;
		7719: Delta = 39'sb111111111111111111111110111110000000000;
		11212: Delta = 39'sb000000000000000000000010000010000000000;
		4673: Delta = 39'sb111111111111111111111110000010000000000;
		9164: Delta = 39'sb000000000000000000000001111110000000000;
		2625: Delta = 39'sb111111111111111111111101111110000000000;
		7563: Delta = 39'sb000000000000000000000100000010000000000;
		8322: Delta = 39'sb111111111111111111111100000010000000000;
		5515: Delta = 39'sb000000000000000000000011111110000000000;
		6274: Delta = 39'sb111111111111111111111011111110000000000;
		265: Delta = 39'sb000000000000000000001000000010000000000;
		1783: Delta = 39'sb111111111111111111111000000010000000000;
		12054: Delta = 39'sb000000000000000000000111111110000000000;
		13572: Delta = 39'sb111111111111111111110111111110000000000;
		13343: Delta = 39'sb000000000000000000010000000010000000000;
		2542: Delta = 39'sb111111111111111111110000000010000000000;
		11295: Delta = 39'sb000000000000000000001111111110000000000;
		494: Delta = 39'sb111111111111111111101111111110000000000;
		11825: Delta = 39'sb000000000000000000100000000010000000000;
		4060: Delta = 39'sb111111111111111111100000000010000000000;
		9777: Delta = 39'sb000000000000000000011111111110000000000;
		2012: Delta = 39'sb111111111111111111011111111110000000000;
		8789: Delta = 39'sb000000000000000001000000000010000000000;
		7096: Delta = 39'sb111111111111111111000000000010000000000;
		6741: Delta = 39'sb000000000000000000111111111110000000000;
		5048: Delta = 39'sb111111111111111110111111111110000000000;
		2717: Delta = 39'sb000000000000000010000000000010000000000;
		13168: Delta = 39'sb111111111111111110000000000010000000000;
		669: Delta = 39'sb000000000000000001111111111110000000000;
		11120: Delta = 39'sb111111111111111101111111111110000000000;
		4410: Delta = 39'sb000000000000000100000000000010000000000;
		11475: Delta = 39'sb111111111111111100000000000010000000000;
		2362: Delta = 39'sb000000000000000011111111111110000000000;
		9427: Delta = 39'sb111111111111111011111111111110000000000;
		7796: Delta = 39'sb000000000000001000000000000010000000000;
		8089: Delta = 39'sb111111111111111000000000000010000000000;
		5748: Delta = 39'sb000000000000000111111111111110000000000;
		6041: Delta = 39'sb111111111111110111111111111110000000000;
		731: Delta = 39'sb000000000000010000000000000010000000000;
		1317: Delta = 39'sb111111111111110000000000000010000000000;
		12520: Delta = 39'sb000000000000001111111111111110000000000;
		13106: Delta = 39'sb111111111111101111111111111110000000000;
		438: Delta = 39'sb000000000000100000000000000010000000000;
		1610: Delta = 39'sb111111111111100000000000000010000000000;
		12227: Delta = 39'sb000000000000011111111111111110000000000;
		13399: Delta = 39'sb111111111111011111111111111110000000000;
		13689: Delta = 39'sb000000000001000000000000000010000000000;
		2196: Delta = 39'sb111111111111000000000000000010000000000;
		11641: Delta = 39'sb000000000000111111111111111110000000000;
		148: Delta = 39'sb111111111110111111111111111110000000000;
		12517: Delta = 39'sb000000000010000000000000000010000000000;
		3368: Delta = 39'sb111111111110000000000000000010000000000;
		10469: Delta = 39'sb000000000001111111111111111110000000000;
		1320: Delta = 39'sb111111111101111111111111111110000000000;
		10173: Delta = 39'sb000000000100000000000000000010000000000;
		5712: Delta = 39'sb111111111100000000000000000010000000000;
		8125: Delta = 39'sb000000000011111111111111111110000000000;
		3664: Delta = 39'sb111111111011111111111111111110000000000;
		5485: Delta = 39'sb000000001000000000000000000010000000000;
		10400: Delta = 39'sb111111111000000000000000000010000000000;
		3437: Delta = 39'sb000000000111111111111111111110000000000;
		8352: Delta = 39'sb111111110111111111111111111110000000000;
		9946: Delta = 39'sb000000010000000000000000000010000000000;
		5939: Delta = 39'sb111111110000000000000000000010000000000;
		7898: Delta = 39'sb000000001111111111111111111110000000000;
		3891: Delta = 39'sb111111101111111111111111111110000000000;
		5031: Delta = 39'sb000000100000000000000000000010000000000;
		10854: Delta = 39'sb111111100000000000000000000010000000000;
		2983: Delta = 39'sb000000011111111111111111111110000000000;
		8806: Delta = 39'sb111111011111111111111111111110000000000;
		9038: Delta = 39'sb000001000000000000000000000010000000000;
		6847: Delta = 39'sb111111000000000000000000000010000000000;
		6990: Delta = 39'sb000000111111111111111111111110000000000;
		4799: Delta = 39'sb111110111111111111111111111110000000000;
		3215: Delta = 39'sb000010000000000000000000000010000000000;
		12670: Delta = 39'sb111110000000000000000000000010000000000;
		1167: Delta = 39'sb000001111111111111111111111110000000000;
		10622: Delta = 39'sb111101111111111111111111111110000000000;
		5406: Delta = 39'sb000100000000000000000000000010000000000;
		10479: Delta = 39'sb111100000000000000000000000010000000000;
		3358: Delta = 39'sb000011111111111111111111111110000000000;
		8431: Delta = 39'sb111011111111111111111111111110000000000;
		9788: Delta = 39'sb001000000000000000000000000010000000000;
		6097: Delta = 39'sb111000000000000000000000000010000000000;
		7740: Delta = 39'sb000111111111111111111111111110000000000;
		4049: Delta = 39'sb110111111111111111111111111110000000000;
		4715: Delta = 39'sb010000000000000000000000000010000000000;
		11170: Delta = 39'sb110000000000000000000000000010000000000;
		2667: Delta = 39'sb001111111111111111111111111110000000000;
		9122: Delta = 39'sb101111111111111111111111111110000000000;
		6144: Delta = 39'sb000000000000000000000000001100000000000;
		7693: Delta = 39'sb111111111111111111111111110100000000000;
		10240: Delta = 39'sb000000000000000000000000010100000000000;
		3597: Delta = 39'sb111111111111111111111111101100000000000;
		4595: Delta = 39'sb000000000000000000000000100100000000000;
		13338: Delta = 39'sb111111111111111111111111100100000000000;
		499: Delta = 39'sb000000000000000000000000011100000000000;
		9242: Delta = 39'sb111111111111111111111111011100000000000;
		7142: Delta = 39'sb000000000000000000000001000100000000000;
		10791: Delta = 39'sb111111111111111111111111000100000000000;
		3046: Delta = 39'sb000000000000000000000000111100000000000;
		6695: Delta = 39'sb111111111111111111111110111100000000000;
		12236: Delta = 39'sb000000000000000000000010000100000000000;
		5697: Delta = 39'sb111111111111111111111110000100000000000;
		8140: Delta = 39'sb000000000000000000000001111100000000000;
		1601: Delta = 39'sb111111111111111111111101111100000000000;
		8587: Delta = 39'sb000000000000000000000100000100000000000;
		9346: Delta = 39'sb111111111111111111111100000100000000000;
		4491: Delta = 39'sb000000000000000000000011111100000000000;
		5250: Delta = 39'sb111111111111111111111011111100000000000;
		1289: Delta = 39'sb000000000000000000001000000100000000000;
		2807: Delta = 39'sb111111111111111111111000000100000000000;
		11030: Delta = 39'sb000000000000000000000111111100000000000;
		12548: Delta = 39'sb111111111111111111110111111100000000000;
		530: Delta = 39'sb000000000000000000010000000100000000000;
		3566: Delta = 39'sb111111111111111111110000000100000000000;
		10271: Delta = 39'sb000000000000000000001111111100000000000;
		13307: Delta = 39'sb111111111111111111101111111100000000000;
		12849: Delta = 39'sb000000000000000000100000000100000000000;
		5084: Delta = 39'sb111111111111111111100000000100000000000;
		8753: Delta = 39'sb000000000000000000011111111100000000000;
		988: Delta = 39'sb111111111111111111011111111100000000000;
		9813: Delta = 39'sb000000000000000001000000000100000000000;
		8120: Delta = 39'sb111111111111111111000000000100000000000;
		5717: Delta = 39'sb000000000000000000111111111100000000000;
		4024: Delta = 39'sb111111111111111110111111111100000000000;
		3741: Delta = 39'sb000000000000000010000000000100000000000;
		355: Delta = 39'sb111111111111111110000000000100000000000;
		13482: Delta = 39'sb000000000000000001111111111100000000000;
		10096: Delta = 39'sb111111111111111101111111111100000000000;
		5434: Delta = 39'sb000000000000000100000000000100000000000;
		12499: Delta = 39'sb111111111111111100000000000100000000000;
		1338: Delta = 39'sb000000000000000011111111111100000000000;
		8403: Delta = 39'sb111111111111111011111111111100000000000;
		8820: Delta = 39'sb000000000000001000000000000100000000000;
		9113: Delta = 39'sb111111111111111000000000000100000000000;
		4724: Delta = 39'sb000000000000000111111111111100000000000;
		5017: Delta = 39'sb111111111111110111111111111100000000000;
		1755: Delta = 39'sb000000000000010000000000000100000000000;
		2341: Delta = 39'sb111111111111110000000000000100000000000;
		11496: Delta = 39'sb000000000000001111111111111100000000000;
		12082: Delta = 39'sb111111111111101111111111111100000000000;
		1462: Delta = 39'sb000000000000100000000000000100000000000;
		2634: Delta = 39'sb111111111111100000000000000100000000000;
		11203: Delta = 39'sb000000000000011111111111111100000000000;
		12375: Delta = 39'sb111111111111011111111111111100000000000;
		876: Delta = 39'sb000000000001000000000000000100000000000;
		3220: Delta = 39'sb111111111111000000000000000100000000000;
		10617: Delta = 39'sb000000000000111111111111111100000000000;
		12961: Delta = 39'sb111111111110111111111111111100000000000;
		13541: Delta = 39'sb000000000010000000000000000100000000000;
		4392: Delta = 39'sb111111111110000000000000000100000000000;
		9445: Delta = 39'sb000000000001111111111111111100000000000;
		296: Delta = 39'sb111111111101111111111111111100000000000;
		11197: Delta = 39'sb000000000100000000000000000100000000000;
		6736: Delta = 39'sb111111111100000000000000000100000000000;
		7101: Delta = 39'sb000000000011111111111111111100000000000;
		2640: Delta = 39'sb111111111011111111111111111100000000000;
		6509: Delta = 39'sb000000001000000000000000000100000000000;
		11424: Delta = 39'sb111111111000000000000000000100000000000;
		2413: Delta = 39'sb000000000111111111111111111100000000000;
		7328: Delta = 39'sb111111110111111111111111111100000000000;
		10970: Delta = 39'sb000000010000000000000000000100000000000;
		6963: Delta = 39'sb111111110000000000000000000100000000000;
		6874: Delta = 39'sb000000001111111111111111111100000000000;
		2867: Delta = 39'sb111111101111111111111111111100000000000;
		6055: Delta = 39'sb000000100000000000000000000100000000000;
		11878: Delta = 39'sb111111100000000000000000000100000000000;
		1959: Delta = 39'sb000000011111111111111111111100000000000;
		7782: Delta = 39'sb111111011111111111111111111100000000000;
		10062: Delta = 39'sb000001000000000000000000000100000000000;
		7871: Delta = 39'sb111111000000000000000000000100000000000;
		5966: Delta = 39'sb000000111111111111111111111100000000000;
		3775: Delta = 39'sb111110111111111111111111111100000000000;
		4239: Delta = 39'sb000010000000000000000000000100000000000;
		13694: Delta = 39'sb111110000000000000000000000100000000000;
		143: Delta = 39'sb000001111111111111111111111100000000000;
		9598: Delta = 39'sb111101111111111111111111111100000000000;
		6430: Delta = 39'sb000100000000000000000000000100000000000;
		11503: Delta = 39'sb111100000000000000000000000100000000000;
		2334: Delta = 39'sb000011111111111111111111111100000000000;
		7407: Delta = 39'sb111011111111111111111111111100000000000;
		10812: Delta = 39'sb001000000000000000000000000100000000000;
		7121: Delta = 39'sb111000000000000000000000000100000000000;
		6716: Delta = 39'sb000111111111111111111111111100000000000;
		3025: Delta = 39'sb110111111111111111111111111100000000000;
		5739: Delta = 39'sb010000000000000000000000000100000000000;
		12194: Delta = 39'sb110000000000000000000000000100000000000;
		1643: Delta = 39'sb001111111111111111111111111100000000000;
		8098: Delta = 39'sb101111111111111111111111111100000000000;
		12288: Delta = 39'sb000000000000000000000000011000000000000;
		1549: Delta = 39'sb111111111111111111111111101000000000000;
		6643: Delta = 39'sb000000000000000000000000101000000000000;
		7194: Delta = 39'sb111111111111111111111111011000000000000;
		9190: Delta = 39'sb000000000000000000000001001000000000000;
		12839: Delta = 39'sb111111111111111111111111001000000000000;
		998: Delta = 39'sb000000000000000000000000111000000000000;
		4647: Delta = 39'sb111111111111111111111110111000000000000;
		447: Delta = 39'sb000000000000000000000010001000000000000;
		7745: Delta = 39'sb111111111111111111111110001000000000000;
		6092: Delta = 39'sb000000000000000000000001111000000000000;
		13390: Delta = 39'sb111111111111111111111101111000000000000;
		10635: Delta = 39'sb000000000000000000000100001000000000000;
		11394: Delta = 39'sb111111111111111111111100001000000000000;
		2443: Delta = 39'sb000000000000000000000011111000000000000;
		3202: Delta = 39'sb111111111111111111111011111000000000000;
		3337: Delta = 39'sb000000000000000000001000001000000000000;
		4855: Delta = 39'sb111111111111111111111000001000000000000;
		8982: Delta = 39'sb000000000000000000000111111000000000000;
		10500: Delta = 39'sb111111111111111111110111111000000000000;
		2578: Delta = 39'sb000000000000000000010000001000000000000;
		5614: Delta = 39'sb111111111111111111110000001000000000000;
		8223: Delta = 39'sb000000000000000000001111111000000000000;
		11259: Delta = 39'sb111111111111111111101111111000000000000;
		1060: Delta = 39'sb000000000000000000100000001000000000000;
		7132: Delta = 39'sb111111111111111111100000001000000000000;
		6705: Delta = 39'sb000000000000000000011111111000000000000;
		12777: Delta = 39'sb111111111111111111011111111000000000000;
		11861: Delta = 39'sb000000000000000001000000001000000000000;
		10168: Delta = 39'sb111111111111111111000000001000000000000;
		3669: Delta = 39'sb000000000000000000111111111000000000000;
		1976: Delta = 39'sb111111111111111110111111111000000000000;
		5789: Delta = 39'sb000000000000000010000000001000000000000;
		2403: Delta = 39'sb111111111111111110000000001000000000000;
		11434: Delta = 39'sb000000000000000001111111111000000000000;
		8048: Delta = 39'sb111111111111111101111111111000000000000;
		7482: Delta = 39'sb000000000000000100000000001000000000000;
		710: Delta = 39'sb111111111111111100000000001000000000000;
		13127: Delta = 39'sb000000000000000011111111111000000000000;
		6355: Delta = 39'sb111111111111111011111111111000000000000;
		10868: Delta = 39'sb000000000000001000000000001000000000000;
		11161: Delta = 39'sb111111111111111000000000001000000000000;
		2676: Delta = 39'sb000000000000000111111111111000000000000;
		2969: Delta = 39'sb111111111111110111111111111000000000000;
		3803: Delta = 39'sb000000000000010000000000001000000000000;
		4389: Delta = 39'sb111111111111110000000000001000000000000;
		9448: Delta = 39'sb000000000000001111111111111000000000000;
		10034: Delta = 39'sb111111111111101111111111111000000000000;
		3510: Delta = 39'sb000000000000100000000000001000000000000;
		4682: Delta = 39'sb111111111111100000000000001000000000000;
		9155: Delta = 39'sb000000000000011111111111111000000000000;
		10327: Delta = 39'sb111111111111011111111111111000000000000;
		2924: Delta = 39'sb000000000001000000000000001000000000000;
		5268: Delta = 39'sb111111111111000000000000001000000000000;
		8569: Delta = 39'sb000000000000111111111111111000000000000;
		10913: Delta = 39'sb111111111110111111111111111000000000000;
		1752: Delta = 39'sb000000000010000000000000001000000000000;
		6440: Delta = 39'sb111111111110000000000000001000000000000;
		7397: Delta = 39'sb000000000001111111111111111000000000000;
		12085: Delta = 39'sb111111111101111111111111111000000000000;
		13245: Delta = 39'sb000000000100000000000000001000000000000;
		8784: Delta = 39'sb111111111100000000000000001000000000000;
		5053: Delta = 39'sb000000000011111111111111111000000000000;
		592: Delta = 39'sb111111111011111111111111111000000000000;
		8557: Delta = 39'sb000000001000000000000000001000000000000;
		13472: Delta = 39'sb111111111000000000000000001000000000000;
		365: Delta = 39'sb000000000111111111111111111000000000000;
		5280: Delta = 39'sb111111110111111111111111111000000000000;
		13018: Delta = 39'sb000000010000000000000000001000000000000;
		9011: Delta = 39'sb111111110000000000000000001000000000000;
		4826: Delta = 39'sb000000001111111111111111111000000000000;
		819: Delta = 39'sb111111101111111111111111111000000000000;
		8103: Delta = 39'sb000000100000000000000000001000000000000;
		89: Delta = 39'sb111111100000000000000000001000000000000;
		13748: Delta = 39'sb000000011111111111111111111000000000000;
		5734: Delta = 39'sb111111011111111111111111111000000000000;
		12110: Delta = 39'sb000001000000000000000000001000000000000;
		9919: Delta = 39'sb111111000000000000000000001000000000000;
		3918: Delta = 39'sb000000111111111111111111111000000000000;
		1727: Delta = 39'sb111110111111111111111111111000000000000;
		6287: Delta = 39'sb000010000000000000000000001000000000000;
		1905: Delta = 39'sb111110000000000000000000001000000000000;
		11932: Delta = 39'sb000001111111111111111111111000000000000;
		7550: Delta = 39'sb111101111111111111111111111000000000000;
		8478: Delta = 39'sb000100000000000000000000001000000000000;
		13551: Delta = 39'sb111100000000000000000000001000000000000;
		286: Delta = 39'sb000011111111111111111111111000000000000;
		5359: Delta = 39'sb111011111111111111111111111000000000000;
		12860: Delta = 39'sb001000000000000000000000001000000000000;
		9169: Delta = 39'sb111000000000000000000000001000000000000;
		4668: Delta = 39'sb000111111111111111111111111000000000000;
		977: Delta = 39'sb110111111111111111111111111000000000000;
		7787: Delta = 39'sb010000000000000000000000001000000000000;
		405: Delta = 39'sb110000000000000000000000001000000000000;
		13432: Delta = 39'sb001111111111111111111111111000000000000;
		6050: Delta = 39'sb101111111111111111111111111000000000000;
		10739: Delta = 39'sb000000000000000000000000110000000000000;
		3098: Delta = 39'sb111111111111111111111111010000000000000;
		13286: Delta = 39'sb000000000000000000000001010000000000000;
		551: Delta = 39'sb111111111111111111111110110000000000000;
		4543: Delta = 39'sb000000000000000000000010010000000000000;
		11841: Delta = 39'sb111111111111111111111110010000000000000;
		1996: Delta = 39'sb000000000000000000000001110000000000000;
		9294: Delta = 39'sb111111111111111111111101110000000000000;
		894: Delta = 39'sb000000000000000000000100010000000000000;
		1653: Delta = 39'sb111111111111111111111100010000000000000;
		12184: Delta = 39'sb000000000000000000000011110000000000000;
		12943: Delta = 39'sb111111111111111111111011110000000000000;
		7433: Delta = 39'sb000000000000000000001000010000000000000;
		8951: Delta = 39'sb111111111111111111111000010000000000000;
		4886: Delta = 39'sb000000000000000000000111110000000000000;
		6404: Delta = 39'sb111111111111111111110111110000000000000;
		6674: Delta = 39'sb000000000000000000010000010000000000000;
		9710: Delta = 39'sb111111111111111111110000010000000000000;
		4127: Delta = 39'sb000000000000000000001111110000000000000;
		7163: Delta = 39'sb111111111111111111101111110000000000000;
		5156: Delta = 39'sb000000000000000000100000010000000000000;
		11228: Delta = 39'sb111111111111111111100000010000000000000;
		2609: Delta = 39'sb000000000000000000011111110000000000000;
		8681: Delta = 39'sb111111111111111111011111110000000000000;
		2120: Delta = 39'sb000000000000000001000000010000000000000;
		427: Delta = 39'sb111111111111111111000000010000000000000;
		13410: Delta = 39'sb000000000000000000111111110000000000000;
		11717: Delta = 39'sb111111111111111110111111110000000000000;
		9885: Delta = 39'sb000000000000000010000000010000000000000;
		6499: Delta = 39'sb111111111111111110000000010000000000000;
		7338: Delta = 39'sb000000000000000001111111110000000000000;
		3952: Delta = 39'sb111111111111111101111111110000000000000;
		11578: Delta = 39'sb000000000000000100000000010000000000000;
		4806: Delta = 39'sb111111111111111100000000010000000000000;
		9031: Delta = 39'sb000000000000000011111111110000000000000;
		2259: Delta = 39'sb111111111111111011111111110000000000000;
		1127: Delta = 39'sb000000000000001000000000010000000000000;
		1420: Delta = 39'sb111111111111111000000000010000000000000;
		12417: Delta = 39'sb000000000000000111111111110000000000000;
		12710: Delta = 39'sb111111111111110111111111110000000000000;
		7899: Delta = 39'sb000000000000010000000000010000000000000;
		8485: Delta = 39'sb111111111111110000000000010000000000000;
		5352: Delta = 39'sb000000000000001111111111110000000000000;
		5938: Delta = 39'sb111111111111101111111111110000000000000;
		7606: Delta = 39'sb000000000000100000000000010000000000000;
		8778: Delta = 39'sb111111111111100000000000010000000000000;
		5059: Delta = 39'sb000000000000011111111111110000000000000;
		6231: Delta = 39'sb111111111111011111111111110000000000000;
		7020: Delta = 39'sb000000000001000000000000010000000000000;
		9364: Delta = 39'sb111111111111000000000000010000000000000;
		4473: Delta = 39'sb000000000000111111111111110000000000000;
		6817: Delta = 39'sb111111111110111111111111110000000000000;
		5848: Delta = 39'sb000000000010000000000000010000000000000;
		10536: Delta = 39'sb111111111110000000000000010000000000000;
		3301: Delta = 39'sb000000000001111111111111110000000000000;
		7989: Delta = 39'sb111111111101111111111111110000000000000;
		3504: Delta = 39'sb000000000100000000000000010000000000000;
		12880: Delta = 39'sb111111111100000000000000010000000000000;
		957: Delta = 39'sb000000000011111111111111110000000000000;
		10333: Delta = 39'sb111111111011111111111111110000000000000;
		12653: Delta = 39'sb000000001000000000000000010000000000000;
		3731: Delta = 39'sb111111111000000000000000010000000000000;
		10106: Delta = 39'sb000000000111111111111111110000000000000;
		1184: Delta = 39'sb111111110111111111111111110000000000000;
		3277: Delta = 39'sb000000010000000000000000010000000000000;
		13107: Delta = 39'sb111111110000000000000000010000000000000;
		730: Delta = 39'sb000000001111111111111111110000000000000;
		10560: Delta = 39'sb111111101111111111111111110000000000000;
		12199: Delta = 39'sb000000100000000000000000010000000000000;
		4185: Delta = 39'sb111111100000000000000000010000000000000;
		9652: Delta = 39'sb000000011111111111111111110000000000000;
		1638: Delta = 39'sb111111011111111111111111110000000000000;
		2369: Delta = 39'sb000001000000000000000000010000000000000;
		178: Delta = 39'sb111111000000000000000000010000000000000;
		13659: Delta = 39'sb000000111111111111111111110000000000000;
		11468: Delta = 39'sb111110111111111111111111110000000000000;
		10383: Delta = 39'sb000010000000000000000000010000000000000;
		6001: Delta = 39'sb111110000000000000000000010000000000000;
		7836: Delta = 39'sb000001111111111111111111110000000000000;
		3454: Delta = 39'sb111101111111111111111111110000000000000;
		12574: Delta = 39'sb000100000000000000000000010000000000000;
		3810: Delta = 39'sb111100000000000000000000010000000000000;
		10027: Delta = 39'sb000011111111111111111111110000000000000;
		1263: Delta = 39'sb111011111111111111111111110000000000000;
		3119: Delta = 39'sb001000000000000000000000010000000000000;
		13265: Delta = 39'sb111000000000000000000000010000000000000;
		572: Delta = 39'sb000111111111111111111111110000000000000;
		10718: Delta = 39'sb110111111111111111111111110000000000000;
		11883: Delta = 39'sb010000000000000000000000010000000000000;
		4501: Delta = 39'sb110000000000000000000000010000000000000;
		9336: Delta = 39'sb001111111111111111111111110000000000000;
		1954: Delta = 39'sb101111111111111111111111110000000000000;
		7641: Delta = 39'sb000000000000000000000001100000000000000;
		6196: Delta = 39'sb111111111111111111111110100000000000000;
		12735: Delta = 39'sb000000000000000000000010100000000000000;
		1102: Delta = 39'sb111111111111111111111101100000000000000;
		9086: Delta = 39'sb000000000000000000000100100000000000000;
		9845: Delta = 39'sb111111111111111111111100100000000000000;
		3992: Delta = 39'sb000000000000000000000011100000000000000;
		4751: Delta = 39'sb111111111111111111111011100000000000000;
		1788: Delta = 39'sb000000000000000000001000100000000000000;
		3306: Delta = 39'sb111111111111111111111000100000000000000;
		10531: Delta = 39'sb000000000000000000000111100000000000000;
		12049: Delta = 39'sb111111111111111111110111100000000000000;
		1029: Delta = 39'sb000000000000000000010000100000000000000;
		4065: Delta = 39'sb111111111111111111110000100000000000000;
		9772: Delta = 39'sb000000000000000000001111100000000000000;
		12808: Delta = 39'sb111111111111111111101111100000000000000;
		13348: Delta = 39'sb000000000000000000100000100000000000000;
		5583: Delta = 39'sb111111111111111111100000100000000000000;
		8254: Delta = 39'sb000000000000000000011111100000000000000;
		489: Delta = 39'sb111111111111111111011111100000000000000;
		10312: Delta = 39'sb000000000000000001000000100000000000000;
		8619: Delta = 39'sb111111111111111111000000100000000000000;
		5218: Delta = 39'sb000000000000000000111111100000000000000;
		3525: Delta = 39'sb111111111111111110111111100000000000000;
		4240: Delta = 39'sb000000000000000010000000100000000000000;
		854: Delta = 39'sb111111111111111110000000100000000000000;
		12983: Delta = 39'sb000000000000000001111111100000000000000;
		9597: Delta = 39'sb111111111111111101111111100000000000000;
		5933: Delta = 39'sb000000000000000100000000100000000000000;
		12998: Delta = 39'sb111111111111111100000000100000000000000;
		839: Delta = 39'sb000000000000000011111111100000000000000;
		7904: Delta = 39'sb111111111111111011111111100000000000000;
		9319: Delta = 39'sb000000000000001000000000100000000000000;
		9612: Delta = 39'sb111111111111111000000000100000000000000;
		4225: Delta = 39'sb000000000000000111111111100000000000000;
		4518: Delta = 39'sb111111111111110111111111100000000000000;
		2254: Delta = 39'sb000000000000010000000000100000000000000;
		2840: Delta = 39'sb111111111111110000000000100000000000000;
		10997: Delta = 39'sb000000000000001111111111100000000000000;
		11583: Delta = 39'sb111111111111101111111111100000000000000;
		1961: Delta = 39'sb000000000000100000000000100000000000000;
		3133: Delta = 39'sb111111111111100000000000100000000000000;
		10704: Delta = 39'sb000000000000011111111111100000000000000;
		11876: Delta = 39'sb111111111111011111111111100000000000000;
		1375: Delta = 39'sb000000000001000000000000100000000000000;
		3719: Delta = 39'sb111111111111000000000000100000000000000;
		10118: Delta = 39'sb000000000000111111111111100000000000000;
		12462: Delta = 39'sb111111111110111111111111100000000000000;
		203: Delta = 39'sb000000000010000000000000100000000000000;
		4891: Delta = 39'sb111111111110000000000000100000000000000;
		8946: Delta = 39'sb000000000001111111111111100000000000000;
		13634: Delta = 39'sb111111111101111111111111100000000000000;
		11696: Delta = 39'sb000000000100000000000000100000000000000;
		7235: Delta = 39'sb111111111100000000000000100000000000000;
		6602: Delta = 39'sb000000000011111111111111100000000000000;
		2141: Delta = 39'sb111111111011111111111111100000000000000;
		7008: Delta = 39'sb000000001000000000000000100000000000000;
		11923: Delta = 39'sb111111111000000000000000100000000000000;
		1914: Delta = 39'sb000000000111111111111111100000000000000;
		6829: Delta = 39'sb111111110111111111111111100000000000000;
		11469: Delta = 39'sb000000010000000000000000100000000000000;
		7462: Delta = 39'sb111111110000000000000000100000000000000;
		6375: Delta = 39'sb000000001111111111111111100000000000000;
		2368: Delta = 39'sb111111101111111111111111100000000000000;
		6554: Delta = 39'sb000000100000000000000000100000000000000;
		12377: Delta = 39'sb111111100000000000000000100000000000000;
		1460: Delta = 39'sb000000011111111111111111100000000000000;
		7283: Delta = 39'sb111111011111111111111111100000000000000;
		10561: Delta = 39'sb000001000000000000000000100000000000000;
		8370: Delta = 39'sb111111000000000000000000100000000000000;
		5467: Delta = 39'sb000000111111111111111111100000000000000;
		3276: Delta = 39'sb111110111111111111111111100000000000000;
		4738: Delta = 39'sb000010000000000000000000100000000000000;
		356: Delta = 39'sb111110000000000000000000100000000000000;
		13481: Delta = 39'sb000001111111111111111111100000000000000;
		9099: Delta = 39'sb111101111111111111111111100000000000000;
		6929: Delta = 39'sb000100000000000000000000100000000000000;
		12002: Delta = 39'sb111100000000000000000000100000000000000;
		1835: Delta = 39'sb000011111111111111111111100000000000000;
		6908: Delta = 39'sb111011111111111111111111100000000000000;
		11311: Delta = 39'sb001000000000000000000000100000000000000;
		7620: Delta = 39'sb111000000000000000000000100000000000000;
		6217: Delta = 39'sb000111111111111111111111100000000000000;
		2526: Delta = 39'sb110111111111111111111111100000000000000;
		6238: Delta = 39'sb010000000000000000000000100000000000000;
		12693: Delta = 39'sb110000000000000000000000100000000000000;
		1144: Delta = 39'sb001111111111111111111111100000000000000;
		7599: Delta = 39'sb101111111111111111111111100000000000000;
		1445: Delta = 39'sb000000000000000000000011000000000000000;
		12392: Delta = 39'sb111111111111111111111101000000000000000;
		11633: Delta = 39'sb000000000000000000000101000000000000000;
		2204: Delta = 39'sb111111111111111111111011000000000000000;
		4335: Delta = 39'sb000000000000000000001001000000000000000;
		5853: Delta = 39'sb111111111111111111111001000000000000000;
		7984: Delta = 39'sb000000000000000000000111000000000000000;
		9502: Delta = 39'sb111111111111111111110111000000000000000;
		3576: Delta = 39'sb000000000000000000010001000000000000000;
		6612: Delta = 39'sb111111111111111111110001000000000000000;
		7225: Delta = 39'sb000000000000000000001111000000000000000;
		10261: Delta = 39'sb111111111111111111101111000000000000000;
		2058: Delta = 39'sb000000000000000000100001000000000000000;
		8130: Delta = 39'sb111111111111111111100001000000000000000;
		5707: Delta = 39'sb000000000000000000011111000000000000000;
		11779: Delta = 39'sb111111111111111111011111000000000000000;
		12859: Delta = 39'sb000000000000000001000001000000000000000;
		11166: Delta = 39'sb111111111111111111000001000000000000000;
		2671: Delta = 39'sb000000000000000000111111000000000000000;
		978: Delta = 39'sb111111111111111110111111000000000000000;
		6787: Delta = 39'sb000000000000000010000001000000000000000;
		3401: Delta = 39'sb111111111111111110000001000000000000000;
		10436: Delta = 39'sb000000000000000001111111000000000000000;
		7050: Delta = 39'sb111111111111111101111111000000000000000;
		8480: Delta = 39'sb000000000000000100000001000000000000000;
		1708: Delta = 39'sb111111111111111100000001000000000000000;
		12129: Delta = 39'sb000000000000000011111111000000000000000;
		5357: Delta = 39'sb111111111111111011111111000000000000000;
		11866: Delta = 39'sb000000000000001000000001000000000000000;
		12159: Delta = 39'sb111111111111111000000001000000000000000;
		1678: Delta = 39'sb000000000000000111111111000000000000000;
		1971: Delta = 39'sb111111111111110111111111000000000000000;
		4801: Delta = 39'sb000000000000010000000001000000000000000;
		5387: Delta = 39'sb111111111111110000000001000000000000000;
		8450: Delta = 39'sb000000000000001111111111000000000000000;
		9036: Delta = 39'sb111111111111101111111111000000000000000;
		4508: Delta = 39'sb000000000000100000000001000000000000000;
		5680: Delta = 39'sb111111111111100000000001000000000000000;
		8157: Delta = 39'sb000000000000011111111111000000000000000;
		9329: Delta = 39'sb111111111111011111111111000000000000000;
		3922: Delta = 39'sb000000000001000000000001000000000000000;
		6266: Delta = 39'sb111111111111000000000001000000000000000;
		7571: Delta = 39'sb000000000000111111111111000000000000000;
		9915: Delta = 39'sb111111111110111111111111000000000000000;
		2750: Delta = 39'sb000000000010000000000001000000000000000;
		7438: Delta = 39'sb111111111110000000000001000000000000000;
		6399: Delta = 39'sb000000000001111111111111000000000000000;
		11087: Delta = 39'sb111111111101111111111111000000000000000;
		406: Delta = 39'sb000000000100000000000001000000000000000;
		9782: Delta = 39'sb111111111100000000000001000000000000000;
		4055: Delta = 39'sb000000000011111111111111000000000000000;
		13431: Delta = 39'sb111111111011111111111111000000000000000;
		9555: Delta = 39'sb000000001000000000000001000000000000000;
		633: Delta = 39'sb111111111000000000000001000000000000000;
		13204: Delta = 39'sb000000000111111111111111000000000000000;
		4282: Delta = 39'sb111111110111111111111111000000000000000;
		179: Delta = 39'sb000000010000000000000001000000000000000;
		10009: Delta = 39'sb111111110000000000000001000000000000000;
		3828: Delta = 39'sb000000001111111111111111000000000000000;
		13658: Delta = 39'sb111111101111111111111111000000000000000;
		9101: Delta = 39'sb000000100000000000000001000000000000000;
		1087: Delta = 39'sb111111100000000000000001000000000000000;
		12750: Delta = 39'sb000000011111111111111111000000000000000;
		4736: Delta = 39'sb111111011111111111111111000000000000000;
		13108: Delta = 39'sb000001000000000000000001000000000000000;
		10917: Delta = 39'sb111111000000000000000001000000000000000;
		2920: Delta = 39'sb000000111111111111111111000000000000000;
		729: Delta = 39'sb111110111111111111111111000000000000000;
		7285: Delta = 39'sb000010000000000000000001000000000000000;
		2903: Delta = 39'sb111110000000000000000001000000000000000;
		10934: Delta = 39'sb000001111111111111111111000000000000000;
		6552: Delta = 39'sb111101111111111111111111000000000000000;
		9476: Delta = 39'sb000100000000000000000001000000000000000;
		712: Delta = 39'sb111100000000000000000001000000000000000;
		13125: Delta = 39'sb000011111111111111111111000000000000000;
		4361: Delta = 39'sb111011111111111111111111000000000000000;
		21: Delta = 39'sb001000000000000000000001000000000000000;
		10167: Delta = 39'sb111000000000000000000001000000000000000;
		3670: Delta = 39'sb000111111111111111111111000000000000000;
		13816: Delta = 39'sb110111111111111111111111000000000000000;
		8785: Delta = 39'sb010000000000000000000001000000000000000;
		1403: Delta = 39'sb110000000000000000000001000000000000000;
		12434: Delta = 39'sb001111111111111111111111000000000000000;
		5052: Delta = 39'sb101111111111111111111111000000000000000;
		2890: Delta = 39'sb000000000000000000000110000000000000000;
		10947: Delta = 39'sb111111111111111111111010000000000000000;
		9429: Delta = 39'sb000000000000000000001010000000000000000;
		4408: Delta = 39'sb111111111111111111110110000000000000000;
		8670: Delta = 39'sb000000000000000000010010000000000000000;
		11706: Delta = 39'sb111111111111111111110010000000000000000;
		2131: Delta = 39'sb000000000000000000001110000000000000000;
		5167: Delta = 39'sb111111111111111111101110000000000000000;
		7152: Delta = 39'sb000000000000000000100010000000000000000;
		13224: Delta = 39'sb111111111111111111100010000000000000000;
		613: Delta = 39'sb000000000000000000011110000000000000000;
		6685: Delta = 39'sb111111111111111111011110000000000000000;
		4116: Delta = 39'sb000000000000000001000010000000000000000;
		2423: Delta = 39'sb111111111111111111000010000000000000000;
		11414: Delta = 39'sb000000000000000000111110000000000000000;
		9721: Delta = 39'sb111111111111111110111110000000000000000;
		11881: Delta = 39'sb000000000000000010000010000000000000000;
		8495: Delta = 39'sb111111111111111110000010000000000000000;
		5342: Delta = 39'sb000000000000000001111110000000000000000;
		1956: Delta = 39'sb111111111111111101111110000000000000000;
		13574: Delta = 39'sb000000000000000100000010000000000000000;
		6802: Delta = 39'sb111111111111111100000010000000000000000;
		7035: Delta = 39'sb000000000000000011111110000000000000000;
		263: Delta = 39'sb111111111111111011111110000000000000000;
		3123: Delta = 39'sb000000000000001000000010000000000000000;
		3416: Delta = 39'sb111111111111111000000010000000000000000;
		10421: Delta = 39'sb000000000000000111111110000000000000000;
		10714: Delta = 39'sb111111111111110111111110000000000000000;
		9895: Delta = 39'sb000000000000010000000010000000000000000;
		10481: Delta = 39'sb111111111111110000000010000000000000000;
		3356: Delta = 39'sb000000000000001111111110000000000000000;
		3942: Delta = 39'sb111111111111101111111110000000000000000;
		9602: Delta = 39'sb000000000000100000000010000000000000000;
		10774: Delta = 39'sb111111111111100000000010000000000000000;
		3063: Delta = 39'sb000000000000011111111110000000000000000;
		4235: Delta = 39'sb111111111111011111111110000000000000000;
		9016: Delta = 39'sb000000000001000000000010000000000000000;
		11360: Delta = 39'sb111111111111000000000010000000000000000;
		2477: Delta = 39'sb000000000000111111111110000000000000000;
		4821: Delta = 39'sb111111111110111111111110000000000000000;
		7844: Delta = 39'sb000000000010000000000010000000000000000;
		12532: Delta = 39'sb111111111110000000000010000000000000000;
		1305: Delta = 39'sb000000000001111111111110000000000000000;
		5993: Delta = 39'sb111111111101111111111110000000000000000;
		5500: Delta = 39'sb000000000100000000000010000000000000000;
		1039: Delta = 39'sb111111111100000000000010000000000000000;
		12798: Delta = 39'sb000000000011111111111110000000000000000;
		8337: Delta = 39'sb111111111011111111111110000000000000000;
		812: Delta = 39'sb000000001000000000000010000000000000000;
		5727: Delta = 39'sb111111111000000000000010000000000000000;
		8110: Delta = 39'sb000000000111111111111110000000000000000;
		13025: Delta = 39'sb111111110111111111111110000000000000000;
		5273: Delta = 39'sb000000010000000000000010000000000000000;
		1266: Delta = 39'sb111111110000000000000010000000000000000;
		12571: Delta = 39'sb000000001111111111111110000000000000000;
		8564: Delta = 39'sb111111101111111111111110000000000000000;
		358: Delta = 39'sb000000100000000000000010000000000000000;
		6181: Delta = 39'sb111111100000000000000010000000000000000;
		7656: Delta = 39'sb000000011111111111111110000000000000000;
		13479: Delta = 39'sb111111011111111111111110000000000000000;
		4365: Delta = 39'sb000001000000000000000010000000000000000;
		2174: Delta = 39'sb111111000000000000000010000000000000000;
		11663: Delta = 39'sb000000111111111111111110000000000000000;
		9472: Delta = 39'sb111110111111111111111110000000000000000;
		12379: Delta = 39'sb000010000000000000000010000000000000000;
		7997: Delta = 39'sb111110000000000000000010000000000000000;
		5840: Delta = 39'sb000001111111111111111110000000000000000;
		1458: Delta = 39'sb111101111111111111111110000000000000000;
		733: Delta = 39'sb000100000000000000000010000000000000000;
		5806: Delta = 39'sb111100000000000000000010000000000000000;
		8031: Delta = 39'sb000011111111111111111110000000000000000;
		13104: Delta = 39'sb111011111111111111111110000000000000000;
		5115: Delta = 39'sb001000000000000000000010000000000000000;
		1424: Delta = 39'sb111000000000000000000010000000000000000;
		12413: Delta = 39'sb000111111111111111111110000000000000000;
		8722: Delta = 39'sb110111111111111111111110000000000000000;
		42: Delta = 39'sb010000000000000000000010000000000000000;
		6497: Delta = 39'sb110000000000000000000010000000000000000;
		7340: Delta = 39'sb001111111111111111111110000000000000000;
		13795: Delta = 39'sb101111111111111111111110000000000000000;
		5780: Delta = 39'sb000000000000000000001100000000000000000;
		8057: Delta = 39'sb111111111111111111110100000000000000000;
		5021: Delta = 39'sb000000000000000000010100000000000000000;
		8816: Delta = 39'sb111111111111111111101100000000000000000;
		3503: Delta = 39'sb000000000000000000100100000000000000000;
		9575: Delta = 39'sb111111111111111111100100000000000000000;
		4262: Delta = 39'sb000000000000000000011100000000000000000;
		10334: Delta = 39'sb111111111111111111011100000000000000000;
		467: Delta = 39'sb000000000000000001000100000000000000000;
		12611: Delta = 39'sb111111111111111111000100000000000000000;
		1226: Delta = 39'sb000000000000000000111100000000000000000;
		13370: Delta = 39'sb111111111111111110111100000000000000000;
		8232: Delta = 39'sb000000000000000010000100000000000000000;
		4846: Delta = 39'sb111111111111111110000100000000000000000;
		8991: Delta = 39'sb000000000000000001111100000000000000000;
		5605: Delta = 39'sb111111111111111101111100000000000000000;
		9925: Delta = 39'sb000000000000000100000100000000000000000;
		3153: Delta = 39'sb111111111111111100000100000000000000000;
		10684: Delta = 39'sb000000000000000011111100000000000000000;
		3912: Delta = 39'sb111111111111111011111100000000000000000;
		13311: Delta = 39'sb000000000000001000000100000000000000000;
		13604: Delta = 39'sb111111111111111000000100000000000000000;
		233: Delta = 39'sb000000000000000111111100000000000000000;
		526: Delta = 39'sb111111111111110111111100000000000000000;
		6246: Delta = 39'sb000000000000010000000100000000000000000;
		6832: Delta = 39'sb111111111111110000000100000000000000000;
		7005: Delta = 39'sb000000000000001111111100000000000000000;
		7591: Delta = 39'sb111111111111101111111100000000000000000;
		5953: Delta = 39'sb000000000000100000000100000000000000000;
		7125: Delta = 39'sb111111111111100000000100000000000000000;
		6712: Delta = 39'sb000000000000011111111100000000000000000;
		7884: Delta = 39'sb111111111111011111111100000000000000000;
		5367: Delta = 39'sb000000000001000000000100000000000000000;
		7711: Delta = 39'sb111111111111000000000100000000000000000;
		6126: Delta = 39'sb000000000000111111111100000000000000000;
		8470: Delta = 39'sb111111111110111111111100000000000000000;
		4195: Delta = 39'sb000000000010000000000100000000000000000;
		8883: Delta = 39'sb111111111110000000000100000000000000000;
		4954: Delta = 39'sb000000000001111111111100000000000000000;
		9642: Delta = 39'sb111111111101111111111100000000000000000;
		1851: Delta = 39'sb000000000100000000000100000000000000000;
		11227: Delta = 39'sb111111111100000000000100000000000000000;
		2610: Delta = 39'sb000000000011111111111100000000000000000;
		11986: Delta = 39'sb111111111011111111111100000000000000000;
		11000: Delta = 39'sb000000001000000000000100000000000000000;
		2078: Delta = 39'sb111111111000000000000100000000000000000;
		11759: Delta = 39'sb000000000111111111111100000000000000000;
		2837: Delta = 39'sb111111110111111111111100000000000000000;
		1624: Delta = 39'sb000000010000000000000100000000000000000;
		11454: Delta = 39'sb111111110000000000000100000000000000000;
		2383: Delta = 39'sb000000001111111111111100000000000000000;
		12213: Delta = 39'sb111111101111111111111100000000000000000;
		10546: Delta = 39'sb000000100000000000000100000000000000000;
		2532: Delta = 39'sb111111100000000000000100000000000000000;
		11305: Delta = 39'sb000000011111111111111100000000000000000;
		3291: Delta = 39'sb111111011111111111111100000000000000000;
		716: Delta = 39'sb000001000000000000000100000000000000000;
		12362: Delta = 39'sb111111000000000000000100000000000000000;
		1475: Delta = 39'sb000000111111111111111100000000000000000;
		13121: Delta = 39'sb111110111111111111111100000000000000000;
		8730: Delta = 39'sb000010000000000000000100000000000000000;
		4348: Delta = 39'sb111110000000000000000100000000000000000;
		9489: Delta = 39'sb000001111111111111111100000000000000000;
		5107: Delta = 39'sb111101111111111111111100000000000000000;
		10921: Delta = 39'sb000100000000000000000100000000000000000;
		2157: Delta = 39'sb111100000000000000000100000000000000000;
		11680: Delta = 39'sb000011111111111111111100000000000000000;
		2916: Delta = 39'sb111011111111111111111100000000000000000;
		1466: Delta = 39'sb001000000000000000000100000000000000000;
		11612: Delta = 39'sb111000000000000000000100000000000000000;
		2225: Delta = 39'sb000111111111111111111100000000000000000;
		12371: Delta = 39'sb110111111111111111111100000000000000000;
		10230: Delta = 39'sb010000000000000000000100000000000000000;
		2848: Delta = 39'sb110000000000000000000100000000000000000;
		10989: Delta = 39'sb001111111111111111111100000000000000000;
		3607: Delta = 39'sb101111111111111111111100000000000000000;
		11560: Delta = 39'sb000000000000000000011000000000000000000;
		2277: Delta = 39'sb111111111111111111101000000000000000000;
		10042: Delta = 39'sb000000000000000000101000000000000000000;
		3795: Delta = 39'sb111111111111111111011000000000000000000;
		7006: Delta = 39'sb000000000000000001001000000000000000000;
		5313: Delta = 39'sb111111111111111111001000000000000000000;
		8524: Delta = 39'sb000000000000000000111000000000000000000;
		6831: Delta = 39'sb111111111111111110111000000000000000000;
		934: Delta = 39'sb000000000000000010001000000000000000000;
		11385: Delta = 39'sb111111111111111110001000000000000000000;
		2452: Delta = 39'sb000000000000000001111000000000000000000;
		12903: Delta = 39'sb111111111111111101111000000000000000000;
		2627: Delta = 39'sb000000000000000100001000000000000000000;
		9692: Delta = 39'sb111111111111111100001000000000000000000;
		4145: Delta = 39'sb000000000000000011111000000000000000000;
		11210: Delta = 39'sb111111111111111011111000000000000000000;
		6013: Delta = 39'sb000000000000001000001000000000000000000;
		6306: Delta = 39'sb111111111111111000001000000000000000000;
		7531: Delta = 39'sb000000000000000111111000000000000000000;
		7824: Delta = 39'sb111111111111110111111000000000000000000;
		12785: Delta = 39'sb000000000000010000001000000000000000000;
		13371: Delta = 39'sb111111111111110000001000000000000000000;
		466: Delta = 39'sb000000000000001111111000000000000000000;
		1052: Delta = 39'sb111111111111101111111000000000000000000;
		12492: Delta = 39'sb000000000000100000001000000000000000000;
		13664: Delta = 39'sb111111111111100000001000000000000000000;
		173: Delta = 39'sb000000000000011111111000000000000000000;
		1345: Delta = 39'sb111111111111011111111000000000000000000;
		11906: Delta = 39'sb000000000001000000001000000000000000000;
		413: Delta = 39'sb111111111111000000001000000000000000000;
		13424: Delta = 39'sb000000000000111111111000000000000000000;
		1931: Delta = 39'sb111111111110111111111000000000000000000;
		10734: Delta = 39'sb000000000010000000001000000000000000000;
		1585: Delta = 39'sb111111111110000000001000000000000000000;
		12252: Delta = 39'sb000000000001111111111000000000000000000;
		3103: Delta = 39'sb111111111101111111111000000000000000000;
		8390: Delta = 39'sb000000000100000000001000000000000000000;
		3929: Delta = 39'sb111111111100000000001000000000000000000;
		9908: Delta = 39'sb000000000011111111111000000000000000000;
		5447: Delta = 39'sb111111111011111111111000000000000000000;
		3702: Delta = 39'sb000000001000000000001000000000000000000;
		8617: Delta = 39'sb111111111000000000001000000000000000000;
		5220: Delta = 39'sb000000000111111111111000000000000000000;
		10135: Delta = 39'sb111111110111111111111000000000000000000;
		8163: Delta = 39'sb000000010000000000001000000000000000000;
		4156: Delta = 39'sb111111110000000000001000000000000000000;
		9681: Delta = 39'sb000000001111111111111000000000000000000;
		5674: Delta = 39'sb111111101111111111111000000000000000000;
		3248: Delta = 39'sb000000100000000000001000000000000000000;
		9071: Delta = 39'sb111111100000000000001000000000000000000;
		4766: Delta = 39'sb000000011111111111111000000000000000000;
		10589: Delta = 39'sb111111011111111111111000000000000000000;
		7255: Delta = 39'sb000001000000000000001000000000000000000;
		5064: Delta = 39'sb111111000000000000001000000000000000000;
		8773: Delta = 39'sb000000111111111111111000000000000000000;
		6582: Delta = 39'sb111110111111111111111000000000000000000;
		1432: Delta = 39'sb000010000000000000001000000000000000000;
		10887: Delta = 39'sb111110000000000000001000000000000000000;
		2950: Delta = 39'sb000001111111111111111000000000000000000;
		12405: Delta = 39'sb111101111111111111111000000000000000000;
		3623: Delta = 39'sb000100000000000000001000000000000000000;
		8696: Delta = 39'sb111100000000000000001000000000000000000;
		5141: Delta = 39'sb000011111111111111111000000000000000000;
		10214: Delta = 39'sb111011111111111111111000000000000000000;
		8005: Delta = 39'sb001000000000000000001000000000000000000;
		4314: Delta = 39'sb111000000000000000001000000000000000000;
		9523: Delta = 39'sb000111111111111111111000000000000000000;
		5832: Delta = 39'sb110111111111111111111000000000000000000;
		2932: Delta = 39'sb010000000000000000001000000000000000000;
		9387: Delta = 39'sb110000000000000000001000000000000000000;
		4450: Delta = 39'sb001111111111111111111000000000000000000;
		10905: Delta = 39'sb101111111111111111111000000000000000000;
		9283: Delta = 39'sb000000000000000000110000000000000000000;
		4554: Delta = 39'sb111111111111111111010000000000000000000;
		6247: Delta = 39'sb000000000000000001010000000000000000000;
		7590: Delta = 39'sb111111111111111110110000000000000000000;
		175: Delta = 39'sb000000000000000010010000000000000000000;
		10626: Delta = 39'sb111111111111111110010000000000000000000;
		3211: Delta = 39'sb000000000000000001110000000000000000000;
		13662: Delta = 39'sb111111111111111101110000000000000000000;
		1868: Delta = 39'sb000000000000000100010000000000000000000;
		8933: Delta = 39'sb111111111111111100010000000000000000000;
		4904: Delta = 39'sb000000000000000011110000000000000000000;
		11969: Delta = 39'sb111111111111111011110000000000000000000;
		5254: Delta = 39'sb000000000000001000010000000000000000000;
		5547: Delta = 39'sb111111111111111000010000000000000000000;
		8290: Delta = 39'sb000000000000000111110000000000000000000;
		8583: Delta = 39'sb111111111111110111110000000000000000000;
		12026: Delta = 39'sb000000000000010000010000000000000000000;
		12612: Delta = 39'sb111111111111110000010000000000000000000;
		1225: Delta = 39'sb000000000000001111110000000000000000000;
		1811: Delta = 39'sb111111111111101111110000000000000000000;
		11733: Delta = 39'sb000000000000100000010000000000000000000;
		12905: Delta = 39'sb111111111111100000010000000000000000000;
		932: Delta = 39'sb000000000000011111110000000000000000000;
		2104: Delta = 39'sb111111111111011111110000000000000000000;
		11147: Delta = 39'sb000000000001000000010000000000000000000;
		13491: Delta = 39'sb111111111111000000010000000000000000000;
		346: Delta = 39'sb000000000000111111110000000000000000000;
		2690: Delta = 39'sb111111111110111111110000000000000000000;
		9975: Delta = 39'sb000000000010000000010000000000000000000;
		826: Delta = 39'sb111111111110000000010000000000000000000;
		13011: Delta = 39'sb000000000001111111110000000000000000000;
		3862: Delta = 39'sb111111111101111111110000000000000000000;
		7631: Delta = 39'sb000000000100000000010000000000000000000;
		3170: Delta = 39'sb111111111100000000010000000000000000000;
		10667: Delta = 39'sb000000000011111111110000000000000000000;
		6206: Delta = 39'sb111111111011111111110000000000000000000;
		2943: Delta = 39'sb000000001000000000010000000000000000000;
		7858: Delta = 39'sb111111111000000000010000000000000000000;
		5979: Delta = 39'sb000000000111111111110000000000000000000;
		10894: Delta = 39'sb111111110111111111110000000000000000000;
		7404: Delta = 39'sb000000010000000000010000000000000000000;
		3397: Delta = 39'sb111111110000000000010000000000000000000;
		10440: Delta = 39'sb000000001111111111110000000000000000000;
		6433: Delta = 39'sb111111101111111111110000000000000000000;
		2489: Delta = 39'sb000000100000000000010000000000000000000;
		8312: Delta = 39'sb111111100000000000010000000000000000000;
		5525: Delta = 39'sb000000011111111111110000000000000000000;
		11348: Delta = 39'sb111111011111111111110000000000000000000;
		6496: Delta = 39'sb000001000000000000010000000000000000000;
		4305: Delta = 39'sb111111000000000000010000000000000000000;
		9532: Delta = 39'sb000000111111111111110000000000000000000;
		7341: Delta = 39'sb111110111111111111110000000000000000000;
		673: Delta = 39'sb000010000000000000010000000000000000000;
		10128: Delta = 39'sb111110000000000000010000000000000000000;
		3709: Delta = 39'sb000001111111111111110000000000000000000;
		13164: Delta = 39'sb111101111111111111110000000000000000000;
		2864: Delta = 39'sb000100000000000000010000000000000000000;
		7937: Delta = 39'sb111100000000000000010000000000000000000;
		5900: Delta = 39'sb000011111111111111110000000000000000000;
		10973: Delta = 39'sb111011111111111111110000000000000000000;
		7246: Delta = 39'sb001000000000000000010000000000000000000;
		3555: Delta = 39'sb111000000000000000010000000000000000000;
		10282: Delta = 39'sb000111111111111111110000000000000000000;
		6591: Delta = 39'sb110111111111111111110000000000000000000;
		2173: Delta = 39'sb010000000000000000010000000000000000000;
		8628: Delta = 39'sb110000000000000000010000000000000000000;
		5209: Delta = 39'sb001111111111111111110000000000000000000;
		11664: Delta = 39'sb101111111111111111110000000000000000000;
		4729: Delta = 39'sb000000000000000001100000000000000000000;
		9108: Delta = 39'sb111111111111111110100000000000000000000;
		12494: Delta = 39'sb000000000000000010100000000000000000000;
		1343: Delta = 39'sb111111111111111101100000000000000000000;
		350: Delta = 39'sb000000000000000100100000000000000000000;
		7415: Delta = 39'sb111111111111111100100000000000000000000;
		6422: Delta = 39'sb000000000000000011100000000000000000000;
		13487: Delta = 39'sb111111111111111011100000000000000000000;
		3736: Delta = 39'sb000000000000001000100000000000000000000;
		4029: Delta = 39'sb111111111111111000100000000000000000000;
		9808: Delta = 39'sb000000000000000111100000000000000000000;
		10101: Delta = 39'sb111111111111110111100000000000000000000;
		10508: Delta = 39'sb000000000000010000100000000000000000000;
		11094: Delta = 39'sb111111111111110000100000000000000000000;
		2743: Delta = 39'sb000000000000001111100000000000000000000;
		3329: Delta = 39'sb111111111111101111100000000000000000000;
		10215: Delta = 39'sb000000000000100000100000000000000000000;
		11387: Delta = 39'sb111111111111100000100000000000000000000;
		2450: Delta = 39'sb000000000000011111100000000000000000000;
		3622: Delta = 39'sb111111111111011111100000000000000000000;
		9629: Delta = 39'sb000000000001000000100000000000000000000;
		11973: Delta = 39'sb111111111111000000100000000000000000000;
		1864: Delta = 39'sb000000000000111111100000000000000000000;
		4208: Delta = 39'sb111111111110111111100000000000000000000;
		8457: Delta = 39'sb000000000010000000100000000000000000000;
		13145: Delta = 39'sb111111111110000000100000000000000000000;
		692: Delta = 39'sb000000000001111111100000000000000000000;
		5380: Delta = 39'sb111111111101111111100000000000000000000;
		6113: Delta = 39'sb000000000100000000100000000000000000000;
		1652: Delta = 39'sb111111111100000000100000000000000000000;
		12185: Delta = 39'sb000000000011111111100000000000000000000;
		7724: Delta = 39'sb111111111011111111100000000000000000000;
		1425: Delta = 39'sb000000001000000000100000000000000000000;
		6340: Delta = 39'sb111111111000000000100000000000000000000;
		7497: Delta = 39'sb000000000111111111100000000000000000000;
		12412: Delta = 39'sb111111110111111111100000000000000000000;
		5886: Delta = 39'sb000000010000000000100000000000000000000;
		1879: Delta = 39'sb111111110000000000100000000000000000000;
		11958: Delta = 39'sb000000001111111111100000000000000000000;
		7951: Delta = 39'sb111111101111111111100000000000000000000;
		971: Delta = 39'sb000000100000000000100000000000000000000;
		6794: Delta = 39'sb111111100000000000100000000000000000000;
		7043: Delta = 39'sb000000011111111111100000000000000000000;
		12866: Delta = 39'sb111111011111111111100000000000000000000;
		4978: Delta = 39'sb000001000000000000100000000000000000000;
		2787: Delta = 39'sb111111000000000000100000000000000000000;
		11050: Delta = 39'sb000000111111111111100000000000000000000;
		8859: Delta = 39'sb111110111111111111100000000000000000000;
		12992: Delta = 39'sb000010000000000000100000000000000000000;
		8610: Delta = 39'sb111110000000000000100000000000000000000;
		5227: Delta = 39'sb000001111111111111100000000000000000000;
		845: Delta = 39'sb111101111111111111100000000000000000000;
		1346: Delta = 39'sb000100000000000000100000000000000000000;
		6419: Delta = 39'sb111100000000000000100000000000000000000;
		7418: Delta = 39'sb000011111111111111100000000000000000000;
		12491: Delta = 39'sb111011111111111111100000000000000000000;
		5728: Delta = 39'sb001000000000000000100000000000000000000;
		2037: Delta = 39'sb111000000000000000100000000000000000000;
		11800: Delta = 39'sb000111111111111111100000000000000000000;
		8109: Delta = 39'sb110111111111111111100000000000000000000;
		655: Delta = 39'sb010000000000000000100000000000000000000;
		7110: Delta = 39'sb110000000000000000100000000000000000000;
		6727: Delta = 39'sb001111111111111111100000000000000000000;
		13182: Delta = 39'sb101111111111111111100000000000000000000;
		9458: Delta = 39'sb000000000000000011000000000000000000000;
		4379: Delta = 39'sb111111111111111101000000000000000000000;
		11151: Delta = 39'sb000000000000000101000000000000000000000;
		2686: Delta = 39'sb111111111111111011000000000000000000000;
		700: Delta = 39'sb000000000000001001000000000000000000000;
		993: Delta = 39'sb111111111111111001000000000000000000000;
		12844: Delta = 39'sb000000000000000111000000000000000000000;
		13137: Delta = 39'sb111111111111110111000000000000000000000;
		7472: Delta = 39'sb000000000000010001000000000000000000000;
		8058: Delta = 39'sb111111111111110001000000000000000000000;
		5779: Delta = 39'sb000000000000001111000000000000000000000;
		6365: Delta = 39'sb111111111111101111000000000000000000000;
		7179: Delta = 39'sb000000000000100001000000000000000000000;
		8351: Delta = 39'sb111111111111100001000000000000000000000;
		5486: Delta = 39'sb000000000000011111000000000000000000000;
		6658: Delta = 39'sb111111111111011111000000000000000000000;
		6593: Delta = 39'sb000000000001000001000000000000000000000;
		8937: Delta = 39'sb111111111111000001000000000000000000000;
		4900: Delta = 39'sb000000000000111111000000000000000000000;
		7244: Delta = 39'sb111111111110111111000000000000000000000;
		5421: Delta = 39'sb000000000010000001000000000000000000000;
		10109: Delta = 39'sb111111111110000001000000000000000000000;
		3728: Delta = 39'sb000000000001111111000000000000000000000;
		8416: Delta = 39'sb111111111101111111000000000000000000000;
		3077: Delta = 39'sb000000000100000001000000000000000000000;
		12453: Delta = 39'sb111111111100000001000000000000000000000;
		1384: Delta = 39'sb000000000011111111000000000000000000000;
		10760: Delta = 39'sb111111111011111111000000000000000000000;
		12226: Delta = 39'sb000000001000000001000000000000000000000;
		3304: Delta = 39'sb111111111000000001000000000000000000000;
		10533: Delta = 39'sb000000000111111111000000000000000000000;
		1611: Delta = 39'sb111111110111111111000000000000000000000;
		2850: Delta = 39'sb000000010000000001000000000000000000000;
		12680: Delta = 39'sb111111110000000001000000000000000000000;
		1157: Delta = 39'sb000000001111111111000000000000000000000;
		10987: Delta = 39'sb111111101111111111000000000000000000000;
		11772: Delta = 39'sb000000100000000001000000000000000000000;
		3758: Delta = 39'sb111111100000000001000000000000000000000;
		10079: Delta = 39'sb000000011111111111000000000000000000000;
		2065: Delta = 39'sb111111011111111111000000000000000000000;
		1942: Delta = 39'sb000001000000000001000000000000000000000;
		13588: Delta = 39'sb111111000000000001000000000000000000000;
		249: Delta = 39'sb000000111111111111000000000000000000000;
		11895: Delta = 39'sb111110111111111111000000000000000000000;
		9956: Delta = 39'sb000010000000000001000000000000000000000;
		5574: Delta = 39'sb111110000000000001000000000000000000000;
		8263: Delta = 39'sb000001111111111111000000000000000000000;
		3881: Delta = 39'sb111101111111111111000000000000000000000;
		12147: Delta = 39'sb000100000000000001000000000000000000000;
		3383: Delta = 39'sb111100000000000001000000000000000000000;
		10454: Delta = 39'sb000011111111111111000000000000000000000;
		1690: Delta = 39'sb111011111111111111000000000000000000000;
		2692: Delta = 39'sb001000000000000001000000000000000000000;
		12838: Delta = 39'sb111000000000000001000000000000000000000;
		999: Delta = 39'sb000111111111111111000000000000000000000;
		11145: Delta = 39'sb110111111111111111000000000000000000000;
		11456: Delta = 39'sb010000000000000001000000000000000000000;
		4074: Delta = 39'sb110000000000000001000000000000000000000;
		9763: Delta = 39'sb001111111111111111000000000000000000000;
		2381: Delta = 39'sb101111111111111111000000000000000000000;
		5079: Delta = 39'sb000000000000000110000000000000000000000;
		8758: Delta = 39'sb111111111111111010000000000000000000000;
		8465: Delta = 39'sb000000000000001010000000000000000000000;
		5372: Delta = 39'sb111111111111110110000000000000000000000;
		1400: Delta = 39'sb000000000000010010000000000000000000000;
		1986: Delta = 39'sb111111111111110010000000000000000000000;
		11851: Delta = 39'sb000000000000001110000000000000000000000;
		12437: Delta = 39'sb111111111111101110000000000000000000000;
		1107: Delta = 39'sb000000000000100010000000000000000000000;
		2279: Delta = 39'sb111111111111100010000000000000000000000;
		11558: Delta = 39'sb000000000000011110000000000000000000000;
		12730: Delta = 39'sb111111111111011110000000000000000000000;
		521: Delta = 39'sb000000000001000010000000000000000000000;
		2865: Delta = 39'sb111111111111000010000000000000000000000;
		10972: Delta = 39'sb000000000000111110000000000000000000000;
		13316: Delta = 39'sb111111111110111110000000000000000000000;
		13186: Delta = 39'sb000000000010000010000000000000000000000;
		4037: Delta = 39'sb111111111110000010000000000000000000000;
		9800: Delta = 39'sb000000000001111110000000000000000000000;
		651: Delta = 39'sb111111111101111110000000000000000000000;
		10842: Delta = 39'sb000000000100000010000000000000000000000;
		6381: Delta = 39'sb111111111100000010000000000000000000000;
		7456: Delta = 39'sb000000000011111110000000000000000000000;
		2995: Delta = 39'sb111111111011111110000000000000000000000;
		6154: Delta = 39'sb000000001000000010000000000000000000000;
		11069: Delta = 39'sb111111111000000010000000000000000000000;
		2768: Delta = 39'sb000000000111111110000000000000000000000;
		7683: Delta = 39'sb111111110111111110000000000000000000000;
		10615: Delta = 39'sb000000010000000010000000000000000000000;
		6608: Delta = 39'sb111111110000000010000000000000000000000;
		7229: Delta = 39'sb000000001111111110000000000000000000000;
		3222: Delta = 39'sb111111101111111110000000000000000000000;
		5700: Delta = 39'sb000000100000000010000000000000000000000;
		11523: Delta = 39'sb111111100000000010000000000000000000000;
		2314: Delta = 39'sb000000011111111110000000000000000000000;
		8137: Delta = 39'sb111111011111111110000000000000000000000;
		9707: Delta = 39'sb000001000000000010000000000000000000000;
		7516: Delta = 39'sb111111000000000010000000000000000000000;
		6321: Delta = 39'sb000000111111111110000000000000000000000;
		4130: Delta = 39'sb111110111111111110000000000000000000000;
		3884: Delta = 39'sb000010000000000010000000000000000000000;
		13339: Delta = 39'sb111110000000000010000000000000000000000;
		498: Delta = 39'sb000001111111111110000000000000000000000;
		9953: Delta = 39'sb111101111111111110000000000000000000000;
		6075: Delta = 39'sb000100000000000010000000000000000000000;
		11148: Delta = 39'sb111100000000000010000000000000000000000;
		2689: Delta = 39'sb000011111111111110000000000000000000000;
		7762: Delta = 39'sb111011111111111110000000000000000000000;
		10457: Delta = 39'sb001000000000000010000000000000000000000;
		6766: Delta = 39'sb111000000000000010000000000000000000000;
		7071: Delta = 39'sb000111111111111110000000000000000000000;
		3380: Delta = 39'sb110111111111111110000000000000000000000;
		5384: Delta = 39'sb010000000000000010000000000000000000000;
		11839: Delta = 39'sb110000000000000010000000000000000000000;
		1998: Delta = 39'sb001111111111111110000000000000000000000;
		8453: Delta = 39'sb101111111111111110000000000000000000000;
		10158: Delta = 39'sb000000000000001100000000000000000000000;
		3679: Delta = 39'sb111111111111110100000000000000000000000;
		3093: Delta = 39'sb000000000000010100000000000000000000000;
		10744: Delta = 39'sb111111111111101100000000000000000000000;
		2800: Delta = 39'sb000000000000100100000000000000000000000;
		3972: Delta = 39'sb111111111111100100000000000000000000000;
		9865: Delta = 39'sb000000000000011100000000000000000000000;
		11037: Delta = 39'sb111111111111011100000000000000000000000;
		2214: Delta = 39'sb000000000001000100000000000000000000000;
		4558: Delta = 39'sb111111111111000100000000000000000000000;
		9279: Delta = 39'sb000000000000111100000000000000000000000;
		11623: Delta = 39'sb111111111110111100000000000000000000000;
		1042: Delta = 39'sb000000000010000100000000000000000000000;
		5730: Delta = 39'sb111111111110000100000000000000000000000;
		8107: Delta = 39'sb000000000001111100000000000000000000000;
		12795: Delta = 39'sb111111111101111100000000000000000000000;
		12535: Delta = 39'sb000000000100000100000000000000000000000;
		8074: Delta = 39'sb111111111100000100000000000000000000000;
		5763: Delta = 39'sb000000000011111100000000000000000000000;
		1302: Delta = 39'sb111111111011111100000000000000000000000;
		7847: Delta = 39'sb000000001000000100000000000000000000000;
		12762: Delta = 39'sb111111111000000100000000000000000000000;
		1075: Delta = 39'sb000000000111111100000000000000000000000;
		5990: Delta = 39'sb111111110111111100000000000000000000000;
		12308: Delta = 39'sb000000010000000100000000000000000000000;
		8301: Delta = 39'sb111111110000000100000000000000000000000;
		5536: Delta = 39'sb000000001111111100000000000000000000000;
		1529: Delta = 39'sb111111101111111100000000000000000000000;
		7393: Delta = 39'sb000000100000000100000000000000000000000;
		13216: Delta = 39'sb111111100000000100000000000000000000000;
		621: Delta = 39'sb000000011111111100000000000000000000000;
		6444: Delta = 39'sb111111011111111100000000000000000000000;
		11400: Delta = 39'sb000001000000000100000000000000000000000;
		9209: Delta = 39'sb111111000000000100000000000000000000000;
		4628: Delta = 39'sb000000111111111100000000000000000000000;
		2437: Delta = 39'sb111110111111111100000000000000000000000;
		5577: Delta = 39'sb000010000000000100000000000000000000000;
		1195: Delta = 39'sb111110000000000100000000000000000000000;
		12642: Delta = 39'sb000001111111111100000000000000000000000;
		8260: Delta = 39'sb111101111111111100000000000000000000000;
		7768: Delta = 39'sb000100000000000100000000000000000000000;
		12841: Delta = 39'sb111100000000000100000000000000000000000;
		996: Delta = 39'sb000011111111111100000000000000000000000;
		6069: Delta = 39'sb111011111111111100000000000000000000000;
		12150: Delta = 39'sb001000000000000100000000000000000000000;
		8459: Delta = 39'sb111000000000000100000000000000000000000;
		5378: Delta = 39'sb000111111111111100000000000000000000000;
		1687: Delta = 39'sb110111111111111100000000000000000000000;
		7077: Delta = 39'sb010000000000000100000000000000000000000;
		13532: Delta = 39'sb110000000000000100000000000000000000000;
		305: Delta = 39'sb001111111111111100000000000000000000000;
		6760: Delta = 39'sb101111111111111100000000000000000000000;
		6479: Delta = 39'sb000000000000011000000000000000000000000;
		7358: Delta = 39'sb111111111111101000000000000000000000000;
		6186: Delta = 39'sb000000000000101000000000000000000000000;
		7651: Delta = 39'sb111111111111011000000000000000000000000;
		5600: Delta = 39'sb000000000001001000000000000000000000000;
		7944: Delta = 39'sb111111111111001000000000000000000000000;
		5893: Delta = 39'sb000000000000111000000000000000000000000;
		8237: Delta = 39'sb111111111110111000000000000000000000000;
		4428: Delta = 39'sb000000000010001000000000000000000000000;
		9116: Delta = 39'sb111111111110001000000000000000000000000;
		4721: Delta = 39'sb000000000001111000000000000000000000000;
		9409: Delta = 39'sb111111111101111000000000000000000000000;
		2084: Delta = 39'sb000000000100001000000000000000000000000;
		11460: Delta = 39'sb111111111100001000000000000000000000000;
		2377: Delta = 39'sb000000000011111000000000000000000000000;
		11753: Delta = 39'sb111111111011111000000000000000000000000;
		11233: Delta = 39'sb000000001000001000000000000000000000000;
		2311: Delta = 39'sb111111111000001000000000000000000000000;
		11526: Delta = 39'sb000000000111111000000000000000000000000;
		2604: Delta = 39'sb111111110111111000000000000000000000000;
		1857: Delta = 39'sb000000010000001000000000000000000000000;
		11687: Delta = 39'sb111111110000001000000000000000000000000;
		2150: Delta = 39'sb000000001111111000000000000000000000000;
		11980: Delta = 39'sb111111101111111000000000000000000000000;
		10779: Delta = 39'sb000000100000001000000000000000000000000;
		2765: Delta = 39'sb111111100000001000000000000000000000000;
		11072: Delta = 39'sb000000011111111000000000000000000000000;
		3058: Delta = 39'sb111111011111111000000000000000000000000;
		949: Delta = 39'sb000001000000001000000000000000000000000;
		12595: Delta = 39'sb111111000000001000000000000000000000000;
		1242: Delta = 39'sb000000111111111000000000000000000000000;
		12888: Delta = 39'sb111110111111111000000000000000000000000;
		8963: Delta = 39'sb000010000000001000000000000000000000000;
		4581: Delta = 39'sb111110000000001000000000000000000000000;
		9256: Delta = 39'sb000001111111111000000000000000000000000;
		4874: Delta = 39'sb111101111111111000000000000000000000000;
		11154: Delta = 39'sb000100000000001000000000000000000000000;
		2390: Delta = 39'sb111100000000001000000000000000000000000;
		11447: Delta = 39'sb000011111111111000000000000000000000000;
		2683: Delta = 39'sb111011111111111000000000000000000000000;
		1699: Delta = 39'sb001000000000001000000000000000000000000;
		11845: Delta = 39'sb111000000000001000000000000000000000000;
		1992: Delta = 39'sb000111111111111000000000000000000000000;
		12138: Delta = 39'sb110111111111111000000000000000000000000;
		10463: Delta = 39'sb010000000000001000000000000000000000000;
		3081: Delta = 39'sb110000000000001000000000000000000000000;
		10756: Delta = 39'sb001111111111111000000000000000000000000;
		3374: Delta = 39'sb101111111111111000000000000000000000000;
		12958: Delta = 39'sb000000000000110000000000000000000000000;
		879: Delta = 39'sb111111111111010000000000000000000000000;
		12372: Delta = 39'sb000000000001010000000000000000000000000;
		1465: Delta = 39'sb111111111110110000000000000000000000000;
		11200: Delta = 39'sb000000000010010000000000000000000000000;
		2051: Delta = 39'sb111111111110010000000000000000000000000;
		11786: Delta = 39'sb000000000001110000000000000000000000000;
		2637: Delta = 39'sb111111111101110000000000000000000000000;
		8856: Delta = 39'sb000000000100010000000000000000000000000;
		4395: Delta = 39'sb111111111100010000000000000000000000000;
		9442: Delta = 39'sb000000000011110000000000000000000000000;
		4981: Delta = 39'sb111111111011110000000000000000000000000;
		4168: Delta = 39'sb000000001000010000000000000000000000000;
		9083: Delta = 39'sb111111111000010000000000000000000000000;
		4754: Delta = 39'sb000000000111110000000000000000000000000;
		9669: Delta = 39'sb111111110111110000000000000000000000000;
		8629: Delta = 39'sb000000010000010000000000000000000000000;
		4622: Delta = 39'sb111111110000010000000000000000000000000;
		9215: Delta = 39'sb000000001111110000000000000000000000000;
		5208: Delta = 39'sb111111101111110000000000000000000000000;
		3714: Delta = 39'sb000000100000010000000000000000000000000;
		9537: Delta = 39'sb111111100000010000000000000000000000000;
		4300: Delta = 39'sb000000011111110000000000000000000000000;
		10123: Delta = 39'sb111111011111110000000000000000000000000;
		7721: Delta = 39'sb000001000000010000000000000000000000000;
		5530: Delta = 39'sb111111000000010000000000000000000000000;
		8307: Delta = 39'sb000000111111110000000000000000000000000;
		6116: Delta = 39'sb111110111111110000000000000000000000000;
		1898: Delta = 39'sb000010000000010000000000000000000000000;
		11353: Delta = 39'sb111110000000010000000000000000000000000;
		2484: Delta = 39'sb000001111111110000000000000000000000000;
		11939: Delta = 39'sb111101111111110000000000000000000000000;
		4089: Delta = 39'sb000100000000010000000000000000000000000;
		9162: Delta = 39'sb111100000000010000000000000000000000000;
		4675: Delta = 39'sb000011111111110000000000000000000000000;
		9748: Delta = 39'sb111011111111110000000000000000000000000;
		8471: Delta = 39'sb001000000000010000000000000000000000000;
		4780: Delta = 39'sb111000000000010000000000000000000000000;
		9057: Delta = 39'sb000111111111110000000000000000000000000;
		5366: Delta = 39'sb110111111111110000000000000000000000000;
		3398: Delta = 39'sb010000000000010000000000000000000000000;
		9853: Delta = 39'sb110000000000010000000000000000000000000;
		3984: Delta = 39'sb001111111111110000000000000000000000000;
		10439: Delta = 39'sb101111111111110000000000000000000000000;
		12079: Delta = 39'sb000000000001100000000000000000000000000;
		1758: Delta = 39'sb111111111110100000000000000000000000000;
		10907: Delta = 39'sb000000000010100000000000000000000000000;
		2930: Delta = 39'sb111111111101100000000000000000000000000;
		8563: Delta = 39'sb000000000100100000000000000000000000000;
		4102: Delta = 39'sb111111111100100000000000000000000000000;
		9735: Delta = 39'sb000000000011100000000000000000000000000;
		5274: Delta = 39'sb111111111011100000000000000000000000000;
		3875: Delta = 39'sb000000001000100000000000000000000000000;
		8790: Delta = 39'sb111111111000100000000000000000000000000;
		5047: Delta = 39'sb000000000111100000000000000000000000000;
		9962: Delta = 39'sb111111110111100000000000000000000000000;
		8336: Delta = 39'sb000000010000100000000000000000000000000;
		4329: Delta = 39'sb111111110000100000000000000000000000000;
		9508: Delta = 39'sb000000001111100000000000000000000000000;
		5501: Delta = 39'sb111111101111100000000000000000000000000;
		3421: Delta = 39'sb000000100000100000000000000000000000000;
		9244: Delta = 39'sb111111100000100000000000000000000000000;
		4593: Delta = 39'sb000000011111100000000000000000000000000;
		10416: Delta = 39'sb111111011111100000000000000000000000000;
		7428: Delta = 39'sb000001000000100000000000000000000000000;
		5237: Delta = 39'sb111111000000100000000000000000000000000;
		8600: Delta = 39'sb000000111111100000000000000000000000000;
		6409: Delta = 39'sb111110111111100000000000000000000000000;
		1605: Delta = 39'sb000010000000100000000000000000000000000;
		11060: Delta = 39'sb111110000000100000000000000000000000000;
		2777: Delta = 39'sb000001111111100000000000000000000000000;
		12232: Delta = 39'sb111101111111100000000000000000000000000;
		3796: Delta = 39'sb000100000000100000000000000000000000000;
		8869: Delta = 39'sb111100000000100000000000000000000000000;
		4968: Delta = 39'sb000011111111100000000000000000000000000;
		10041: Delta = 39'sb111011111111100000000000000000000000000;
		8178: Delta = 39'sb001000000000100000000000000000000000000;
		4487: Delta = 39'sb111000000000100000000000000000000000000;
		9350: Delta = 39'sb000111111111100000000000000000000000000;
		5659: Delta = 39'sb110111111111100000000000000000000000000;
		3105: Delta = 39'sb010000000000100000000000000000000000000;
		9560: Delta = 39'sb110000000000100000000000000000000000000;
		4277: Delta = 39'sb001111111111100000000000000000000000000;
		10732: Delta = 39'sb101111111111100000000000000000000000000;
		10321: Delta = 39'sb000000000011000000000000000000000000000;
		3516: Delta = 39'sb111111111101000000000000000000000000000;
		7977: Delta = 39'sb000000000101000000000000000000000000000;
		5860: Delta = 39'sb111111111011000000000000000000000000000;
		3289: Delta = 39'sb000000001001000000000000000000000000000;
		8204: Delta = 39'sb111111111001000000000000000000000000000;
		5633: Delta = 39'sb000000000111000000000000000000000000000;
		10548: Delta = 39'sb111111110111000000000000000000000000000;
		7750: Delta = 39'sb000000010001000000000000000000000000000;
		3743: Delta = 39'sb111111110001000000000000000000000000000;
		10094: Delta = 39'sb000000001111000000000000000000000000000;
		6087: Delta = 39'sb111111101111000000000000000000000000000;
		2835: Delta = 39'sb000000100001000000000000000000000000000;
		8658: Delta = 39'sb111111100001000000000000000000000000000;
		5179: Delta = 39'sb000000011111000000000000000000000000000;
		11002: Delta = 39'sb111111011111000000000000000000000000000;
		6842: Delta = 39'sb000001000001000000000000000000000000000;
		4651: Delta = 39'sb111111000001000000000000000000000000000;
		9186: Delta = 39'sb000000111111000000000000000000000000000;
		6995: Delta = 39'sb111110111111000000000000000000000000000;
		1019: Delta = 39'sb000010000001000000000000000000000000000;
		10474: Delta = 39'sb111110000001000000000000000000000000000;
		3363: Delta = 39'sb000001111111000000000000000000000000000;
		12818: Delta = 39'sb111101111111000000000000000000000000000;
		3210: Delta = 39'sb000100000001000000000000000000000000000;
		8283: Delta = 39'sb111100000001000000000000000000000000000;
		5554: Delta = 39'sb000011111111000000000000000000000000000;
		10627: Delta = 39'sb111011111111000000000000000000000000000;
		7592: Delta = 39'sb001000000001000000000000000000000000000;
		3901: Delta = 39'sb111000000001000000000000000000000000000;
		9936: Delta = 39'sb000111111111000000000000000000000000000;
		6245: Delta = 39'sb110111111111000000000000000000000000000;
		2519: Delta = 39'sb010000000001000000000000000000000000000;
		8974: Delta = 39'sb110000000001000000000000000000000000000;
		4863: Delta = 39'sb001111111111000000000000000000000000000;
		11318: Delta = 39'sb101111111111000000000000000000000000000;
		6805: Delta = 39'sb000000000110000000000000000000000000000;
		7032: Delta = 39'sb111111111010000000000000000000000000000;
		2117: Delta = 39'sb000000001010000000000000000000000000000;
		11720: Delta = 39'sb111111110110000000000000000000000000000;
		6578: Delta = 39'sb000000010010000000000000000000000000000;
		2571: Delta = 39'sb111111110010000000000000000000000000000;
		11266: Delta = 39'sb000000001110000000000000000000000000000;
		7259: Delta = 39'sb111111101110000000000000000000000000000;
		1663: Delta = 39'sb000000100010000000000000000000000000000;
		7486: Delta = 39'sb111111100010000000000000000000000000000;
		6351: Delta = 39'sb000000011110000000000000000000000000000;
		12174: Delta = 39'sb111111011110000000000000000000000000000;
		5670: Delta = 39'sb000001000010000000000000000000000000000;
		3479: Delta = 39'sb111111000010000000000000000000000000000;
		10358: Delta = 39'sb000000111110000000000000000000000000000;
		8167: Delta = 39'sb111110111110000000000000000000000000000;
		13684: Delta = 39'sb000010000010000000000000000000000000000;
		9302: Delta = 39'sb111110000010000000000000000000000000000;
		4535: Delta = 39'sb000001111110000000000000000000000000000;
		153: Delta = 39'sb111101111110000000000000000000000000000;
		2038: Delta = 39'sb000100000010000000000000000000000000000;
		7111: Delta = 39'sb111100000010000000000000000000000000000;
		6726: Delta = 39'sb000011111110000000000000000000000000000;
		11799: Delta = 39'sb111011111110000000000000000000000000000;
		6420: Delta = 39'sb001000000010000000000000000000000000000;
		2729: Delta = 39'sb111000000010000000000000000000000000000;
		11108: Delta = 39'sb000111111110000000000000000000000000000;
		7417: Delta = 39'sb110111111110000000000000000000000000000;
		1347: Delta = 39'sb010000000010000000000000000000000000000;
		7802: Delta = 39'sb110000000010000000000000000000000000000;
		6035: Delta = 39'sb001111111110000000000000000000000000000;
		12490: Delta = 39'sb101111111110000000000000000000000000000;
		13610: Delta = 39'sb000000001100000000000000000000000000000;
		227: Delta = 39'sb111111110100000000000000000000000000000;
		4234: Delta = 39'sb000000010100000000000000000000000000000;
		9603: Delta = 39'sb111111101100000000000000000000000000000;
		13156: Delta = 39'sb000000100100000000000000000000000000000;
		5142: Delta = 39'sb111111100100000000000000000000000000000;
		8695: Delta = 39'sb000000011100000000000000000000000000000;
		681: Delta = 39'sb111111011100000000000000000000000000000;
		3326: Delta = 39'sb000001000100000000000000000000000000000;
		1135: Delta = 39'sb111111000100000000000000000000000000000;
		12702: Delta = 39'sb000000111100000000000000000000000000000;
		10511: Delta = 39'sb111110111100000000000000000000000000000;
		11340: Delta = 39'sb000010000100000000000000000000000000000;
		6958: Delta = 39'sb111110000100000000000000000000000000000;
		6879: Delta = 39'sb000001111100000000000000000000000000000;
		2497: Delta = 39'sb111101111100000000000000000000000000000;
		13531: Delta = 39'sb000100000100000000000000000000000000000;
		4767: Delta = 39'sb111100000100000000000000000000000000000;
		9070: Delta = 39'sb000011111100000000000000000000000000000;
		306: Delta = 39'sb111011111100000000000000000000000000000;
		4076: Delta = 39'sb001000000100000000000000000000000000000;
		385: Delta = 39'sb111000000100000000000000000000000000000;
		13452: Delta = 39'sb000111111100000000000000000000000000000;
		9761: Delta = 39'sb110111111100000000000000000000000000000;
		12840: Delta = 39'sb010000000100000000000000000000000000000;
		5458: Delta = 39'sb110000000100000000000000000000000000000;
		8379: Delta = 39'sb001111111100000000000000000000000000000;
		997: Delta = 39'sb101111111100000000000000000000000000000;
		13383: Delta = 39'sb000000011000000000000000000000000000000;
		454: Delta = 39'sb111111101000000000000000000000000000000;
		8468: Delta = 39'sb000000101000000000000000000000000000000;
		5369: Delta = 39'sb111111011000000000000000000000000000000;
		12475: Delta = 39'sb000001001000000000000000000000000000000;
		10284: Delta = 39'sb111111001000000000000000000000000000000;
		3553: Delta = 39'sb000000111000000000000000000000000000000;
		1362: Delta = 39'sb111110111000000000000000000000000000000;
		6652: Delta = 39'sb000010001000000000000000000000000000000;
		2270: Delta = 39'sb111110001000000000000000000000000000000;
		11567: Delta = 39'sb000001111000000000000000000000000000000;
		7185: Delta = 39'sb111101111000000000000000000000000000000;
		8843: Delta = 39'sb000100001000000000000000000000000000000;
		79: Delta = 39'sb111100001000000000000000000000000000000;
		13758: Delta = 39'sb000011111000000000000000000000000000000;
		4994: Delta = 39'sb111011111000000000000000000000000000000;
		13225: Delta = 39'sb001000001000000000000000000000000000000;
		9534: Delta = 39'sb111000001000000000000000000000000000000;
		4303: Delta = 39'sb000111111000000000000000000000000000000;
		612: Delta = 39'sb110111111000000000000000000000000000000;
		8152: Delta = 39'sb010000001000000000000000000000000000000;
		770: Delta = 39'sb110000001000000000000000000000000000000;
		13067: Delta = 39'sb001111111000000000000000000000000000000;
		5685: Delta = 39'sb101111111000000000000000000000000000000;
		12929: Delta = 39'sb000000110000000000000000000000000000000;
		908: Delta = 39'sb111111010000000000000000000000000000000;
		3099: Delta = 39'sb000001010000000000000000000000000000000;
		10738: Delta = 39'sb111110110000000000000000000000000000000;
		11113: Delta = 39'sb000010010000000000000000000000000000000;
		6731: Delta = 39'sb111110010000000000000000000000000000000;
		7106: Delta = 39'sb000001110000000000000000000000000000000;
		2724: Delta = 39'sb111101110000000000000000000000000000000;
		13304: Delta = 39'sb000100010000000000000000000000000000000;
		4540: Delta = 39'sb111100010000000000000000000000000000000;
		9297: Delta = 39'sb000011110000000000000000000000000000000;
		533: Delta = 39'sb111011110000000000000000000000000000000;
		3849: Delta = 39'sb001000010000000000000000000000000000000;
		158: Delta = 39'sb111000010000000000000000000000000000000;
		13679: Delta = 39'sb000111110000000000000000000000000000000;
		9988: Delta = 39'sb110111110000000000000000000000000000000;
		12613: Delta = 39'sb010000010000000000000000000000000000000;
		5231: Delta = 39'sb110000010000000000000000000000000000000;
		8606: Delta = 39'sb001111110000000000000000000000000000000;
		1224: Delta = 39'sb101111110000000000000000000000000000000;
		12021: Delta = 39'sb000001100000000000000000000000000000000;
		1816: Delta = 39'sb111110100000000000000000000000000000000;
		6198: Delta = 39'sb000010100000000000000000000000000000000;
		7639: Delta = 39'sb111101100000000000000000000000000000000;
		8389: Delta = 39'sb000100100000000000000000000000000000000;
		13462: Delta = 39'sb111100100000000000000000000000000000000;
		375: Delta = 39'sb000011100000000000000000000000000000000;
		5448: Delta = 39'sb111011100000000000000000000000000000000;
		12771: Delta = 39'sb001000100000000000000000000000000000000;
		9080: Delta = 39'sb111000100000000000000000000000000000000;
		4757: Delta = 39'sb000111100000000000000000000000000000000;
		1066: Delta = 39'sb110111100000000000000000000000000000000;
		7698: Delta = 39'sb010000100000000000000000000000000000000;
		316: Delta = 39'sb110000100000000000000000000000000000000;
		13521: Delta = 39'sb001111100000000000000000000000000000000;
		6139: Delta = 39'sb101111100000000000000000000000000000000;
		10205: Delta = 39'sb000011000000000000000000000000000000000;
		3632: Delta = 39'sb111101000000000000000000000000000000000;
		12396: Delta = 39'sb000101000000000000000000000000000000000;
		1441: Delta = 39'sb111011000000000000000000000000000000000;
		2941: Delta = 39'sb001001000000000000000000000000000000000;
		13087: Delta = 39'sb111001000000000000000000000000000000000;
		750: Delta = 39'sb000111000000000000000000000000000000000;
		10896: Delta = 39'sb110111000000000000000000000000000000000;
		11705: Delta = 39'sb010001000000000000000000000000000000000;
		4323: Delta = 39'sb110001000000000000000000000000000000000;
		9514: Delta = 39'sb001111000000000000000000000000000000000;
		2132: Delta = 39'sb101111000000000000000000000000000000000;
		6573: Delta = 39'sb000110000000000000000000000000000000000;
		7264: Delta = 39'sb111010000000000000000000000000000000000;
		10955: Delta = 39'sb001010000000000000000000000000000000000;
		2882: Delta = 39'sb110110000000000000000000000000000000000;
		5882: Delta = 39'sb010010000000000000000000000000000000000;
		12337: Delta = 39'sb110010000000000000000000000000000000000;
		1500: Delta = 39'sb001110000000000000000000000000000000000;
		7955: Delta = 39'sb101110000000000000000000000000000000000;
		13146: Delta = 39'sb001100000000000000000000000000000000000;
		691: Delta = 39'sb110100000000000000000000000000000000000;
		8073: Delta = 39'sb010100000000000000000000000000000000000;
		5764: Delta = 39'sb101100000000000000000000000000000000000;
		12455: Delta = 39'sb011000000000000000000000000000000000000;
		1382: Delta = 39'sb101000000000000000000000000000000000000;
		default: Delta =39'sb0;
	endcase
end

assign N = (W - Delta) / A;

endmodule

// Product (AN) Code SEC_LUT_Decoder
// SEC_LUT_Decoder20bits.v
// Received codeword W = AN + e, e is single arithmetic weight error (AWE), +2^i or -2^i.
module SEC_LUT_Decoder20bits(W, N);
input 	[32:0]	W;
output	[19:0]	N;
parameter A = 6311;

wire 	[19:0]	Q;
wire 	[12:0]	R;
assign Q = W / A;
assign R = W - (A * Q);

reg	signed	[33:0]	Delta;
always@(*) begin
	case(R)
		1: Delta = 34'sb0000000000000000000000000000000001;
		6310: Delta = 34'sb1111111111111111111111111111111111;
		2: Delta = 34'sb0000000000000000000000000000000010;
		6309: Delta = 34'sb1111111111111111111111111111111110;
		4: Delta = 34'sb0000000000000000000000000000000100;
		6307: Delta = 34'sb1111111111111111111111111111111100;
		8: Delta = 34'sb0000000000000000000000000000001000;
		6303: Delta = 34'sb1111111111111111111111111111111000;
		16: Delta = 34'sb0000000000000000000000000000010000;
		6295: Delta = 34'sb1111111111111111111111111111110000;
		32: Delta = 34'sb0000000000000000000000000000100000;
		6279: Delta = 34'sb1111111111111111111111111111100000;
		64: Delta = 34'sb0000000000000000000000000001000000;
		6247: Delta = 34'sb1111111111111111111111111111000000;
		128: Delta = 34'sb0000000000000000000000000010000000;
		6183: Delta = 34'sb1111111111111111111111111110000000;
		256: Delta = 34'sb0000000000000000000000000100000000;
		6055: Delta = 34'sb1111111111111111111111111100000000;
		512: Delta = 34'sb0000000000000000000000001000000000;
		5799: Delta = 34'sb1111111111111111111111111000000000;
		1024: Delta = 34'sb0000000000000000000000010000000000;
		5287: Delta = 34'sb1111111111111111111111110000000000;
		2048: Delta = 34'sb0000000000000000000000100000000000;
		4263: Delta = 34'sb1111111111111111111111100000000000;
		4096: Delta = 34'sb0000000000000000000001000000000000;
		2215: Delta = 34'sb1111111111111111111111000000000000;
		1881: Delta = 34'sb0000000000000000000010000000000000;
		4430: Delta = 34'sb1111111111111111111110000000000000;
		3762: Delta = 34'sb0000000000000000000100000000000000;
		2549: Delta = 34'sb1111111111111111111100000000000000;
		1213: Delta = 34'sb0000000000000000001000000000000000;
		5098: Delta = 34'sb1111111111111111111000000000000000;
		2426: Delta = 34'sb0000000000000000010000000000000000;
		3885: Delta = 34'sb1111111111111111110000000000000000;
		4852: Delta = 34'sb0000000000000000100000000000000000;
		1459: Delta = 34'sb1111111111111111100000000000000000;
		3393: Delta = 34'sb0000000000000001000000000000000000;
		2918: Delta = 34'sb1111111111111111000000000000000000;
		475: Delta = 34'sb0000000000000010000000000000000000;
		5836: Delta = 34'sb1111111111111110000000000000000000;
		950: Delta = 34'sb0000000000000100000000000000000000;
		5361: Delta = 34'sb1111111111111100000000000000000000;
		1900: Delta = 34'sb0000000000001000000000000000000000;
		4411: Delta = 34'sb1111111111111000000000000000000000;
		3800: Delta = 34'sb0000000000010000000000000000000000;
		2511: Delta = 34'sb1111111111110000000000000000000000;
		1289: Delta = 34'sb0000000000100000000000000000000000;
		5022: Delta = 34'sb1111111111100000000000000000000000;
		2578: Delta = 34'sb0000000001000000000000000000000000;
		3733: Delta = 34'sb1111111111000000000000000000000000;
		5156: Delta = 34'sb0000000010000000000000000000000000;
		1155: Delta = 34'sb1111111110000000000000000000000000;
		4001: Delta = 34'sb0000000100000000000000000000000000;
		2310: Delta = 34'sb1111111100000000000000000000000000;
		1691: Delta = 34'sb0000001000000000000000000000000000;
		4620: Delta = 34'sb1111111000000000000000000000000000;
		3382: Delta = 34'sb0000010000000000000000000000000000;
		2929: Delta = 34'sb1111110000000000000000000000000000;
		453: Delta = 34'sb0000100000000000000000000000000000;
		5858: Delta = 34'sb1111100000000000000000000000000000;
		906: Delta = 34'sb0001000000000000000000000000000000;
		5405: Delta = 34'sb1111000000000000000000000000000000;
		1812: Delta = 34'sb0010000000000000000000000000000000;
		4499: Delta = 34'sb1110000000000000000000000000000000;
		3624: Delta = 34'sb0100000000000000000000000000000000;
		2687: Delta = 34'sb1100000000000000000000000000000000;
		default: Delta =34'sb0;
	endcase
end

assign N = (W - Delta) / A;

endmodule

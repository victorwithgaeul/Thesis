// Product (AN) Code SEC l-LUT
// SEC_lLUT16bits.v
// Received single error location l, output remainder r.
module SEC_lLUT16bits(l, r);
input	signed	[5:0]	l;
output	reg	[12:0]	r;
always@(*) begin
	case(l)
		1: r = 1;
		-1: r = 4546;
		2: r = 2;
		-2: r = 4545;
		3: r = 4;
		-3: r = 4543;
		4: r = 8;
		-4: r = 4539;
		5: r = 16;
		-5: r = 4531;
		6: r = 32;
		-6: r = 4515;
		7: r = 64;
		-7: r = 4483;
		8: r = 128;
		-8: r = 4419;
		9: r = 256;
		-9: r = 4291;
		10: r = 512;
		-10: r = 4035;
		11: r = 1024;
		-11: r = 3523;
		12: r = 2048;
		-12: r = 2499;
		13: r = 4096;
		-13: r = 451;
		14: r = 3645;
		-14: r = 902;
		15: r = 2743;
		-15: r = 1804;
		16: r = 939;
		-16: r = 3608;
		17: r = 1878;
		-17: r = 2669;
		18: r = 3756;
		-18: r = 791;
		19: r = 2965;
		-19: r = 1582;
		20: r = 1383;
		-20: r = 3164;
		21: r = 2766;
		-21: r = 1781;
		22: r = 985;
		-22: r = 3562;
		23: r = 1970;
		-23: r = 2577;
		24: r = 3940;
		-24: r = 607;
		25: r = 3333;
		-25: r = 1214;
		26: r = 2119;
		-26: r = 2428;
		27: r = 4238;
		-27: r = 309;
		28: r = 3929;
		-28: r = 618;
		29: r = 3311;
		-29: r = 1236;
		default: r = 0;
	endcase
end

endmodule

// Product (AN) Code DEC_LUT_Decoder
// DEC_LUT_Decoder12bits.v
// Received codeword W = AN + E, E is double AWE (E = e1 + e2), +2^i or -2^i.
module DEC_LUT_Decoder12bits(W, N);
input 	[23:0]	W;
output	[11:0]	N;
parameter A = 3349;

wire 	[11:0]	Q;
wire 	[11:0]	R;
assign Q = W / A;
assign R = W - (A * Q);

reg	signed	[24:0]	Delta;
always@(*) begin
	case(R)
		1: Delta = 25'sb0000000000000000000000001;
		3348: Delta = 25'sb1111111111111111111111111;
		2: Delta = 25'sb0000000000000000000000010;
		3347: Delta = 25'sb1111111111111111111111110;
		4: Delta = 25'sb0000000000000000000000100;
		3345: Delta = 25'sb1111111111111111111111100;
		8: Delta = 25'sb0000000000000000000001000;
		3341: Delta = 25'sb1111111111111111111111000;
		16: Delta = 25'sb0000000000000000000010000;
		3333: Delta = 25'sb1111111111111111111110000;
		32: Delta = 25'sb0000000000000000000100000;
		3317: Delta = 25'sb1111111111111111111100000;
		64: Delta = 25'sb0000000000000000001000000;
		3285: Delta = 25'sb1111111111111111111000000;
		128: Delta = 25'sb0000000000000000010000000;
		3221: Delta = 25'sb1111111111111111110000000;
		256: Delta = 25'sb0000000000000000100000000;
		3093: Delta = 25'sb1111111111111111100000000;
		512: Delta = 25'sb0000000000000001000000000;
		2837: Delta = 25'sb1111111111111111000000000;
		1024: Delta = 25'sb0000000000000010000000000;
		2325: Delta = 25'sb1111111111111110000000000;
		2048: Delta = 25'sb0000000000000100000000000;
		1301: Delta = 25'sb1111111111111100000000000;
		747: Delta = 25'sb0000000000001000000000000;
		2602: Delta = 25'sb1111111111111000000000000;
		1494: Delta = 25'sb0000000000010000000000000;
		1855: Delta = 25'sb1111111111110000000000000;
		2988: Delta = 25'sb0000000000100000000000000;
		361: Delta = 25'sb1111111111100000000000000;
		2627: Delta = 25'sb0000000001000000000000000;
		722: Delta = 25'sb1111111111000000000000000;
		1905: Delta = 25'sb0000000010000000000000000;
		1444: Delta = 25'sb1111111110000000000000000;
		461: Delta = 25'sb0000000100000000000000000;
		2888: Delta = 25'sb1111111100000000000000000;
		922: Delta = 25'sb0000001000000000000000000;
		2427: Delta = 25'sb1111111000000000000000000;
		1844: Delta = 25'sb0000010000000000000000000;
		1505: Delta = 25'sb1111110000000000000000000;
		339: Delta = 25'sb0000100000000000000000000;
		3010: Delta = 25'sb1111100000000000000000000;
		678: Delta = 25'sb0001000000000000000000000;
		2671: Delta = 25'sb1111000000000000000000000;
		1356: Delta = 25'sb0010000000000000000000000;
		1993: Delta = 25'sb1110000000000000000000000;
		2712: Delta = 25'sb0100000000000000000000000;
		637: Delta = 25'sb1100000000000000000000000;
		3: Delta = 25'sb0000000000000000000000011;
		3346: Delta = 25'sb1111111111111111111111101;
		5: Delta = 25'sb0000000000000000000000101;
		3344: Delta = 25'sb1111111111111111111111011;
		9: Delta = 25'sb0000000000000000000001001;
		3342: Delta = 25'sb1111111111111111111111001;
		7: Delta = 25'sb0000000000000000000000111;
		3340: Delta = 25'sb1111111111111111111110111;
		17: Delta = 25'sb0000000000000000000010001;
		3334: Delta = 25'sb1111111111111111111110001;
		15: Delta = 25'sb0000000000000000000001111;
		3332: Delta = 25'sb1111111111111111111101111;
		33: Delta = 25'sb0000000000000000000100001;
		3318: Delta = 25'sb1111111111111111111100001;
		31: Delta = 25'sb0000000000000000000011111;
		3316: Delta = 25'sb1111111111111111111011111;
		65: Delta = 25'sb0000000000000000001000001;
		3286: Delta = 25'sb1111111111111111111000001;
		63: Delta = 25'sb0000000000000000000111111;
		3284: Delta = 25'sb1111111111111111110111111;
		129: Delta = 25'sb0000000000000000010000001;
		3222: Delta = 25'sb1111111111111111110000001;
		127: Delta = 25'sb0000000000000000001111111;
		3220: Delta = 25'sb1111111111111111101111111;
		257: Delta = 25'sb0000000000000000100000001;
		3094: Delta = 25'sb1111111111111111100000001;
		255: Delta = 25'sb0000000000000000011111111;
		3092: Delta = 25'sb1111111111111111011111111;
		513: Delta = 25'sb0000000000000001000000001;
		2838: Delta = 25'sb1111111111111111000000001;
		511: Delta = 25'sb0000000000000000111111111;
		2836: Delta = 25'sb1111111111111110111111111;
		1025: Delta = 25'sb0000000000000010000000001;
		2326: Delta = 25'sb1111111111111110000000001;
		1023: Delta = 25'sb0000000000000001111111111;
		2324: Delta = 25'sb1111111111111101111111111;
		2049: Delta = 25'sb0000000000000100000000001;
		1302: Delta = 25'sb1111111111111100000000001;
		2047: Delta = 25'sb0000000000000011111111111;
		1300: Delta = 25'sb1111111111111011111111111;
		748: Delta = 25'sb0000000000001000000000001;
		2603: Delta = 25'sb1111111111111000000000001;
		746: Delta = 25'sb0000000000000111111111111;
		2601: Delta = 25'sb1111111111110111111111111;
		1495: Delta = 25'sb0000000000010000000000001;
		1856: Delta = 25'sb1111111111110000000000001;
		1493: Delta = 25'sb0000000000001111111111111;
		1854: Delta = 25'sb1111111111101111111111111;
		2989: Delta = 25'sb0000000000100000000000001;
		362: Delta = 25'sb1111111111100000000000001;
		2987: Delta = 25'sb0000000000011111111111111;
		360: Delta = 25'sb1111111111011111111111111;
		2628: Delta = 25'sb0000000001000000000000001;
		723: Delta = 25'sb1111111111000000000000001;
		2626: Delta = 25'sb0000000000111111111111111;
		721: Delta = 25'sb1111111110111111111111111;
		1906: Delta = 25'sb0000000010000000000000001;
		1445: Delta = 25'sb1111111110000000000000001;
		1904: Delta = 25'sb0000000001111111111111111;
		1443: Delta = 25'sb1111111101111111111111111;
		462: Delta = 25'sb0000000100000000000000001;
		2889: Delta = 25'sb1111111100000000000000001;
		460: Delta = 25'sb0000000011111111111111111;
		2887: Delta = 25'sb1111111011111111111111111;
		923: Delta = 25'sb0000001000000000000000001;
		2428: Delta = 25'sb1111111000000000000000001;
		921: Delta = 25'sb0000000111111111111111111;
		2426: Delta = 25'sb1111110111111111111111111;
		1845: Delta = 25'sb0000010000000000000000001;
		1506: Delta = 25'sb1111110000000000000000001;
		1843: Delta = 25'sb0000001111111111111111111;
		1504: Delta = 25'sb1111101111111111111111111;
		340: Delta = 25'sb0000100000000000000000001;
		3011: Delta = 25'sb1111100000000000000000001;
		338: Delta = 25'sb0000011111111111111111111;
		3009: Delta = 25'sb1111011111111111111111111;
		679: Delta = 25'sb0001000000000000000000001;
		2672: Delta = 25'sb1111000000000000000000001;
		677: Delta = 25'sb0000111111111111111111111;
		2670: Delta = 25'sb1110111111111111111111111;
		1357: Delta = 25'sb0010000000000000000000001;
		1994: Delta = 25'sb1110000000000000000000001;
		1355: Delta = 25'sb0001111111111111111111111;
		1992: Delta = 25'sb1101111111111111111111111;
		2713: Delta = 25'sb0100000000000000000000001;
		638: Delta = 25'sb1100000000000000000000001;
		2711: Delta = 25'sb0011111111111111111111111;
		636: Delta = 25'sb1011111111111111111111111;
		6: Delta = 25'sb0000000000000000000000110;
		3343: Delta = 25'sb1111111111111111111111010;
		10: Delta = 25'sb0000000000000000000001010;
		3339: Delta = 25'sb1111111111111111111110110;
		18: Delta = 25'sb0000000000000000000010010;
		3335: Delta = 25'sb1111111111111111111110010;
		14: Delta = 25'sb0000000000000000000001110;
		3331: Delta = 25'sb1111111111111111111101110;
		34: Delta = 25'sb0000000000000000000100010;
		3319: Delta = 25'sb1111111111111111111100010;
		30: Delta = 25'sb0000000000000000000011110;
		3315: Delta = 25'sb1111111111111111111011110;
		66: Delta = 25'sb0000000000000000001000010;
		3287: Delta = 25'sb1111111111111111111000010;
		62: Delta = 25'sb0000000000000000000111110;
		3283: Delta = 25'sb1111111111111111110111110;
		130: Delta = 25'sb0000000000000000010000010;
		3223: Delta = 25'sb1111111111111111110000010;
		126: Delta = 25'sb0000000000000000001111110;
		3219: Delta = 25'sb1111111111111111101111110;
		258: Delta = 25'sb0000000000000000100000010;
		3095: Delta = 25'sb1111111111111111100000010;
		254: Delta = 25'sb0000000000000000011111110;
		3091: Delta = 25'sb1111111111111111011111110;
		514: Delta = 25'sb0000000000000001000000010;
		2839: Delta = 25'sb1111111111111111000000010;
		510: Delta = 25'sb0000000000000000111111110;
		2835: Delta = 25'sb1111111111111110111111110;
		1026: Delta = 25'sb0000000000000010000000010;
		2327: Delta = 25'sb1111111111111110000000010;
		1022: Delta = 25'sb0000000000000001111111110;
		2323: Delta = 25'sb1111111111111101111111110;
		2050: Delta = 25'sb0000000000000100000000010;
		1303: Delta = 25'sb1111111111111100000000010;
		2046: Delta = 25'sb0000000000000011111111110;
		1299: Delta = 25'sb1111111111111011111111110;
		749: Delta = 25'sb0000000000001000000000010;
		2604: Delta = 25'sb1111111111111000000000010;
		745: Delta = 25'sb0000000000000111111111110;
		2600: Delta = 25'sb1111111111110111111111110;
		1496: Delta = 25'sb0000000000010000000000010;
		1857: Delta = 25'sb1111111111110000000000010;
		1492: Delta = 25'sb0000000000001111111111110;
		1853: Delta = 25'sb1111111111101111111111110;
		2990: Delta = 25'sb0000000000100000000000010;
		363: Delta = 25'sb1111111111100000000000010;
		2986: Delta = 25'sb0000000000011111111111110;
		359: Delta = 25'sb1111111111011111111111110;
		2629: Delta = 25'sb0000000001000000000000010;
		724: Delta = 25'sb1111111111000000000000010;
		2625: Delta = 25'sb0000000000111111111111110;
		720: Delta = 25'sb1111111110111111111111110;
		1907: Delta = 25'sb0000000010000000000000010;
		1446: Delta = 25'sb1111111110000000000000010;
		1903: Delta = 25'sb0000000001111111111111110;
		1442: Delta = 25'sb1111111101111111111111110;
		463: Delta = 25'sb0000000100000000000000010;
		2890: Delta = 25'sb1111111100000000000000010;
		459: Delta = 25'sb0000000011111111111111110;
		2886: Delta = 25'sb1111111011111111111111110;
		924: Delta = 25'sb0000001000000000000000010;
		2429: Delta = 25'sb1111111000000000000000010;
		920: Delta = 25'sb0000000111111111111111110;
		2425: Delta = 25'sb1111110111111111111111110;
		1846: Delta = 25'sb0000010000000000000000010;
		1507: Delta = 25'sb1111110000000000000000010;
		1842: Delta = 25'sb0000001111111111111111110;
		1503: Delta = 25'sb1111101111111111111111110;
		341: Delta = 25'sb0000100000000000000000010;
		3012: Delta = 25'sb1111100000000000000000010;
		337: Delta = 25'sb0000011111111111111111110;
		3008: Delta = 25'sb1111011111111111111111110;
		680: Delta = 25'sb0001000000000000000000010;
		2673: Delta = 25'sb1111000000000000000000010;
		676: Delta = 25'sb0000111111111111111111110;
		2669: Delta = 25'sb1110111111111111111111110;
		1358: Delta = 25'sb0010000000000000000000010;
		1995: Delta = 25'sb1110000000000000000000010;
		1354: Delta = 25'sb0001111111111111111111110;
		1991: Delta = 25'sb1101111111111111111111110;
		2714: Delta = 25'sb0100000000000000000000010;
		639: Delta = 25'sb1100000000000000000000010;
		2710: Delta = 25'sb0011111111111111111111110;
		635: Delta = 25'sb1011111111111111111111110;
		12: Delta = 25'sb0000000000000000000001100;
		3337: Delta = 25'sb1111111111111111111110100;
		20: Delta = 25'sb0000000000000000000010100;
		3329: Delta = 25'sb1111111111111111111101100;
		36: Delta = 25'sb0000000000000000000100100;
		3321: Delta = 25'sb1111111111111111111100100;
		28: Delta = 25'sb0000000000000000000011100;
		3313: Delta = 25'sb1111111111111111111011100;
		68: Delta = 25'sb0000000000000000001000100;
		3289: Delta = 25'sb1111111111111111111000100;
		60: Delta = 25'sb0000000000000000000111100;
		3281: Delta = 25'sb1111111111111111110111100;
		132: Delta = 25'sb0000000000000000010000100;
		3225: Delta = 25'sb1111111111111111110000100;
		124: Delta = 25'sb0000000000000000001111100;
		3217: Delta = 25'sb1111111111111111101111100;
		260: Delta = 25'sb0000000000000000100000100;
		3097: Delta = 25'sb1111111111111111100000100;
		252: Delta = 25'sb0000000000000000011111100;
		3089: Delta = 25'sb1111111111111111011111100;
		516: Delta = 25'sb0000000000000001000000100;
		2841: Delta = 25'sb1111111111111111000000100;
		508: Delta = 25'sb0000000000000000111111100;
		2833: Delta = 25'sb1111111111111110111111100;
		1028: Delta = 25'sb0000000000000010000000100;
		2329: Delta = 25'sb1111111111111110000000100;
		1020: Delta = 25'sb0000000000000001111111100;
		2321: Delta = 25'sb1111111111111101111111100;
		2052: Delta = 25'sb0000000000000100000000100;
		1305: Delta = 25'sb1111111111111100000000100;
		2044: Delta = 25'sb0000000000000011111111100;
		1297: Delta = 25'sb1111111111111011111111100;
		751: Delta = 25'sb0000000000001000000000100;
		2606: Delta = 25'sb1111111111111000000000100;
		743: Delta = 25'sb0000000000000111111111100;
		2598: Delta = 25'sb1111111111110111111111100;
		1498: Delta = 25'sb0000000000010000000000100;
		1859: Delta = 25'sb1111111111110000000000100;
		1490: Delta = 25'sb0000000000001111111111100;
		1851: Delta = 25'sb1111111111101111111111100;
		2992: Delta = 25'sb0000000000100000000000100;
		365: Delta = 25'sb1111111111100000000000100;
		2984: Delta = 25'sb0000000000011111111111100;
		357: Delta = 25'sb1111111111011111111111100;
		2631: Delta = 25'sb0000000001000000000000100;
		726: Delta = 25'sb1111111111000000000000100;
		2623: Delta = 25'sb0000000000111111111111100;
		718: Delta = 25'sb1111111110111111111111100;
		1909: Delta = 25'sb0000000010000000000000100;
		1448: Delta = 25'sb1111111110000000000000100;
		1901: Delta = 25'sb0000000001111111111111100;
		1440: Delta = 25'sb1111111101111111111111100;
		465: Delta = 25'sb0000000100000000000000100;
		2892: Delta = 25'sb1111111100000000000000100;
		457: Delta = 25'sb0000000011111111111111100;
		2884: Delta = 25'sb1111111011111111111111100;
		926: Delta = 25'sb0000001000000000000000100;
		2431: Delta = 25'sb1111111000000000000000100;
		918: Delta = 25'sb0000000111111111111111100;
		2423: Delta = 25'sb1111110111111111111111100;
		1848: Delta = 25'sb0000010000000000000000100;
		1509: Delta = 25'sb1111110000000000000000100;
		1840: Delta = 25'sb0000001111111111111111100;
		1501: Delta = 25'sb1111101111111111111111100;
		343: Delta = 25'sb0000100000000000000000100;
		3014: Delta = 25'sb1111100000000000000000100;
		335: Delta = 25'sb0000011111111111111111100;
		3006: Delta = 25'sb1111011111111111111111100;
		682: Delta = 25'sb0001000000000000000000100;
		2675: Delta = 25'sb1111000000000000000000100;
		674: Delta = 25'sb0000111111111111111111100;
		2667: Delta = 25'sb1110111111111111111111100;
		1360: Delta = 25'sb0010000000000000000000100;
		1997: Delta = 25'sb1110000000000000000000100;
		1352: Delta = 25'sb0001111111111111111111100;
		1989: Delta = 25'sb1101111111111111111111100;
		2716: Delta = 25'sb0100000000000000000000100;
		641: Delta = 25'sb1100000000000000000000100;
		2708: Delta = 25'sb0011111111111111111111100;
		633: Delta = 25'sb1011111111111111111111100;
		24: Delta = 25'sb0000000000000000000011000;
		3325: Delta = 25'sb1111111111111111111101000;
		40: Delta = 25'sb0000000000000000000101000;
		3309: Delta = 25'sb1111111111111111111011000;
		72: Delta = 25'sb0000000000000000001001000;
		3293: Delta = 25'sb1111111111111111111001000;
		56: Delta = 25'sb0000000000000000000111000;
		3277: Delta = 25'sb1111111111111111110111000;
		136: Delta = 25'sb0000000000000000010001000;
		3229: Delta = 25'sb1111111111111111110001000;
		120: Delta = 25'sb0000000000000000001111000;
		3213: Delta = 25'sb1111111111111111101111000;
		264: Delta = 25'sb0000000000000000100001000;
		3101: Delta = 25'sb1111111111111111100001000;
		248: Delta = 25'sb0000000000000000011111000;
		3085: Delta = 25'sb1111111111111111011111000;
		520: Delta = 25'sb0000000000000001000001000;
		2845: Delta = 25'sb1111111111111111000001000;
		504: Delta = 25'sb0000000000000000111111000;
		2829: Delta = 25'sb1111111111111110111111000;
		1032: Delta = 25'sb0000000000000010000001000;
		2333: Delta = 25'sb1111111111111110000001000;
		1016: Delta = 25'sb0000000000000001111111000;
		2317: Delta = 25'sb1111111111111101111111000;
		2056: Delta = 25'sb0000000000000100000001000;
		1309: Delta = 25'sb1111111111111100000001000;
		2040: Delta = 25'sb0000000000000011111111000;
		1293: Delta = 25'sb1111111111111011111111000;
		755: Delta = 25'sb0000000000001000000001000;
		2610: Delta = 25'sb1111111111111000000001000;
		739: Delta = 25'sb0000000000000111111111000;
		2594: Delta = 25'sb1111111111110111111111000;
		1502: Delta = 25'sb0000000000010000000001000;
		1863: Delta = 25'sb1111111111110000000001000;
		1486: Delta = 25'sb0000000000001111111111000;
		1847: Delta = 25'sb1111111111101111111111000;
		2996: Delta = 25'sb0000000000100000000001000;
		369: Delta = 25'sb1111111111100000000001000;
		2980: Delta = 25'sb0000000000011111111111000;
		353: Delta = 25'sb1111111111011111111111000;
		2635: Delta = 25'sb0000000001000000000001000;
		730: Delta = 25'sb1111111111000000000001000;
		2619: Delta = 25'sb0000000000111111111111000;
		714: Delta = 25'sb1111111110111111111111000;
		1913: Delta = 25'sb0000000010000000000001000;
		1452: Delta = 25'sb1111111110000000000001000;
		1897: Delta = 25'sb0000000001111111111111000;
		1436: Delta = 25'sb1111111101111111111111000;
		469: Delta = 25'sb0000000100000000000001000;
		2896: Delta = 25'sb1111111100000000000001000;
		453: Delta = 25'sb0000000011111111111111000;
		2880: Delta = 25'sb1111111011111111111111000;
		930: Delta = 25'sb0000001000000000000001000;
		2435: Delta = 25'sb1111111000000000000001000;
		914: Delta = 25'sb0000000111111111111111000;
		2419: Delta = 25'sb1111110111111111111111000;
		1852: Delta = 25'sb0000010000000000000001000;
		1513: Delta = 25'sb1111110000000000000001000;
		1836: Delta = 25'sb0000001111111111111111000;
		1497: Delta = 25'sb1111101111111111111111000;
		347: Delta = 25'sb0000100000000000000001000;
		3018: Delta = 25'sb1111100000000000000001000;
		331: Delta = 25'sb0000011111111111111111000;
		3002: Delta = 25'sb1111011111111111111111000;
		686: Delta = 25'sb0001000000000000000001000;
		2679: Delta = 25'sb1111000000000000000001000;
		670: Delta = 25'sb0000111111111111111111000;
		2663: Delta = 25'sb1110111111111111111111000;
		1364: Delta = 25'sb0010000000000000000001000;
		2001: Delta = 25'sb1110000000000000000001000;
		1348: Delta = 25'sb0001111111111111111111000;
		1985: Delta = 25'sb1101111111111111111111000;
		2720: Delta = 25'sb0100000000000000000001000;
		645: Delta = 25'sb1100000000000000000001000;
		2704: Delta = 25'sb0011111111111111111111000;
		629: Delta = 25'sb1011111111111111111111000;
		48: Delta = 25'sb0000000000000000000110000;
		3301: Delta = 25'sb1111111111111111111010000;
		80: Delta = 25'sb0000000000000000001010000;
		3269: Delta = 25'sb1111111111111111110110000;
		144: Delta = 25'sb0000000000000000010010000;
		3237: Delta = 25'sb1111111111111111110010000;
		112: Delta = 25'sb0000000000000000001110000;
		3205: Delta = 25'sb1111111111111111101110000;
		272: Delta = 25'sb0000000000000000100010000;
		3109: Delta = 25'sb1111111111111111100010000;
		240: Delta = 25'sb0000000000000000011110000;
		3077: Delta = 25'sb1111111111111111011110000;
		528: Delta = 25'sb0000000000000001000010000;
		2853: Delta = 25'sb1111111111111111000010000;
		496: Delta = 25'sb0000000000000000111110000;
		2821: Delta = 25'sb1111111111111110111110000;
		1040: Delta = 25'sb0000000000000010000010000;
		2341: Delta = 25'sb1111111111111110000010000;
		1008: Delta = 25'sb0000000000000001111110000;
		2309: Delta = 25'sb1111111111111101111110000;
		2064: Delta = 25'sb0000000000000100000010000;
		1317: Delta = 25'sb1111111111111100000010000;
		2032: Delta = 25'sb0000000000000011111110000;
		1285: Delta = 25'sb1111111111111011111110000;
		763: Delta = 25'sb0000000000001000000010000;
		2618: Delta = 25'sb1111111111111000000010000;
		731: Delta = 25'sb0000000000000111111110000;
		2586: Delta = 25'sb1111111111110111111110000;
		1510: Delta = 25'sb0000000000010000000010000;
		1871: Delta = 25'sb1111111111110000000010000;
		1478: Delta = 25'sb0000000000001111111110000;
		1839: Delta = 25'sb1111111111101111111110000;
		3004: Delta = 25'sb0000000000100000000010000;
		377: Delta = 25'sb1111111111100000000010000;
		2972: Delta = 25'sb0000000000011111111110000;
		345: Delta = 25'sb1111111111011111111110000;
		2643: Delta = 25'sb0000000001000000000010000;
		738: Delta = 25'sb1111111111000000000010000;
		2611: Delta = 25'sb0000000000111111111110000;
		706: Delta = 25'sb1111111110111111111110000;
		1921: Delta = 25'sb0000000010000000000010000;
		1460: Delta = 25'sb1111111110000000000010000;
		1889: Delta = 25'sb0000000001111111111110000;
		1428: Delta = 25'sb1111111101111111111110000;
		477: Delta = 25'sb0000000100000000000010000;
		2904: Delta = 25'sb1111111100000000000010000;
		445: Delta = 25'sb0000000011111111111110000;
		2872: Delta = 25'sb1111111011111111111110000;
		938: Delta = 25'sb0000001000000000000010000;
		2443: Delta = 25'sb1111111000000000000010000;
		906: Delta = 25'sb0000000111111111111110000;
		2411: Delta = 25'sb1111110111111111111110000;
		1860: Delta = 25'sb0000010000000000000010000;
		1521: Delta = 25'sb1111110000000000000010000;
		1828: Delta = 25'sb0000001111111111111110000;
		1489: Delta = 25'sb1111101111111111111110000;
		355: Delta = 25'sb0000100000000000000010000;
		3026: Delta = 25'sb1111100000000000000010000;
		323: Delta = 25'sb0000011111111111111110000;
		2994: Delta = 25'sb1111011111111111111110000;
		694: Delta = 25'sb0001000000000000000010000;
		2687: Delta = 25'sb1111000000000000000010000;
		662: Delta = 25'sb0000111111111111111110000;
		2655: Delta = 25'sb1110111111111111111110000;
		1372: Delta = 25'sb0010000000000000000010000;
		2009: Delta = 25'sb1110000000000000000010000;
		1340: Delta = 25'sb0001111111111111111110000;
		1977: Delta = 25'sb1101111111111111111110000;
		2728: Delta = 25'sb0100000000000000000010000;
		653: Delta = 25'sb1100000000000000000010000;
		2696: Delta = 25'sb0011111111111111111110000;
		621: Delta = 25'sb1011111111111111111110000;
		96: Delta = 25'sb0000000000000000001100000;
		3253: Delta = 25'sb1111111111111111110100000;
		160: Delta = 25'sb0000000000000000010100000;
		3189: Delta = 25'sb1111111111111111101100000;
		288: Delta = 25'sb0000000000000000100100000;
		3125: Delta = 25'sb1111111111111111100100000;
		224: Delta = 25'sb0000000000000000011100000;
		3061: Delta = 25'sb1111111111111111011100000;
		544: Delta = 25'sb0000000000000001000100000;
		2869: Delta = 25'sb1111111111111111000100000;
		480: Delta = 25'sb0000000000000000111100000;
		2805: Delta = 25'sb1111111111111110111100000;
		1056: Delta = 25'sb0000000000000010000100000;
		2357: Delta = 25'sb1111111111111110000100000;
		992: Delta = 25'sb0000000000000001111100000;
		2293: Delta = 25'sb1111111111111101111100000;
		2080: Delta = 25'sb0000000000000100000100000;
		1333: Delta = 25'sb1111111111111100000100000;
		2016: Delta = 25'sb0000000000000011111100000;
		1269: Delta = 25'sb1111111111111011111100000;
		779: Delta = 25'sb0000000000001000000100000;
		2634: Delta = 25'sb1111111111111000000100000;
		715: Delta = 25'sb0000000000000111111100000;
		2570: Delta = 25'sb1111111111110111111100000;
		1526: Delta = 25'sb0000000000010000000100000;
		1887: Delta = 25'sb1111111111110000000100000;
		1462: Delta = 25'sb0000000000001111111100000;
		1823: Delta = 25'sb1111111111101111111100000;
		3020: Delta = 25'sb0000000000100000000100000;
		393: Delta = 25'sb1111111111100000000100000;
		2956: Delta = 25'sb0000000000011111111100000;
		329: Delta = 25'sb1111111111011111111100000;
		2659: Delta = 25'sb0000000001000000000100000;
		754: Delta = 25'sb1111111111000000000100000;
		2595: Delta = 25'sb0000000000111111111100000;
		690: Delta = 25'sb1111111110111111111100000;
		1937: Delta = 25'sb0000000010000000000100000;
		1476: Delta = 25'sb1111111110000000000100000;
		1873: Delta = 25'sb0000000001111111111100000;
		1412: Delta = 25'sb1111111101111111111100000;
		493: Delta = 25'sb0000000100000000000100000;
		2920: Delta = 25'sb1111111100000000000100000;
		429: Delta = 25'sb0000000011111111111100000;
		2856: Delta = 25'sb1111111011111111111100000;
		954: Delta = 25'sb0000001000000000000100000;
		2459: Delta = 25'sb1111111000000000000100000;
		890: Delta = 25'sb0000000111111111111100000;
		2395: Delta = 25'sb1111110111111111111100000;
		1876: Delta = 25'sb0000010000000000000100000;
		1537: Delta = 25'sb1111110000000000000100000;
		1812: Delta = 25'sb0000001111111111111100000;
		1473: Delta = 25'sb1111101111111111111100000;
		371: Delta = 25'sb0000100000000000000100000;
		3042: Delta = 25'sb1111100000000000000100000;
		307: Delta = 25'sb0000011111111111111100000;
		2978: Delta = 25'sb1111011111111111111100000;
		710: Delta = 25'sb0001000000000000000100000;
		2703: Delta = 25'sb1111000000000000000100000;
		646: Delta = 25'sb0000111111111111111100000;
		2639: Delta = 25'sb1110111111111111111100000;
		1388: Delta = 25'sb0010000000000000000100000;
		2025: Delta = 25'sb1110000000000000000100000;
		1324: Delta = 25'sb0001111111111111111100000;
		1961: Delta = 25'sb1101111111111111111100000;
		2744: Delta = 25'sb0100000000000000000100000;
		669: Delta = 25'sb1100000000000000000100000;
		2680: Delta = 25'sb0011111111111111111100000;
		605: Delta = 25'sb1011111111111111111100000;
		192: Delta = 25'sb0000000000000000011000000;
		3157: Delta = 25'sb1111111111111111101000000;
		320: Delta = 25'sb0000000000000000101000000;
		3029: Delta = 25'sb1111111111111111011000000;
		576: Delta = 25'sb0000000000000001001000000;
		2901: Delta = 25'sb1111111111111111001000000;
		448: Delta = 25'sb0000000000000000111000000;
		2773: Delta = 25'sb1111111111111110111000000;
		1088: Delta = 25'sb0000000000000010001000000;
		2389: Delta = 25'sb1111111111111110001000000;
		960: Delta = 25'sb0000000000000001111000000;
		2261: Delta = 25'sb1111111111111101111000000;
		2112: Delta = 25'sb0000000000000100001000000;
		1365: Delta = 25'sb1111111111111100001000000;
		1984: Delta = 25'sb0000000000000011111000000;
		1237: Delta = 25'sb1111111111111011111000000;
		811: Delta = 25'sb0000000000001000001000000;
		2666: Delta = 25'sb1111111111111000001000000;
		683: Delta = 25'sb0000000000000111111000000;
		2538: Delta = 25'sb1111111111110111111000000;
		1558: Delta = 25'sb0000000000010000001000000;
		1919: Delta = 25'sb1111111111110000001000000;
		1430: Delta = 25'sb0000000000001111111000000;
		1791: Delta = 25'sb1111111111101111111000000;
		3052: Delta = 25'sb0000000000100000001000000;
		425: Delta = 25'sb1111111111100000001000000;
		2924: Delta = 25'sb0000000000011111111000000;
		297: Delta = 25'sb1111111111011111111000000;
		2691: Delta = 25'sb0000000001000000001000000;
		786: Delta = 25'sb1111111111000000001000000;
		2563: Delta = 25'sb0000000000111111111000000;
		658: Delta = 25'sb1111111110111111111000000;
		1969: Delta = 25'sb0000000010000000001000000;
		1508: Delta = 25'sb1111111110000000001000000;
		1841: Delta = 25'sb0000000001111111111000000;
		1380: Delta = 25'sb1111111101111111111000000;
		525: Delta = 25'sb0000000100000000001000000;
		2952: Delta = 25'sb1111111100000000001000000;
		397: Delta = 25'sb0000000011111111111000000;
		2824: Delta = 25'sb1111111011111111111000000;
		986: Delta = 25'sb0000001000000000001000000;
		2491: Delta = 25'sb1111111000000000001000000;
		858: Delta = 25'sb0000000111111111111000000;
		2363: Delta = 25'sb1111110111111111111000000;
		1908: Delta = 25'sb0000010000000000001000000;
		1569: Delta = 25'sb1111110000000000001000000;
		1780: Delta = 25'sb0000001111111111111000000;
		1441: Delta = 25'sb1111101111111111111000000;
		403: Delta = 25'sb0000100000000000001000000;
		3074: Delta = 25'sb1111100000000000001000000;
		275: Delta = 25'sb0000011111111111111000000;
		2946: Delta = 25'sb1111011111111111111000000;
		742: Delta = 25'sb0001000000000000001000000;
		2735: Delta = 25'sb1111000000000000001000000;
		614: Delta = 25'sb0000111111111111111000000;
		2607: Delta = 25'sb1110111111111111111000000;
		1420: Delta = 25'sb0010000000000000001000000;
		2057: Delta = 25'sb1110000000000000001000000;
		1292: Delta = 25'sb0001111111111111111000000;
		1929: Delta = 25'sb1101111111111111111000000;
		2776: Delta = 25'sb0100000000000000001000000;
		701: Delta = 25'sb1100000000000000001000000;
		2648: Delta = 25'sb0011111111111111111000000;
		573: Delta = 25'sb1011111111111111111000000;
		384: Delta = 25'sb0000000000000000110000000;
		2965: Delta = 25'sb1111111111111111010000000;
		640: Delta = 25'sb0000000000000001010000000;
		2709: Delta = 25'sb1111111111111110110000000;
		1152: Delta = 25'sb0000000000000010010000000;
		2453: Delta = 25'sb1111111111111110010000000;
		896: Delta = 25'sb0000000000000001110000000;
		2197: Delta = 25'sb1111111111111101110000000;
		2176: Delta = 25'sb0000000000000100010000000;
		1429: Delta = 25'sb1111111111111100010000000;
		1920: Delta = 25'sb0000000000000011110000000;
		1173: Delta = 25'sb1111111111111011110000000;
		875: Delta = 25'sb0000000000001000010000000;
		2730: Delta = 25'sb1111111111111000010000000;
		619: Delta = 25'sb0000000000000111110000000;
		2474: Delta = 25'sb1111111111110111110000000;
		1622: Delta = 25'sb0000000000010000010000000;
		1983: Delta = 25'sb1111111111110000010000000;
		1366: Delta = 25'sb0000000000001111110000000;
		1727: Delta = 25'sb1111111111101111110000000;
		3116: Delta = 25'sb0000000000100000010000000;
		489: Delta = 25'sb1111111111100000010000000;
		2860: Delta = 25'sb0000000000011111110000000;
		233: Delta = 25'sb1111111111011111110000000;
		2755: Delta = 25'sb0000000001000000010000000;
		850: Delta = 25'sb1111111111000000010000000;
		2499: Delta = 25'sb0000000000111111110000000;
		594: Delta = 25'sb1111111110111111110000000;
		2033: Delta = 25'sb0000000010000000010000000;
		1572: Delta = 25'sb1111111110000000010000000;
		1777: Delta = 25'sb0000000001111111110000000;
		1316: Delta = 25'sb1111111101111111110000000;
		589: Delta = 25'sb0000000100000000010000000;
		3016: Delta = 25'sb1111111100000000010000000;
		333: Delta = 25'sb0000000011111111110000000;
		2760: Delta = 25'sb1111111011111111110000000;
		1050: Delta = 25'sb0000001000000000010000000;
		2555: Delta = 25'sb1111111000000000010000000;
		794: Delta = 25'sb0000000111111111110000000;
		2299: Delta = 25'sb1111110111111111110000000;
		1972: Delta = 25'sb0000010000000000010000000;
		1633: Delta = 25'sb1111110000000000010000000;
		1716: Delta = 25'sb0000001111111111110000000;
		1377: Delta = 25'sb1111101111111111110000000;
		467: Delta = 25'sb0000100000000000010000000;
		3138: Delta = 25'sb1111100000000000010000000;
		211: Delta = 25'sb0000011111111111110000000;
		2882: Delta = 25'sb1111011111111111110000000;
		806: Delta = 25'sb0001000000000000010000000;
		2799: Delta = 25'sb1111000000000000010000000;
		550: Delta = 25'sb0000111111111111110000000;
		2543: Delta = 25'sb1110111111111111110000000;
		1484: Delta = 25'sb0010000000000000010000000;
		2121: Delta = 25'sb1110000000000000010000000;
		1228: Delta = 25'sb0001111111111111110000000;
		1865: Delta = 25'sb1101111111111111110000000;
		2840: Delta = 25'sb0100000000000000010000000;
		765: Delta = 25'sb1100000000000000010000000;
		2584: Delta = 25'sb0011111111111111110000000;
		509: Delta = 25'sb1011111111111111110000000;
		768: Delta = 25'sb0000000000000001100000000;
		2581: Delta = 25'sb1111111111111110100000000;
		1280: Delta = 25'sb0000000000000010100000000;
		2069: Delta = 25'sb1111111111111101100000000;
		2304: Delta = 25'sb0000000000000100100000000;
		1557: Delta = 25'sb1111111111111100100000000;
		1792: Delta = 25'sb0000000000000011100000000;
		1045: Delta = 25'sb1111111111111011100000000;
		1003: Delta = 25'sb0000000000001000100000000;
		2858: Delta = 25'sb1111111111111000100000000;
		491: Delta = 25'sb0000000000000111100000000;
		2346: Delta = 25'sb1111111111110111100000000;
		1750: Delta = 25'sb0000000000010000100000000;
		2111: Delta = 25'sb1111111111110000100000000;
		1238: Delta = 25'sb0000000000001111100000000;
		1599: Delta = 25'sb1111111111101111100000000;
		3244: Delta = 25'sb0000000000100000100000000;
		617: Delta = 25'sb1111111111100000100000000;
		2732: Delta = 25'sb0000000000011111100000000;
		105: Delta = 25'sb1111111111011111100000000;
		2883: Delta = 25'sb0000000001000000100000000;
		978: Delta = 25'sb1111111111000000100000000;
		2371: Delta = 25'sb0000000000111111100000000;
		466: Delta = 25'sb1111111110111111100000000;
		2161: Delta = 25'sb0000000010000000100000000;
		1700: Delta = 25'sb1111111110000000100000000;
		1649: Delta = 25'sb0000000001111111100000000;
		1188: Delta = 25'sb1111111101111111100000000;
		717: Delta = 25'sb0000000100000000100000000;
		3144: Delta = 25'sb1111111100000000100000000;
		205: Delta = 25'sb0000000011111111100000000;
		2632: Delta = 25'sb1111111011111111100000000;
		1178: Delta = 25'sb0000001000000000100000000;
		2683: Delta = 25'sb1111111000000000100000000;
		666: Delta = 25'sb0000000111111111100000000;
		2171: Delta = 25'sb1111110111111111100000000;
		2100: Delta = 25'sb0000010000000000100000000;
		1761: Delta = 25'sb1111110000000000100000000;
		1588: Delta = 25'sb0000001111111111100000000;
		1249: Delta = 25'sb1111101111111111100000000;
		595: Delta = 25'sb0000100000000000100000000;
		3266: Delta = 25'sb1111100000000000100000000;
		83: Delta = 25'sb0000011111111111100000000;
		2754: Delta = 25'sb1111011111111111100000000;
		934: Delta = 25'sb0001000000000000100000000;
		2927: Delta = 25'sb1111000000000000100000000;
		422: Delta = 25'sb0000111111111111100000000;
		2415: Delta = 25'sb1110111111111111100000000;
		1612: Delta = 25'sb0010000000000000100000000;
		2249: Delta = 25'sb1110000000000000100000000;
		1100: Delta = 25'sb0001111111111111100000000;
		1737: Delta = 25'sb1101111111111111100000000;
		2968: Delta = 25'sb0100000000000000100000000;
		893: Delta = 25'sb1100000000000000100000000;
		2456: Delta = 25'sb0011111111111111100000000;
		381: Delta = 25'sb1011111111111111100000000;
		1536: Delta = 25'sb0000000000000011000000000;
		1813: Delta = 25'sb1111111111111101000000000;
		2560: Delta = 25'sb0000000000000101000000000;
		789: Delta = 25'sb1111111111111011000000000;
		1259: Delta = 25'sb0000000000001001000000000;
		3114: Delta = 25'sb1111111111111001000000000;
		235: Delta = 25'sb0000000000000111000000000;
		2090: Delta = 25'sb1111111111110111000000000;
		2006: Delta = 25'sb0000000000010001000000000;
		2367: Delta = 25'sb1111111111110001000000000;
		982: Delta = 25'sb0000000000001111000000000;
		1343: Delta = 25'sb1111111111101111000000000;
		151: Delta = 25'sb0000000000100001000000000;
		873: Delta = 25'sb1111111111100001000000000;
		2476: Delta = 25'sb0000000000011111000000000;
		3198: Delta = 25'sb1111111111011111000000000;
		3139: Delta = 25'sb0000000001000001000000000;
		1234: Delta = 25'sb1111111111000001000000000;
		2115: Delta = 25'sb0000000000111111000000000;
		210: Delta = 25'sb1111111110111111000000000;
		2417: Delta = 25'sb0000000010000001000000000;
		1956: Delta = 25'sb1111111110000001000000000;
		1393: Delta = 25'sb0000000001111111000000000;
		932: Delta = 25'sb1111111101111111000000000;
		973: Delta = 25'sb0000000100000001000000000;
		51: Delta = 25'sb1111111100000001000000000;
		3298: Delta = 25'sb0000000011111111000000000;
		2376: Delta = 25'sb1111111011111111000000000;
		1434: Delta = 25'sb0000001000000001000000000;
		2939: Delta = 25'sb1111111000000001000000000;
		410: Delta = 25'sb0000000111111111000000000;
		1915: Delta = 25'sb1111110111111111000000000;
		2356: Delta = 25'sb0000010000000001000000000;
		2017: Delta = 25'sb1111110000000001000000000;
		1332: Delta = 25'sb0000001111111111000000000;
		993: Delta = 25'sb1111101111111111000000000;
		851: Delta = 25'sb0000100000000001000000000;
		173: Delta = 25'sb1111100000000001000000000;
		3176: Delta = 25'sb0000011111111111000000000;
		2498: Delta = 25'sb1111011111111111000000000;
		1190: Delta = 25'sb0001000000000001000000000;
		3183: Delta = 25'sb1111000000000001000000000;
		166: Delta = 25'sb0000111111111111000000000;
		2159: Delta = 25'sb1110111111111111000000000;
		1868: Delta = 25'sb0010000000000001000000000;
		2505: Delta = 25'sb1110000000000001000000000;
		844: Delta = 25'sb0001111111111111000000000;
		1481: Delta = 25'sb1101111111111111000000000;
		3224: Delta = 25'sb0100000000000001000000000;
		1149: Delta = 25'sb1100000000000001000000000;
		2200: Delta = 25'sb0011111111111111000000000;
		125: Delta = 25'sb1011111111111111000000000;
		3072: Delta = 25'sb0000000000000110000000000;
		277: Delta = 25'sb1111111111111010000000000;
		1771: Delta = 25'sb0000000000001010000000000;
		1578: Delta = 25'sb1111111111110110000000000;
		2518: Delta = 25'sb0000000000010010000000000;
		2879: Delta = 25'sb1111111111110010000000000;
		470: Delta = 25'sb0000000000001110000000000;
		831: Delta = 25'sb1111111111101110000000000;
		663: Delta = 25'sb0000000000100010000000000;
		1385: Delta = 25'sb1111111111100010000000000;
		1964: Delta = 25'sb0000000000011110000000000;
		2686: Delta = 25'sb1111111111011110000000000;
		302: Delta = 25'sb0000000001000010000000000;
		1746: Delta = 25'sb1111111111000010000000000;
		1603: Delta = 25'sb0000000000111110000000000;
		3047: Delta = 25'sb1111111110111110000000000;
		2929: Delta = 25'sb0000000010000010000000000;
		2468: Delta = 25'sb1111111110000010000000000;
		881: Delta = 25'sb0000000001111110000000000;
		420: Delta = 25'sb1111111101111110000000000;
		1485: Delta = 25'sb0000000100000010000000000;
		563: Delta = 25'sb1111111100000010000000000;
		2786: Delta = 25'sb0000000011111110000000000;
		1864: Delta = 25'sb1111111011111110000000000;
		1946: Delta = 25'sb0000001000000010000000000;
		102: Delta = 25'sb1111111000000010000000000;
		3247: Delta = 25'sb0000000111111110000000000;
		1403: Delta = 25'sb1111110111111110000000000;
		2868: Delta = 25'sb0000010000000010000000000;
		2529: Delta = 25'sb1111110000000010000000000;
		820: Delta = 25'sb0000001111111110000000000;
		481: Delta = 25'sb1111101111111110000000000;
		1363: Delta = 25'sb0000100000000010000000000;
		685: Delta = 25'sb1111100000000010000000000;
		2664: Delta = 25'sb0000011111111110000000000;
		1986: Delta = 25'sb1111011111111110000000000;
		1702: Delta = 25'sb0001000000000010000000000;
		346: Delta = 25'sb1111000000000010000000000;
		3003: Delta = 25'sb0000111111111110000000000;
		1647: Delta = 25'sb1110111111111110000000000;
		2380: Delta = 25'sb0010000000000010000000000;
		3017: Delta = 25'sb1110000000000010000000000;
		332: Delta = 25'sb0001111111111110000000000;
		969: Delta = 25'sb1101111111111110000000000;
		387: Delta = 25'sb0100000000000010000000000;
		1661: Delta = 25'sb1100000000000010000000000;
		1688: Delta = 25'sb0011111111111110000000000;
		2962: Delta = 25'sb1011111111111110000000000;
		2795: Delta = 25'sb0000000000001100000000000;
		554: Delta = 25'sb1111111111110100000000000;
		193: Delta = 25'sb0000000000010100000000000;
		3156: Delta = 25'sb1111111111101100000000000;
		1687: Delta = 25'sb0000000000100100000000000;
		2409: Delta = 25'sb1111111111100100000000000;
		940: Delta = 25'sb0000000000011100000000000;
		1662: Delta = 25'sb1111111111011100000000000;
		1326: Delta = 25'sb0000000001000100000000000;
		2770: Delta = 25'sb1111111111000100000000000;
		579: Delta = 25'sb0000000000111100000000000;
		2023: Delta = 25'sb1111111110111100000000000;
		604: Delta = 25'sb0000000010000100000000000;
		143: Delta = 25'sb1111111110000100000000000;
		3206: Delta = 25'sb0000000001111100000000000;
		2745: Delta = 25'sb1111111101111100000000000;
		2509: Delta = 25'sb0000000100000100000000000;
		1587: Delta = 25'sb1111111100000100000000000;
		1762: Delta = 25'sb0000000011111100000000000;
		840: Delta = 25'sb1111111011111100000000000;
		2970: Delta = 25'sb0000001000000100000000000;
		1126: Delta = 25'sb1111111000000100000000000;
		2223: Delta = 25'sb0000000111111100000000000;
		379: Delta = 25'sb1111110111111100000000000;
		543: Delta = 25'sb0000010000000100000000000;
		204: Delta = 25'sb1111110000000100000000000;
		3145: Delta = 25'sb0000001111111100000000000;
		2806: Delta = 25'sb1111101111111100000000000;
		2387: Delta = 25'sb0000100000000100000000000;
		1709: Delta = 25'sb1111100000000100000000000;
		1640: Delta = 25'sb0000011111111100000000000;
		962: Delta = 25'sb1111011111111100000000000;
		2726: Delta = 25'sb0001000000000100000000000;
		1370: Delta = 25'sb1111000000000100000000000;
		1979: Delta = 25'sb0000111111111100000000000;
		623: Delta = 25'sb1110111111111100000000000;
		55: Delta = 25'sb0010000000000100000000000;
		692: Delta = 25'sb1110000000000100000000000;
		2657: Delta = 25'sb0001111111111100000000000;
		3294: Delta = 25'sb1101111111111100000000000;
		1411: Delta = 25'sb0100000000000100000000000;
		2685: Delta = 25'sb1100000000000100000000000;
		664: Delta = 25'sb0011111111111100000000000;
		1938: Delta = 25'sb1011111111111100000000000;
		2241: Delta = 25'sb0000000000011000000000000;
		1108: Delta = 25'sb1111111111101000000000000;
		386: Delta = 25'sb0000000000101000000000000;
		2963: Delta = 25'sb1111111111011000000000000;
		25: Delta = 25'sb0000000001001000000000000;
		1469: Delta = 25'sb1111111111001000000000000;
		1880: Delta = 25'sb0000000000111000000000000;
		3324: Delta = 25'sb1111111110111000000000000;
		2652: Delta = 25'sb0000000010001000000000000;
		2191: Delta = 25'sb1111111110001000000000000;
		1158: Delta = 25'sb0000000001111000000000000;
		697: Delta = 25'sb1111111101111000000000000;
		1208: Delta = 25'sb0000000100001000000000000;
		286: Delta = 25'sb1111111100001000000000000;
		3063: Delta = 25'sb0000000011111000000000000;
		2141: Delta = 25'sb1111111011111000000000000;
		1669: Delta = 25'sb0000001000001000000000000;
		3174: Delta = 25'sb1111111000001000000000000;
		175: Delta = 25'sb0000000111111000000000000;
		1680: Delta = 25'sb1111110111111000000000000;
		2591: Delta = 25'sb0000010000001000000000000;
		2252: Delta = 25'sb1111110000001000000000000;
		1097: Delta = 25'sb0000001111111000000000000;
		758: Delta = 25'sb1111101111111000000000000;
		1086: Delta = 25'sb0000100000001000000000000;
		408: Delta = 25'sb1111100000001000000000000;
		2941: Delta = 25'sb0000011111111000000000000;
		2263: Delta = 25'sb1111011111111000000000000;
		1425: Delta = 25'sb0001000000001000000000000;
		69: Delta = 25'sb1111000000001000000000000;
		3280: Delta = 25'sb0000111111111000000000000;
		1924: Delta = 25'sb1110111111111000000000000;
		2103: Delta = 25'sb0010000000001000000000000;
		2740: Delta = 25'sb1110000000001000000000000;
		609: Delta = 25'sb0001111111111000000000000;
		1246: Delta = 25'sb1101111111111000000000000;
		110: Delta = 25'sb0100000000001000000000000;
		1384: Delta = 25'sb1100000000001000000000000;
		1965: Delta = 25'sb0011111111111000000000000;
		3239: Delta = 25'sb1011111111111000000000000;
		1133: Delta = 25'sb0000000000110000000000000;
		2216: Delta = 25'sb1111111111010000000000000;
		772: Delta = 25'sb0000000001010000000000000;
		2577: Delta = 25'sb1111111110110000000000000;
		50: Delta = 25'sb0000000010010000000000000;
		2938: Delta = 25'sb1111111110010000000000000;
		411: Delta = 25'sb0000000001110000000000000;
		3299: Delta = 25'sb1111111101110000000000000;
		1955: Delta = 25'sb0000000100010000000000000;
		1033: Delta = 25'sb1111111100010000000000000;
		2316: Delta = 25'sb0000000011110000000000000;
		1394: Delta = 25'sb1111111011110000000000000;
		2416: Delta = 25'sb0000001000010000000000000;
		572: Delta = 25'sb1111111000010000000000000;
		2777: Delta = 25'sb0000000111110000000000000;
		933: Delta = 25'sb1111110111110000000000000;
		3338: Delta = 25'sb0000010000010000000000000;
		2999: Delta = 25'sb1111110000010000000000000;
		350: Delta = 25'sb0000001111110000000000000;
		11: Delta = 25'sb1111101111110000000000000;
		1833: Delta = 25'sb0000100000010000000000000;
		1155: Delta = 25'sb1111100000010000000000000;
		2194: Delta = 25'sb0000011111110000000000000;
		1516: Delta = 25'sb1111011111110000000000000;
		2172: Delta = 25'sb0001000000010000000000000;
		816: Delta = 25'sb1111000000010000000000000;
		2533: Delta = 25'sb0000111111110000000000000;
		1177: Delta = 25'sb1110111111110000000000000;
		2850: Delta = 25'sb0010000000010000000000000;
		138: Delta = 25'sb1110000000010000000000000;
		3211: Delta = 25'sb0001111111110000000000000;
		499: Delta = 25'sb1101111111110000000000000;
		857: Delta = 25'sb0100000000010000000000000;
		2131: Delta = 25'sb1100000000010000000000000;
		1218: Delta = 25'sb0011111111110000000000000;
		2492: Delta = 25'sb1011111111110000000000000;
		2266: Delta = 25'sb0000000001100000000000000;
		1083: Delta = 25'sb1111111110100000000000000;
		1544: Delta = 25'sb0000000010100000000000000;
		1805: Delta = 25'sb1111111101100000000000000;
		100: Delta = 25'sb0000000100100000000000000;
		2527: Delta = 25'sb1111111100100000000000000;
		822: Delta = 25'sb0000000011100000000000000;
		3249: Delta = 25'sb1111111011100000000000000;
		561: Delta = 25'sb0000001000100000000000000;
		2066: Delta = 25'sb1111111000100000000000000;
		1283: Delta = 25'sb0000000111100000000000000;
		2788: Delta = 25'sb1111110111100000000000000;
		1483: Delta = 25'sb0000010000100000000000000;
		1144: Delta = 25'sb1111110000100000000000000;
		2205: Delta = 25'sb0000001111100000000000000;
		1866: Delta = 25'sb1111101111100000000000000;
		3327: Delta = 25'sb0000100000100000000000000;
		2649: Delta = 25'sb1111100000100000000000000;
		700: Delta = 25'sb0000011111100000000000000;
		22: Delta = 25'sb1111011111100000000000000;
		317: Delta = 25'sb0001000000100000000000000;
		2310: Delta = 25'sb1111000000100000000000000;
		1039: Delta = 25'sb0000111111100000000000000;
		3032: Delta = 25'sb1110111111100000000000000;
		995: Delta = 25'sb0010000000100000000000000;
		1632: Delta = 25'sb1110000000100000000000000;
		1717: Delta = 25'sb0001111111100000000000000;
		2354: Delta = 25'sb1101111111100000000000000;
		2351: Delta = 25'sb0100000000100000000000000;
		276: Delta = 25'sb1100000000100000000000000;
		3073: Delta = 25'sb0011111111100000000000000;
		998: Delta = 25'sb1011111111100000000000000;
		1183: Delta = 25'sb0000000011000000000000000;
		2166: Delta = 25'sb1111111101000000000000000;
		3088: Delta = 25'sb0000000101000000000000000;
		261: Delta = 25'sb1111111011000000000000000;
		200: Delta = 25'sb0000001001000000000000000;
		1705: Delta = 25'sb1111111001000000000000000;
		1644: Delta = 25'sb0000000111000000000000000;
		3149: Delta = 25'sb1111110111000000000000000;
		1122: Delta = 25'sb0000010001000000000000000;
		783: Delta = 25'sb1111110001000000000000000;
		2566: Delta = 25'sb0000001111000000000000000;
		2227: Delta = 25'sb1111101111000000000000000;
		2966: Delta = 25'sb0000100001000000000000000;
		2288: Delta = 25'sb1111100001000000000000000;
		1061: Delta = 25'sb0000011111000000000000000;
		383: Delta = 25'sb1111011111000000000000000;
		3305: Delta = 25'sb0001000001000000000000000;
		1949: Delta = 25'sb1111000001000000000000000;
		1400: Delta = 25'sb0000111111000000000000000;
		44: Delta = 25'sb1110111111000000000000000;
		634: Delta = 25'sb0010000001000000000000000;
		1271: Delta = 25'sb1110000001000000000000000;
		2078: Delta = 25'sb0001111111000000000000000;
		2715: Delta = 25'sb1101111111000000000000000;
		1990: Delta = 25'sb0100000001000000000000000;
		3264: Delta = 25'sb1100000001000000000000000;
		85: Delta = 25'sb0011111111000000000000000;
		1359: Delta = 25'sb1011111111000000000000000;
		2366: Delta = 25'sb0000000110000000000000000;
		983: Delta = 25'sb1111111010000000000000000;
		2827: Delta = 25'sb0000001010000000000000000;
		522: Delta = 25'sb1111110110000000000000000;
		400: Delta = 25'sb0000010010000000000000000;
		61: Delta = 25'sb1111110010000000000000000;
		3288: Delta = 25'sb0000001110000000000000000;
		2949: Delta = 25'sb1111101110000000000000000;
		2244: Delta = 25'sb0000100010000000000000000;
		1566: Delta = 25'sb1111100010000000000000000;
		1783: Delta = 25'sb0000011110000000000000000;
		1105: Delta = 25'sb1111011110000000000000000;
		2583: Delta = 25'sb0001000010000000000000000;
		1227: Delta = 25'sb1111000010000000000000000;
		2122: Delta = 25'sb0000111110000000000000000;
		766: Delta = 25'sb1110111110000000000000000;
		3261: Delta = 25'sb0010000010000000000000000;
		549: Delta = 25'sb1110000010000000000000000;
		2800: Delta = 25'sb0001111110000000000000000;
		88: Delta = 25'sb1101111110000000000000000;
		1268: Delta = 25'sb0100000010000000000000000;
		2542: Delta = 25'sb1100000010000000000000000;
		807: Delta = 25'sb0011111110000000000000000;
		2081: Delta = 25'sb1011111110000000000000000;
		1383: Delta = 25'sb0000001100000000000000000;
		1966: Delta = 25'sb1111110100000000000000000;
		2305: Delta = 25'sb0000010100000000000000000;
		1044: Delta = 25'sb1111101100000000000000000;
		800: Delta = 25'sb0000100100000000000000000;
		122: Delta = 25'sb1111100100000000000000000;
		3227: Delta = 25'sb0000011100000000000000000;
		2549: Delta = 25'sb1111011100000000000000000;
		1139: Delta = 25'sb0001000100000000000000000;
		3132: Delta = 25'sb1111000100000000000000000;
		217: Delta = 25'sb0000111100000000000000000;
		2210: Delta = 25'sb1110111100000000000000000;
		1817: Delta = 25'sb0010000100000000000000000;
		2454: Delta = 25'sb1110000100000000000000000;
		895: Delta = 25'sb0001111100000000000000000;
		1532: Delta = 25'sb1101111100000000000000000;
		3173: Delta = 25'sb0100000100000000000000000;
		1098: Delta = 25'sb1100000100000000000000000;
		2251: Delta = 25'sb0011111100000000000000000;
		176: Delta = 25'sb1011111100000000000000000;
		2766: Delta = 25'sb0000011000000000000000000;
		583: Delta = 25'sb1111101000000000000000000;
		1261: Delta = 25'sb0000101000000000000000000;
		2088: Delta = 25'sb1111011000000000000000000;
		1600: Delta = 25'sb0001001000000000000000000;
		244: Delta = 25'sb1111001000000000000000000;
		3105: Delta = 25'sb0000111000000000000000000;
		1749: Delta = 25'sb1110111000000000000000000;
		2278: Delta = 25'sb0010001000000000000000000;
		2915: Delta = 25'sb1110001000000000000000000;
		434: Delta = 25'sb0001111000000000000000000;
		1071: Delta = 25'sb1101111000000000000000000;
		285: Delta = 25'sb0100001000000000000000000;
		1559: Delta = 25'sb1100001000000000000000000;
		1790: Delta = 25'sb0011111000000000000000000;
		3064: Delta = 25'sb1011111000000000000000000;
		2183: Delta = 25'sb0000110000000000000000000;
		1166: Delta = 25'sb1111010000000000000000000;
		2522: Delta = 25'sb0001010000000000000000000;
		827: Delta = 25'sb1110110000000000000000000;
		3200: Delta = 25'sb0010010000000000000000000;
		488: Delta = 25'sb1110010000000000000000000;
		2861: Delta = 25'sb0001110000000000000000000;
		149: Delta = 25'sb1101110000000000000000000;
		1207: Delta = 25'sb0100010000000000000000000;
		2481: Delta = 25'sb1100010000000000000000000;
		868: Delta = 25'sb0011110000000000000000000;
		2142: Delta = 25'sb1011110000000000000000000;
		1017: Delta = 25'sb0001100000000000000000000;
		2332: Delta = 25'sb1110100000000000000000000;
		1695: Delta = 25'sb0010100000000000000000000;
		1654: Delta = 25'sb1101100000000000000000000;
		3051: Delta = 25'sb0100100000000000000000000;
		976: Delta = 25'sb1100100000000000000000000;
		2373: Delta = 25'sb0011100000000000000000000;
		298: Delta = 25'sb1011100000000000000000000;
		2034: Delta = 25'sb0011000000000000000000000;
		1315: Delta = 25'sb1101000000000000000000000;
		41: Delta = 25'sb0101000000000000000000000;
		3308: Delta = 25'sb1011000000000000000000000;
		719: Delta = 25'sb0110000000000000000000000;
		2630: Delta = 25'sb1010000000000000000000000;
		default: Delta =25'sb0;
	endcase
end

assign N = (W - Delta) / A;

endmodule

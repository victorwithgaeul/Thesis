// Product (AN) Code SEC_LUT_Decoder
// SEC_LUT_Decoder12bits.v
// Received codeword W = AN + e, e is single arithmetic weight error (AWE), +2^i or -2^i.
module SEC_LUT_Decoder12bits(W, N);
input 	[23:0]	W;
output	[11:0]	N;
parameter A = 3349;

wire 	[11:0]	Q;
wire 	[11:0]	R;
assign Q = W / A;
assign R = W - (A * Q);

reg	signed	[24:0]	Delta;
always@(*) begin
	case(R)
		1: Delta = 25'sb0000000000000000000000001;
		3348: Delta = 25'sb1111111111111111111111111;
		2: Delta = 25'sb0000000000000000000000010;
		3347: Delta = 25'sb1111111111111111111111110;
		4: Delta = 25'sb0000000000000000000000100;
		3345: Delta = 25'sb1111111111111111111111100;
		8: Delta = 25'sb0000000000000000000001000;
		3341: Delta = 25'sb1111111111111111111111000;
		16: Delta = 25'sb0000000000000000000010000;
		3333: Delta = 25'sb1111111111111111111110000;
		32: Delta = 25'sb0000000000000000000100000;
		3317: Delta = 25'sb1111111111111111111100000;
		64: Delta = 25'sb0000000000000000001000000;
		3285: Delta = 25'sb1111111111111111111000000;
		128: Delta = 25'sb0000000000000000010000000;
		3221: Delta = 25'sb1111111111111111110000000;
		256: Delta = 25'sb0000000000000000100000000;
		3093: Delta = 25'sb1111111111111111100000000;
		512: Delta = 25'sb0000000000000001000000000;
		2837: Delta = 25'sb1111111111111111000000000;
		1024: Delta = 25'sb0000000000000010000000000;
		2325: Delta = 25'sb1111111111111110000000000;
		2048: Delta = 25'sb0000000000000100000000000;
		1301: Delta = 25'sb1111111111111100000000000;
		747: Delta = 25'sb0000000000001000000000000;
		2602: Delta = 25'sb1111111111111000000000000;
		1494: Delta = 25'sb0000000000010000000000000;
		1855: Delta = 25'sb1111111111110000000000000;
		2988: Delta = 25'sb0000000000100000000000000;
		361: Delta = 25'sb1111111111100000000000000;
		2627: Delta = 25'sb0000000001000000000000000;
		722: Delta = 25'sb1111111111000000000000000;
		1905: Delta = 25'sb0000000010000000000000000;
		1444: Delta = 25'sb1111111110000000000000000;
		461: Delta = 25'sb0000000100000000000000000;
		2888: Delta = 25'sb1111111100000000000000000;
		922: Delta = 25'sb0000001000000000000000000;
		2427: Delta = 25'sb1111111000000000000000000;
		1844: Delta = 25'sb0000010000000000000000000;
		1505: Delta = 25'sb1111110000000000000000000;
		339: Delta = 25'sb0000100000000000000000000;
		3010: Delta = 25'sb1111100000000000000000000;
		678: Delta = 25'sb0001000000000000000000000;
		2671: Delta = 25'sb1111000000000000000000000;
		1356: Delta = 25'sb0010000000000000000000000;
		1993: Delta = 25'sb1110000000000000000000000;
		2712: Delta = 25'sb0100000000000000000000000;
		637: Delta = 25'sb1100000000000000000000000;
		default: Delta =25'sb0;
	endcase
end

assign N = (W - Delta) / A;

endmodule

// Product (AN) Code SEC_LUT_Decoder
// SEC_LUT_Decoder8bits.v
// Received codeword W = AN + e, e is single arithmetic weight error (AWE), +2^i or -2^i.
module SEC_LUT_Decoder8bits(W, N);
input 	[18:0]	W;
output	[7:0]	N;
parameter A = 1939;

wire 	[7:0]	Q;
wire 	[10:0]	R;
assign Q = W / A;
assign R = W - (A * Q);

reg	signed	[19:0]	Delta;
always@(*) begin
	case(R)
		1: Delta = 20'sb00000000000000000001;
		1938: Delta = 20'sb11111111111111111111;
		2: Delta = 20'sb00000000000000000010;
		1937: Delta = 20'sb11111111111111111110;
		4: Delta = 20'sb00000000000000000100;
		1935: Delta = 20'sb11111111111111111100;
		8: Delta = 20'sb00000000000000001000;
		1931: Delta = 20'sb11111111111111111000;
		16: Delta = 20'sb00000000000000010000;
		1923: Delta = 20'sb11111111111111110000;
		32: Delta = 20'sb00000000000000100000;
		1907: Delta = 20'sb11111111111111100000;
		64: Delta = 20'sb00000000000001000000;
		1875: Delta = 20'sb11111111111111000000;
		128: Delta = 20'sb00000000000010000000;
		1811: Delta = 20'sb11111111111110000000;
		256: Delta = 20'sb00000000000100000000;
		1683: Delta = 20'sb11111111111100000000;
		512: Delta = 20'sb00000000001000000000;
		1427: Delta = 20'sb11111111111000000000;
		1024: Delta = 20'sb00000000010000000000;
		915: Delta = 20'sb11111111110000000000;
		109: Delta = 20'sb00000000100000000000;
		1830: Delta = 20'sb11111111100000000000;
		218: Delta = 20'sb00000001000000000000;
		1721: Delta = 20'sb11111111000000000000;
		436: Delta = 20'sb00000010000000000000;
		1503: Delta = 20'sb11111110000000000000;
		872: Delta = 20'sb00000100000000000000;
		1067: Delta = 20'sb11111100000000000000;
		1744: Delta = 20'sb00001000000000000000;
		195: Delta = 20'sb11111000000000000000;
		1549: Delta = 20'sb00010000000000000000;
		390: Delta = 20'sb11110000000000000000;
		1159: Delta = 20'sb00100000000000000000;
		780: Delta = 20'sb11100000000000000000;
		379: Delta = 20'sb01000000000000000000;
		1560: Delta = 20'sb11000000000000000000;
		default: Delta =20'sb0;
	endcase
end

assign N = (W - Delta) / A;

endmodule

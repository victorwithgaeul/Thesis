// Product (AN) Code SEC r-LUT
// SEC_rLUT30bits.v
// Received remainder r, output single error location.
module SEC_rLUT30bits(r, l);
input 	[14:0]	r;
output	reg	signed	[6:0]	l;
always@(*) begin
	case(r)
		1: l = +1;
		18612: l = -1;
		2: l = +2;
		18611: l = -2;
		4: l = +3;
		18609: l = -3;
		8: l = +4;
		18605: l = -4;
		16: l = +5;
		18597: l = -5;
		32: l = +6;
		18581: l = -6;
		64: l = +7;
		18549: l = -7;
		128: l = +8;
		18485: l = -8;
		256: l = +9;
		18357: l = -9;
		512: l = +10;
		18101: l = -10;
		1024: l = +11;
		17589: l = -11;
		2048: l = +12;
		16565: l = -12;
		4096: l = +13;
		14517: l = -13;
		8192: l = +14;
		10421: l = -14;
		16384: l = +15;
		2229: l = -15;
		14155: l = +16;
		4458: l = -16;
		9697: l = +17;
		8916: l = -17;
		781: l = +18;
		17832: l = -18;
		1562: l = +19;
		17051: l = -19;
		3124: l = +20;
		15489: l = -20;
		6248: l = +21;
		12365: l = -21;
		12496: l = +22;
		6117: l = -22;
		6379: l = +23;
		12234: l = -23;
		12758: l = +24;
		5855: l = -24;
		6903: l = +25;
		11710: l = -25;
		13806: l = +26;
		4807: l = -26;
		8999: l = +27;
		9614: l = -27;
		17998: l = +28;
		615: l = -28;
		17383: l = +29;
		1230: l = -29;
		16153: l = +30;
		2460: l = -30;
		13693: l = +31;
		4920: l = -31;
		8773: l = +32;
		9840: l = -32;
		17546: l = +33;
		1067: l = -33;
		16479: l = +34;
		2134: l = -34;
		14345: l = +35;
		4268: l = -35;
		10077: l = +36;
		8536: l = -36;
		1541: l = +37;
		17072: l = -37;
		3082: l = +38;
		15531: l = -38;
		6164: l = +39;
		12449: l = -39;
		12328: l = +40;
		6285: l = -40;
		6043: l = +41;
		12570: l = -41;
		12086: l = +42;
		6527: l = -42;
		5559: l = +43;
		13054: l = -43;
		11118: l = +44;
		7495: l = -44;
		3623: l = +45;
		14990: l = -45;
		default: l = 0;
	endcase
end

endmodule

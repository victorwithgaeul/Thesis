// Product (AN) Code SEC l-LUT
// SEC_lLUT30bits.v
// Received single error location l, output remainder r.
module SEC_lLUT30bits(l, r);
input	signed	[6:0]	l;
output	reg	[14:0]	r;
always@(*) begin
	case(l)
		1: r = 1;
		-1: r = 18612;
		2: r = 2;
		-2: r = 18611;
		3: r = 4;
		-3: r = 18609;
		4: r = 8;
		-4: r = 18605;
		5: r = 16;
		-5: r = 18597;
		6: r = 32;
		-6: r = 18581;
		7: r = 64;
		-7: r = 18549;
		8: r = 128;
		-8: r = 18485;
		9: r = 256;
		-9: r = 18357;
		10: r = 512;
		-10: r = 18101;
		11: r = 1024;
		-11: r = 17589;
		12: r = 2048;
		-12: r = 16565;
		13: r = 4096;
		-13: r = 14517;
		14: r = 8192;
		-14: r = 10421;
		15: r = 16384;
		-15: r = 2229;
		16: r = 14155;
		-16: r = 4458;
		17: r = 9697;
		-17: r = 8916;
		18: r = 781;
		-18: r = 17832;
		19: r = 1562;
		-19: r = 17051;
		20: r = 3124;
		-20: r = 15489;
		21: r = 6248;
		-21: r = 12365;
		22: r = 12496;
		-22: r = 6117;
		23: r = 6379;
		-23: r = 12234;
		24: r = 12758;
		-24: r = 5855;
		25: r = 6903;
		-25: r = 11710;
		26: r = 13806;
		-26: r = 4807;
		27: r = 8999;
		-27: r = 9614;
		28: r = 17998;
		-28: r = 615;
		29: r = 17383;
		-29: r = 1230;
		30: r = 16153;
		-30: r = 2460;
		31: r = 13693;
		-31: r = 4920;
		32: r = 8773;
		-32: r = 9840;
		33: r = 17546;
		-33: r = 1067;
		34: r = 16479;
		-34: r = 2134;
		35: r = 14345;
		-35: r = 4268;
		36: r = 10077;
		-36: r = 8536;
		37: r = 1541;
		-37: r = 17072;
		38: r = 3082;
		-38: r = 15531;
		39: r = 6164;
		-39: r = 12449;
		40: r = 12328;
		-40: r = 6285;
		41: r = 6043;
		-41: r = 12570;
		42: r = 12086;
		-42: r = 6527;
		43: r = 5559;
		-43: r = 13054;
		44: r = 11118;
		-44: r = 7495;
		45: r = 3623;
		-45: r = 14990;
		default: r = 0;
	endcase
end

endmodule

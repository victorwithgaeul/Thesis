// Product (AN) Code DEC_LUT_Decoder
// DEC_LUT_Decoder30bits.v
// Received codeword W = AN + E, E is double AWE (E = e1 + e2), +2^i or -2^i.
module DEC_LUT_Decoder30bits_clk(clk, rst_n, W, found, N);

//=========================================================================
//   PARAMETER AND LOCALPARAM FOR FSM
//   W_BITS 要考慮 OVERFLOW 問題
//   N_BITS 也要考慮 OVERFLOW 問題
//=========================================================================
parameter A = 18613 , W_BITS = 46, A_BITS = 15 , N_BITS = 31;

localparam [1:0] idle=2'b00, pre=2'b01,load=2'b10, LUT=2'b11;

reg [1:0] ps;
//==========================================
//   INPUT AND OUTPUT DECLARATION
//==========================================
input   clk, rst_n;
input 	[W_BITS-1:0]	W;
output	reg  [N_BITS-1:0] N;
output  reg  found;

reg 	[N_BITS-1:0]	Q;
reg 	[A_BITS-1:0]	R;

reg	signed	[45:0]	Delta;
always@(*) begin
	case(R)
		1: Delta = 46'sb0000000000000000000000000000000000000000000001;
		18612: Delta = 46'sb1111111111111111111111111111111111111111111111;
		2: Delta = 46'sb0000000000000000000000000000000000000000000010;
		18611: Delta = 46'sb1111111111111111111111111111111111111111111110;
		4: Delta = 46'sb0000000000000000000000000000000000000000000100;
		18609: Delta = 46'sb1111111111111111111111111111111111111111111100;
		8: Delta = 46'sb0000000000000000000000000000000000000000001000;
		18605: Delta = 46'sb1111111111111111111111111111111111111111111000;
		16: Delta = 46'sb0000000000000000000000000000000000000000010000;
		18597: Delta = 46'sb1111111111111111111111111111111111111111110000;
		32: Delta = 46'sb0000000000000000000000000000000000000000100000;
		18581: Delta = 46'sb1111111111111111111111111111111111111111100000;
		64: Delta = 46'sb0000000000000000000000000000000000000001000000;
		18549: Delta = 46'sb1111111111111111111111111111111111111111000000;
		128: Delta = 46'sb0000000000000000000000000000000000000010000000;
		18485: Delta = 46'sb1111111111111111111111111111111111111110000000;
		256: Delta = 46'sb0000000000000000000000000000000000000100000000;
		18357: Delta = 46'sb1111111111111111111111111111111111111100000000;
		512: Delta = 46'sb0000000000000000000000000000000000001000000000;
		18101: Delta = 46'sb1111111111111111111111111111111111111000000000;
		1024: Delta = 46'sb0000000000000000000000000000000000010000000000;
		17589: Delta = 46'sb1111111111111111111111111111111111110000000000;
		2048: Delta = 46'sb0000000000000000000000000000000000100000000000;
		16565: Delta = 46'sb1111111111111111111111111111111111100000000000;
		4096: Delta = 46'sb0000000000000000000000000000000001000000000000;
		14517: Delta = 46'sb1111111111111111111111111111111111000000000000;
		8192: Delta = 46'sb0000000000000000000000000000000010000000000000;
		10421: Delta = 46'sb1111111111111111111111111111111110000000000000;
		16384: Delta = 46'sb0000000000000000000000000000000100000000000000;
		2229: Delta = 46'sb1111111111111111111111111111111100000000000000;
		14155: Delta = 46'sb0000000000000000000000000000001000000000000000;
		4458: Delta = 46'sb1111111111111111111111111111111000000000000000;
		9697: Delta = 46'sb0000000000000000000000000000010000000000000000;
		8916: Delta = 46'sb1111111111111111111111111111110000000000000000;
		781: Delta = 46'sb0000000000000000000000000000100000000000000000;
		17832: Delta = 46'sb1111111111111111111111111111100000000000000000;
		1562: Delta = 46'sb0000000000000000000000000001000000000000000000;
		17051: Delta = 46'sb1111111111111111111111111111000000000000000000;
		3124: Delta = 46'sb0000000000000000000000000010000000000000000000;
		15489: Delta = 46'sb1111111111111111111111111110000000000000000000;
		6248: Delta = 46'sb0000000000000000000000000100000000000000000000;
		12365: Delta = 46'sb1111111111111111111111111100000000000000000000;
		12496: Delta = 46'sb0000000000000000000000001000000000000000000000;
		6117: Delta = 46'sb1111111111111111111111111000000000000000000000;
		6379: Delta = 46'sb0000000000000000000000010000000000000000000000;
		12234: Delta = 46'sb1111111111111111111111110000000000000000000000;
		12758: Delta = 46'sb0000000000000000000000100000000000000000000000;
		5855: Delta = 46'sb1111111111111111111111100000000000000000000000;
		6903: Delta = 46'sb0000000000000000000001000000000000000000000000;
		11710: Delta = 46'sb1111111111111111111111000000000000000000000000;
		13806: Delta = 46'sb0000000000000000000010000000000000000000000000;
		4807: Delta = 46'sb1111111111111111111110000000000000000000000000;
		8999: Delta = 46'sb0000000000000000000100000000000000000000000000;
		9614: Delta = 46'sb1111111111111111111100000000000000000000000000;
		17998: Delta = 46'sb0000000000000000001000000000000000000000000000;
		615: Delta = 46'sb1111111111111111111000000000000000000000000000;
		17383: Delta = 46'sb0000000000000000010000000000000000000000000000;
		1230: Delta = 46'sb1111111111111111110000000000000000000000000000;
		16153: Delta = 46'sb0000000000000000100000000000000000000000000000;
		2460: Delta = 46'sb1111111111111111100000000000000000000000000000;
		13693: Delta = 46'sb0000000000000001000000000000000000000000000000;
		4920: Delta = 46'sb1111111111111111000000000000000000000000000000;
		8773: Delta = 46'sb0000000000000010000000000000000000000000000000;
		9840: Delta = 46'sb1111111111111110000000000000000000000000000000;
		17546: Delta = 46'sb0000000000000100000000000000000000000000000000;
		1067: Delta = 46'sb1111111111111100000000000000000000000000000000;
		16479: Delta = 46'sb0000000000001000000000000000000000000000000000;
		2134: Delta = 46'sb1111111111111000000000000000000000000000000000;
		14345: Delta = 46'sb0000000000010000000000000000000000000000000000;
		4268: Delta = 46'sb1111111111110000000000000000000000000000000000;
		10077: Delta = 46'sb0000000000100000000000000000000000000000000000;
		8536: Delta = 46'sb1111111111100000000000000000000000000000000000;
		1541: Delta = 46'sb0000000001000000000000000000000000000000000000;
		17072: Delta = 46'sb1111111111000000000000000000000000000000000000;
		3082: Delta = 46'sb0000000010000000000000000000000000000000000000;
		15531: Delta = 46'sb1111111110000000000000000000000000000000000000;
		6164: Delta = 46'sb0000000100000000000000000000000000000000000000;
		12449: Delta = 46'sb1111111100000000000000000000000000000000000000;
		12328: Delta = 46'sb0000001000000000000000000000000000000000000000;
		6285: Delta = 46'sb1111111000000000000000000000000000000000000000;
		6043: Delta = 46'sb0000010000000000000000000000000000000000000000;
		12570: Delta = 46'sb1111110000000000000000000000000000000000000000;
		12086: Delta = 46'sb0000100000000000000000000000000000000000000000;
		6527: Delta = 46'sb1111100000000000000000000000000000000000000000;
		5559: Delta = 46'sb0001000000000000000000000000000000000000000000;
		13054: Delta = 46'sb1111000000000000000000000000000000000000000000;
		11118: Delta = 46'sb0010000000000000000000000000000000000000000000;
		7495: Delta = 46'sb1110000000000000000000000000000000000000000000;
		3623: Delta = 46'sb0100000000000000000000000000000000000000000000;
		14990: Delta = 46'sb1100000000000000000000000000000000000000000000;
		3: Delta = 46'sb0000000000000000000000000000000000000000000011;
		18610: Delta = 46'sb1111111111111111111111111111111111111111111101;
		5: Delta = 46'sb0000000000000000000000000000000000000000000101;
		18608: Delta = 46'sb1111111111111111111111111111111111111111111011;
		9: Delta = 46'sb0000000000000000000000000000000000000000001001;
		18606: Delta = 46'sb1111111111111111111111111111111111111111111001;
		7: Delta = 46'sb0000000000000000000000000000000000000000000111;
		18604: Delta = 46'sb1111111111111111111111111111111111111111110111;
		17: Delta = 46'sb0000000000000000000000000000000000000000010001;
		18598: Delta = 46'sb1111111111111111111111111111111111111111110001;
		15: Delta = 46'sb0000000000000000000000000000000000000000001111;
		18596: Delta = 46'sb1111111111111111111111111111111111111111101111;
		33: Delta = 46'sb0000000000000000000000000000000000000000100001;
		18582: Delta = 46'sb1111111111111111111111111111111111111111100001;
		31: Delta = 46'sb0000000000000000000000000000000000000000011111;
		18580: Delta = 46'sb1111111111111111111111111111111111111111011111;
		65: Delta = 46'sb0000000000000000000000000000000000000001000001;
		18550: Delta = 46'sb1111111111111111111111111111111111111111000001;
		63: Delta = 46'sb0000000000000000000000000000000000000000111111;
		18548: Delta = 46'sb1111111111111111111111111111111111111110111111;
		129: Delta = 46'sb0000000000000000000000000000000000000010000001;
		18486: Delta = 46'sb1111111111111111111111111111111111111110000001;
		127: Delta = 46'sb0000000000000000000000000000000000000001111111;
		18484: Delta = 46'sb1111111111111111111111111111111111111101111111;
		257: Delta = 46'sb0000000000000000000000000000000000000100000001;
		18358: Delta = 46'sb1111111111111111111111111111111111111100000001;
		255: Delta = 46'sb0000000000000000000000000000000000000011111111;
		18356: Delta = 46'sb1111111111111111111111111111111111111011111111;
		513: Delta = 46'sb0000000000000000000000000000000000001000000001;
		18102: Delta = 46'sb1111111111111111111111111111111111111000000001;
		511: Delta = 46'sb0000000000000000000000000000000000000111111111;
		18100: Delta = 46'sb1111111111111111111111111111111111110111111111;
		1025: Delta = 46'sb0000000000000000000000000000000000010000000001;
		17590: Delta = 46'sb1111111111111111111111111111111111110000000001;
		1023: Delta = 46'sb0000000000000000000000000000000000001111111111;
		17588: Delta = 46'sb1111111111111111111111111111111111101111111111;
		2049: Delta = 46'sb0000000000000000000000000000000000100000000001;
		16566: Delta = 46'sb1111111111111111111111111111111111100000000001;
		2047: Delta = 46'sb0000000000000000000000000000000000011111111111;
		16564: Delta = 46'sb1111111111111111111111111111111111011111111111;
		4097: Delta = 46'sb0000000000000000000000000000000001000000000001;
		14518: Delta = 46'sb1111111111111111111111111111111111000000000001;
		4095: Delta = 46'sb0000000000000000000000000000000000111111111111;
		14516: Delta = 46'sb1111111111111111111111111111111110111111111111;
		8193: Delta = 46'sb0000000000000000000000000000000010000000000001;
		10422: Delta = 46'sb1111111111111111111111111111111110000000000001;
		8191: Delta = 46'sb0000000000000000000000000000000001111111111111;
		10420: Delta = 46'sb1111111111111111111111111111111101111111111111;
		16385: Delta = 46'sb0000000000000000000000000000000100000000000001;
		2230: Delta = 46'sb1111111111111111111111111111111100000000000001;
		16383: Delta = 46'sb0000000000000000000000000000000011111111111111;
		2228: Delta = 46'sb1111111111111111111111111111111011111111111111;
		14156: Delta = 46'sb0000000000000000000000000000001000000000000001;
		4459: Delta = 46'sb1111111111111111111111111111111000000000000001;
		14154: Delta = 46'sb0000000000000000000000000000000111111111111111;
		4457: Delta = 46'sb1111111111111111111111111111110111111111111111;
		9698: Delta = 46'sb0000000000000000000000000000010000000000000001;
		8917: Delta = 46'sb1111111111111111111111111111110000000000000001;
		9696: Delta = 46'sb0000000000000000000000000000001111111111111111;
		8915: Delta = 46'sb1111111111111111111111111111101111111111111111;
		782: Delta = 46'sb0000000000000000000000000000100000000000000001;
		17833: Delta = 46'sb1111111111111111111111111111100000000000000001;
		780: Delta = 46'sb0000000000000000000000000000011111111111111111;
		17831: Delta = 46'sb1111111111111111111111111111011111111111111111;
		1563: Delta = 46'sb0000000000000000000000000001000000000000000001;
		17052: Delta = 46'sb1111111111111111111111111111000000000000000001;
		1561: Delta = 46'sb0000000000000000000000000000111111111111111111;
		17050: Delta = 46'sb1111111111111111111111111110111111111111111111;
		3125: Delta = 46'sb0000000000000000000000000010000000000000000001;
		15490: Delta = 46'sb1111111111111111111111111110000000000000000001;
		3123: Delta = 46'sb0000000000000000000000000001111111111111111111;
		15488: Delta = 46'sb1111111111111111111111111101111111111111111111;
		6249: Delta = 46'sb0000000000000000000000000100000000000000000001;
		12366: Delta = 46'sb1111111111111111111111111100000000000000000001;
		6247: Delta = 46'sb0000000000000000000000000011111111111111111111;
		12364: Delta = 46'sb1111111111111111111111111011111111111111111111;
		12497: Delta = 46'sb0000000000000000000000001000000000000000000001;
		6118: Delta = 46'sb1111111111111111111111111000000000000000000001;
		12495: Delta = 46'sb0000000000000000000000000111111111111111111111;
		6116: Delta = 46'sb1111111111111111111111110111111111111111111111;
		6380: Delta = 46'sb0000000000000000000000010000000000000000000001;
		12235: Delta = 46'sb1111111111111111111111110000000000000000000001;
		6378: Delta = 46'sb0000000000000000000000001111111111111111111111;
		12233: Delta = 46'sb1111111111111111111111101111111111111111111111;
		12759: Delta = 46'sb0000000000000000000000100000000000000000000001;
		5856: Delta = 46'sb1111111111111111111111100000000000000000000001;
		12757: Delta = 46'sb0000000000000000000000011111111111111111111111;
		5854: Delta = 46'sb1111111111111111111111011111111111111111111111;
		6904: Delta = 46'sb0000000000000000000001000000000000000000000001;
		11711: Delta = 46'sb1111111111111111111111000000000000000000000001;
		6902: Delta = 46'sb0000000000000000000000111111111111111111111111;
		11709: Delta = 46'sb1111111111111111111110111111111111111111111111;
		13807: Delta = 46'sb0000000000000000000010000000000000000000000001;
		4808: Delta = 46'sb1111111111111111111110000000000000000000000001;
		13805: Delta = 46'sb0000000000000000000001111111111111111111111111;
		4806: Delta = 46'sb1111111111111111111101111111111111111111111111;
		9000: Delta = 46'sb0000000000000000000100000000000000000000000001;
		9615: Delta = 46'sb1111111111111111111100000000000000000000000001;
		8998: Delta = 46'sb0000000000000000000011111111111111111111111111;
		9613: Delta = 46'sb1111111111111111111011111111111111111111111111;
		17999: Delta = 46'sb0000000000000000001000000000000000000000000001;
		616: Delta = 46'sb1111111111111111111000000000000000000000000001;
		17997: Delta = 46'sb0000000000000000000111111111111111111111111111;
		614: Delta = 46'sb1111111111111111110111111111111111111111111111;
		17384: Delta = 46'sb0000000000000000010000000000000000000000000001;
		1231: Delta = 46'sb1111111111111111110000000000000000000000000001;
		17382: Delta = 46'sb0000000000000000001111111111111111111111111111;
		1229: Delta = 46'sb1111111111111111101111111111111111111111111111;
		16154: Delta = 46'sb0000000000000000100000000000000000000000000001;
		2461: Delta = 46'sb1111111111111111100000000000000000000000000001;
		16152: Delta = 46'sb0000000000000000011111111111111111111111111111;
		2459: Delta = 46'sb1111111111111111011111111111111111111111111111;
		13694: Delta = 46'sb0000000000000001000000000000000000000000000001;
		4921: Delta = 46'sb1111111111111111000000000000000000000000000001;
		13692: Delta = 46'sb0000000000000000111111111111111111111111111111;
		4919: Delta = 46'sb1111111111111110111111111111111111111111111111;
		8774: Delta = 46'sb0000000000000010000000000000000000000000000001;
		9841: Delta = 46'sb1111111111111110000000000000000000000000000001;
		8772: Delta = 46'sb0000000000000001111111111111111111111111111111;
		9839: Delta = 46'sb1111111111111101111111111111111111111111111111;
		17547: Delta = 46'sb0000000000000100000000000000000000000000000001;
		1068: Delta = 46'sb1111111111111100000000000000000000000000000001;
		17545: Delta = 46'sb0000000000000011111111111111111111111111111111;
		1066: Delta = 46'sb1111111111111011111111111111111111111111111111;
		16480: Delta = 46'sb0000000000001000000000000000000000000000000001;
		2135: Delta = 46'sb1111111111111000000000000000000000000000000001;
		16478: Delta = 46'sb0000000000000111111111111111111111111111111111;
		2133: Delta = 46'sb1111111111110111111111111111111111111111111111;
		14346: Delta = 46'sb0000000000010000000000000000000000000000000001;
		4269: Delta = 46'sb1111111111110000000000000000000000000000000001;
		14344: Delta = 46'sb0000000000001111111111111111111111111111111111;
		4267: Delta = 46'sb1111111111101111111111111111111111111111111111;
		10078: Delta = 46'sb0000000000100000000000000000000000000000000001;
		8537: Delta = 46'sb1111111111100000000000000000000000000000000001;
		10076: Delta = 46'sb0000000000011111111111111111111111111111111111;
		8535: Delta = 46'sb1111111111011111111111111111111111111111111111;
		1542: Delta = 46'sb0000000001000000000000000000000000000000000001;
		17073: Delta = 46'sb1111111111000000000000000000000000000000000001;
		1540: Delta = 46'sb0000000000111111111111111111111111111111111111;
		17071: Delta = 46'sb1111111110111111111111111111111111111111111111;
		3083: Delta = 46'sb0000000010000000000000000000000000000000000001;
		15532: Delta = 46'sb1111111110000000000000000000000000000000000001;
		3081: Delta = 46'sb0000000001111111111111111111111111111111111111;
		15530: Delta = 46'sb1111111101111111111111111111111111111111111111;
		6165: Delta = 46'sb0000000100000000000000000000000000000000000001;
		12450: Delta = 46'sb1111111100000000000000000000000000000000000001;
		6163: Delta = 46'sb0000000011111111111111111111111111111111111111;
		12448: Delta = 46'sb1111111011111111111111111111111111111111111111;
		12329: Delta = 46'sb0000001000000000000000000000000000000000000001;
		6286: Delta = 46'sb1111111000000000000000000000000000000000000001;
		12327: Delta = 46'sb0000000111111111111111111111111111111111111111;
		6284: Delta = 46'sb1111110111111111111111111111111111111111111111;
		6044: Delta = 46'sb0000010000000000000000000000000000000000000001;
		12571: Delta = 46'sb1111110000000000000000000000000000000000000001;
		6042: Delta = 46'sb0000001111111111111111111111111111111111111111;
		12569: Delta = 46'sb1111101111111111111111111111111111111111111111;
		12087: Delta = 46'sb0000100000000000000000000000000000000000000001;
		6528: Delta = 46'sb1111100000000000000000000000000000000000000001;
		12085: Delta = 46'sb0000011111111111111111111111111111111111111111;
		6526: Delta = 46'sb1111011111111111111111111111111111111111111111;
		5560: Delta = 46'sb0001000000000000000000000000000000000000000001;
		13055: Delta = 46'sb1111000000000000000000000000000000000000000001;
		5558: Delta = 46'sb0000111111111111111111111111111111111111111111;
		13053: Delta = 46'sb1110111111111111111111111111111111111111111111;
		11119: Delta = 46'sb0010000000000000000000000000000000000000000001;
		7496: Delta = 46'sb1110000000000000000000000000000000000000000001;
		11117: Delta = 46'sb0001111111111111111111111111111111111111111111;
		7494: Delta = 46'sb1101111111111111111111111111111111111111111111;
		3624: Delta = 46'sb0100000000000000000000000000000000000000000001;
		14991: Delta = 46'sb1100000000000000000000000000000000000000000001;
		3622: Delta = 46'sb0011111111111111111111111111111111111111111111;
		14989: Delta = 46'sb1011111111111111111111111111111111111111111111;
		6: Delta = 46'sb0000000000000000000000000000000000000000000110;
		18607: Delta = 46'sb1111111111111111111111111111111111111111111010;
		10: Delta = 46'sb0000000000000000000000000000000000000000001010;
		18603: Delta = 46'sb1111111111111111111111111111111111111111110110;
		18: Delta = 46'sb0000000000000000000000000000000000000000010010;
		18599: Delta = 46'sb1111111111111111111111111111111111111111110010;
		14: Delta = 46'sb0000000000000000000000000000000000000000001110;
		18595: Delta = 46'sb1111111111111111111111111111111111111111101110;
		34: Delta = 46'sb0000000000000000000000000000000000000000100010;
		18583: Delta = 46'sb1111111111111111111111111111111111111111100010;
		30: Delta = 46'sb0000000000000000000000000000000000000000011110;
		18579: Delta = 46'sb1111111111111111111111111111111111111111011110;
		66: Delta = 46'sb0000000000000000000000000000000000000001000010;
		18551: Delta = 46'sb1111111111111111111111111111111111111111000010;
		62: Delta = 46'sb0000000000000000000000000000000000000000111110;
		18547: Delta = 46'sb1111111111111111111111111111111111111110111110;
		130: Delta = 46'sb0000000000000000000000000000000000000010000010;
		18487: Delta = 46'sb1111111111111111111111111111111111111110000010;
		126: Delta = 46'sb0000000000000000000000000000000000000001111110;
		18483: Delta = 46'sb1111111111111111111111111111111111111101111110;
		258: Delta = 46'sb0000000000000000000000000000000000000100000010;
		18359: Delta = 46'sb1111111111111111111111111111111111111100000010;
		254: Delta = 46'sb0000000000000000000000000000000000000011111110;
		18355: Delta = 46'sb1111111111111111111111111111111111111011111110;
		514: Delta = 46'sb0000000000000000000000000000000000001000000010;
		18103: Delta = 46'sb1111111111111111111111111111111111111000000010;
		510: Delta = 46'sb0000000000000000000000000000000000000111111110;
		18099: Delta = 46'sb1111111111111111111111111111111111110111111110;
		1026: Delta = 46'sb0000000000000000000000000000000000010000000010;
		17591: Delta = 46'sb1111111111111111111111111111111111110000000010;
		1022: Delta = 46'sb0000000000000000000000000000000000001111111110;
		17587: Delta = 46'sb1111111111111111111111111111111111101111111110;
		2050: Delta = 46'sb0000000000000000000000000000000000100000000010;
		16567: Delta = 46'sb1111111111111111111111111111111111100000000010;
		2046: Delta = 46'sb0000000000000000000000000000000000011111111110;
		16563: Delta = 46'sb1111111111111111111111111111111111011111111110;
		4098: Delta = 46'sb0000000000000000000000000000000001000000000010;
		14519: Delta = 46'sb1111111111111111111111111111111111000000000010;
		4094: Delta = 46'sb0000000000000000000000000000000000111111111110;
		14515: Delta = 46'sb1111111111111111111111111111111110111111111110;
		8194: Delta = 46'sb0000000000000000000000000000000010000000000010;
		10423: Delta = 46'sb1111111111111111111111111111111110000000000010;
		8190: Delta = 46'sb0000000000000000000000000000000001111111111110;
		10419: Delta = 46'sb1111111111111111111111111111111101111111111110;
		16386: Delta = 46'sb0000000000000000000000000000000100000000000010;
		2231: Delta = 46'sb1111111111111111111111111111111100000000000010;
		16382: Delta = 46'sb0000000000000000000000000000000011111111111110;
		2227: Delta = 46'sb1111111111111111111111111111111011111111111110;
		14157: Delta = 46'sb0000000000000000000000000000001000000000000010;
		4460: Delta = 46'sb1111111111111111111111111111111000000000000010;
		14153: Delta = 46'sb0000000000000000000000000000000111111111111110;
		4456: Delta = 46'sb1111111111111111111111111111110111111111111110;
		9699: Delta = 46'sb0000000000000000000000000000010000000000000010;
		8918: Delta = 46'sb1111111111111111111111111111110000000000000010;
		9695: Delta = 46'sb0000000000000000000000000000001111111111111110;
		8914: Delta = 46'sb1111111111111111111111111111101111111111111110;
		783: Delta = 46'sb0000000000000000000000000000100000000000000010;
		17834: Delta = 46'sb1111111111111111111111111111100000000000000010;
		779: Delta = 46'sb0000000000000000000000000000011111111111111110;
		17830: Delta = 46'sb1111111111111111111111111111011111111111111110;
		1564: Delta = 46'sb0000000000000000000000000001000000000000000010;
		17053: Delta = 46'sb1111111111111111111111111111000000000000000010;
		1560: Delta = 46'sb0000000000000000000000000000111111111111111110;
		17049: Delta = 46'sb1111111111111111111111111110111111111111111110;
		3126: Delta = 46'sb0000000000000000000000000010000000000000000010;
		15491: Delta = 46'sb1111111111111111111111111110000000000000000010;
		3122: Delta = 46'sb0000000000000000000000000001111111111111111110;
		15487: Delta = 46'sb1111111111111111111111111101111111111111111110;
		6250: Delta = 46'sb0000000000000000000000000100000000000000000010;
		12367: Delta = 46'sb1111111111111111111111111100000000000000000010;
		6246: Delta = 46'sb0000000000000000000000000011111111111111111110;
		12363: Delta = 46'sb1111111111111111111111111011111111111111111110;
		12498: Delta = 46'sb0000000000000000000000001000000000000000000010;
		6119: Delta = 46'sb1111111111111111111111111000000000000000000010;
		12494: Delta = 46'sb0000000000000000000000000111111111111111111110;
		6115: Delta = 46'sb1111111111111111111111110111111111111111111110;
		6381: Delta = 46'sb0000000000000000000000010000000000000000000010;
		12236: Delta = 46'sb1111111111111111111111110000000000000000000010;
		6377: Delta = 46'sb0000000000000000000000001111111111111111111110;
		12232: Delta = 46'sb1111111111111111111111101111111111111111111110;
		12760: Delta = 46'sb0000000000000000000000100000000000000000000010;
		5857: Delta = 46'sb1111111111111111111111100000000000000000000010;
		12756: Delta = 46'sb0000000000000000000000011111111111111111111110;
		5853: Delta = 46'sb1111111111111111111111011111111111111111111110;
		6905: Delta = 46'sb0000000000000000000001000000000000000000000010;
		11712: Delta = 46'sb1111111111111111111111000000000000000000000010;
		6901: Delta = 46'sb0000000000000000000000111111111111111111111110;
		11708: Delta = 46'sb1111111111111111111110111111111111111111111110;
		13808: Delta = 46'sb0000000000000000000010000000000000000000000010;
		4809: Delta = 46'sb1111111111111111111110000000000000000000000010;
		13804: Delta = 46'sb0000000000000000000001111111111111111111111110;
		4805: Delta = 46'sb1111111111111111111101111111111111111111111110;
		9001: Delta = 46'sb0000000000000000000100000000000000000000000010;
		9616: Delta = 46'sb1111111111111111111100000000000000000000000010;
		8997: Delta = 46'sb0000000000000000000011111111111111111111111110;
		9612: Delta = 46'sb1111111111111111111011111111111111111111111110;
		18000: Delta = 46'sb0000000000000000001000000000000000000000000010;
		617: Delta = 46'sb1111111111111111111000000000000000000000000010;
		17996: Delta = 46'sb0000000000000000000111111111111111111111111110;
		613: Delta = 46'sb1111111111111111110111111111111111111111111110;
		17385: Delta = 46'sb0000000000000000010000000000000000000000000010;
		1232: Delta = 46'sb1111111111111111110000000000000000000000000010;
		17381: Delta = 46'sb0000000000000000001111111111111111111111111110;
		1228: Delta = 46'sb1111111111111111101111111111111111111111111110;
		16155: Delta = 46'sb0000000000000000100000000000000000000000000010;
		2462: Delta = 46'sb1111111111111111100000000000000000000000000010;
		16151: Delta = 46'sb0000000000000000011111111111111111111111111110;
		2458: Delta = 46'sb1111111111111111011111111111111111111111111110;
		13695: Delta = 46'sb0000000000000001000000000000000000000000000010;
		4922: Delta = 46'sb1111111111111111000000000000000000000000000010;
		13691: Delta = 46'sb0000000000000000111111111111111111111111111110;
		4918: Delta = 46'sb1111111111111110111111111111111111111111111110;
		8775: Delta = 46'sb0000000000000010000000000000000000000000000010;
		9842: Delta = 46'sb1111111111111110000000000000000000000000000010;
		8771: Delta = 46'sb0000000000000001111111111111111111111111111110;
		9838: Delta = 46'sb1111111111111101111111111111111111111111111110;
		17548: Delta = 46'sb0000000000000100000000000000000000000000000010;
		1069: Delta = 46'sb1111111111111100000000000000000000000000000010;
		17544: Delta = 46'sb0000000000000011111111111111111111111111111110;
		1065: Delta = 46'sb1111111111111011111111111111111111111111111110;
		16481: Delta = 46'sb0000000000001000000000000000000000000000000010;
		2136: Delta = 46'sb1111111111111000000000000000000000000000000010;
		16477: Delta = 46'sb0000000000000111111111111111111111111111111110;
		2132: Delta = 46'sb1111111111110111111111111111111111111111111110;
		14347: Delta = 46'sb0000000000010000000000000000000000000000000010;
		4270: Delta = 46'sb1111111111110000000000000000000000000000000010;
		14343: Delta = 46'sb0000000000001111111111111111111111111111111110;
		4266: Delta = 46'sb1111111111101111111111111111111111111111111110;
		10079: Delta = 46'sb0000000000100000000000000000000000000000000010;
		8538: Delta = 46'sb1111111111100000000000000000000000000000000010;
		10075: Delta = 46'sb0000000000011111111111111111111111111111111110;
		8534: Delta = 46'sb1111111111011111111111111111111111111111111110;
		1543: Delta = 46'sb0000000001000000000000000000000000000000000010;
		17074: Delta = 46'sb1111111111000000000000000000000000000000000010;
		1539: Delta = 46'sb0000000000111111111111111111111111111111111110;
		17070: Delta = 46'sb1111111110111111111111111111111111111111111110;
		3084: Delta = 46'sb0000000010000000000000000000000000000000000010;
		15533: Delta = 46'sb1111111110000000000000000000000000000000000010;
		3080: Delta = 46'sb0000000001111111111111111111111111111111111110;
		15529: Delta = 46'sb1111111101111111111111111111111111111111111110;
		6166: Delta = 46'sb0000000100000000000000000000000000000000000010;
		12451: Delta = 46'sb1111111100000000000000000000000000000000000010;
		6162: Delta = 46'sb0000000011111111111111111111111111111111111110;
		12447: Delta = 46'sb1111111011111111111111111111111111111111111110;
		12330: Delta = 46'sb0000001000000000000000000000000000000000000010;
		6287: Delta = 46'sb1111111000000000000000000000000000000000000010;
		12326: Delta = 46'sb0000000111111111111111111111111111111111111110;
		6283: Delta = 46'sb1111110111111111111111111111111111111111111110;
		6045: Delta = 46'sb0000010000000000000000000000000000000000000010;
		12572: Delta = 46'sb1111110000000000000000000000000000000000000010;
		6041: Delta = 46'sb0000001111111111111111111111111111111111111110;
		12568: Delta = 46'sb1111101111111111111111111111111111111111111110;
		12088: Delta = 46'sb0000100000000000000000000000000000000000000010;
		6529: Delta = 46'sb1111100000000000000000000000000000000000000010;
		12084: Delta = 46'sb0000011111111111111111111111111111111111111110;
		6525: Delta = 46'sb1111011111111111111111111111111111111111111110;
		5561: Delta = 46'sb0001000000000000000000000000000000000000000010;
		13056: Delta = 46'sb1111000000000000000000000000000000000000000010;
		5557: Delta = 46'sb0000111111111111111111111111111111111111111110;
		13052: Delta = 46'sb1110111111111111111111111111111111111111111110;
		11120: Delta = 46'sb0010000000000000000000000000000000000000000010;
		7497: Delta = 46'sb1110000000000000000000000000000000000000000010;
		11116: Delta = 46'sb0001111111111111111111111111111111111111111110;
		7493: Delta = 46'sb1101111111111111111111111111111111111111111110;
		3625: Delta = 46'sb0100000000000000000000000000000000000000000010;
		14992: Delta = 46'sb1100000000000000000000000000000000000000000010;
		3621: Delta = 46'sb0011111111111111111111111111111111111111111110;
		14988: Delta = 46'sb1011111111111111111111111111111111111111111110;
		12: Delta = 46'sb0000000000000000000000000000000000000000001100;
		18601: Delta = 46'sb1111111111111111111111111111111111111111110100;
		20: Delta = 46'sb0000000000000000000000000000000000000000010100;
		18593: Delta = 46'sb1111111111111111111111111111111111111111101100;
		36: Delta = 46'sb0000000000000000000000000000000000000000100100;
		18585: Delta = 46'sb1111111111111111111111111111111111111111100100;
		28: Delta = 46'sb0000000000000000000000000000000000000000011100;
		18577: Delta = 46'sb1111111111111111111111111111111111111111011100;
		68: Delta = 46'sb0000000000000000000000000000000000000001000100;
		18553: Delta = 46'sb1111111111111111111111111111111111111111000100;
		60: Delta = 46'sb0000000000000000000000000000000000000000111100;
		18545: Delta = 46'sb1111111111111111111111111111111111111110111100;
		132: Delta = 46'sb0000000000000000000000000000000000000010000100;
		18489: Delta = 46'sb1111111111111111111111111111111111111110000100;
		124: Delta = 46'sb0000000000000000000000000000000000000001111100;
		18481: Delta = 46'sb1111111111111111111111111111111111111101111100;
		260: Delta = 46'sb0000000000000000000000000000000000000100000100;
		18361: Delta = 46'sb1111111111111111111111111111111111111100000100;
		252: Delta = 46'sb0000000000000000000000000000000000000011111100;
		18353: Delta = 46'sb1111111111111111111111111111111111111011111100;
		516: Delta = 46'sb0000000000000000000000000000000000001000000100;
		18105: Delta = 46'sb1111111111111111111111111111111111111000000100;
		508: Delta = 46'sb0000000000000000000000000000000000000111111100;
		18097: Delta = 46'sb1111111111111111111111111111111111110111111100;
		1028: Delta = 46'sb0000000000000000000000000000000000010000000100;
		17593: Delta = 46'sb1111111111111111111111111111111111110000000100;
		1020: Delta = 46'sb0000000000000000000000000000000000001111111100;
		17585: Delta = 46'sb1111111111111111111111111111111111101111111100;
		2052: Delta = 46'sb0000000000000000000000000000000000100000000100;
		16569: Delta = 46'sb1111111111111111111111111111111111100000000100;
		2044: Delta = 46'sb0000000000000000000000000000000000011111111100;
		16561: Delta = 46'sb1111111111111111111111111111111111011111111100;
		4100: Delta = 46'sb0000000000000000000000000000000001000000000100;
		14521: Delta = 46'sb1111111111111111111111111111111111000000000100;
		4092: Delta = 46'sb0000000000000000000000000000000000111111111100;
		14513: Delta = 46'sb1111111111111111111111111111111110111111111100;
		8196: Delta = 46'sb0000000000000000000000000000000010000000000100;
		10425: Delta = 46'sb1111111111111111111111111111111110000000000100;
		8188: Delta = 46'sb0000000000000000000000000000000001111111111100;
		10417: Delta = 46'sb1111111111111111111111111111111101111111111100;
		16388: Delta = 46'sb0000000000000000000000000000000100000000000100;
		2233: Delta = 46'sb1111111111111111111111111111111100000000000100;
		16380: Delta = 46'sb0000000000000000000000000000000011111111111100;
		2225: Delta = 46'sb1111111111111111111111111111111011111111111100;
		14159: Delta = 46'sb0000000000000000000000000000001000000000000100;
		4462: Delta = 46'sb1111111111111111111111111111111000000000000100;
		14151: Delta = 46'sb0000000000000000000000000000000111111111111100;
		4454: Delta = 46'sb1111111111111111111111111111110111111111111100;
		9701: Delta = 46'sb0000000000000000000000000000010000000000000100;
		8920: Delta = 46'sb1111111111111111111111111111110000000000000100;
		9693: Delta = 46'sb0000000000000000000000000000001111111111111100;
		8912: Delta = 46'sb1111111111111111111111111111101111111111111100;
		785: Delta = 46'sb0000000000000000000000000000100000000000000100;
		17836: Delta = 46'sb1111111111111111111111111111100000000000000100;
		777: Delta = 46'sb0000000000000000000000000000011111111111111100;
		17828: Delta = 46'sb1111111111111111111111111111011111111111111100;
		1566: Delta = 46'sb0000000000000000000000000001000000000000000100;
		17055: Delta = 46'sb1111111111111111111111111111000000000000000100;
		1558: Delta = 46'sb0000000000000000000000000000111111111111111100;
		17047: Delta = 46'sb1111111111111111111111111110111111111111111100;
		3128: Delta = 46'sb0000000000000000000000000010000000000000000100;
		15493: Delta = 46'sb1111111111111111111111111110000000000000000100;
		3120: Delta = 46'sb0000000000000000000000000001111111111111111100;
		15485: Delta = 46'sb1111111111111111111111111101111111111111111100;
		6252: Delta = 46'sb0000000000000000000000000100000000000000000100;
		12369: Delta = 46'sb1111111111111111111111111100000000000000000100;
		6244: Delta = 46'sb0000000000000000000000000011111111111111111100;
		12361: Delta = 46'sb1111111111111111111111111011111111111111111100;
		12500: Delta = 46'sb0000000000000000000000001000000000000000000100;
		6121: Delta = 46'sb1111111111111111111111111000000000000000000100;
		12492: Delta = 46'sb0000000000000000000000000111111111111111111100;
		6113: Delta = 46'sb1111111111111111111111110111111111111111111100;
		6383: Delta = 46'sb0000000000000000000000010000000000000000000100;
		12238: Delta = 46'sb1111111111111111111111110000000000000000000100;
		6375: Delta = 46'sb0000000000000000000000001111111111111111111100;
		12230: Delta = 46'sb1111111111111111111111101111111111111111111100;
		12762: Delta = 46'sb0000000000000000000000100000000000000000000100;
		5859: Delta = 46'sb1111111111111111111111100000000000000000000100;
		12754: Delta = 46'sb0000000000000000000000011111111111111111111100;
		5851: Delta = 46'sb1111111111111111111111011111111111111111111100;
		6907: Delta = 46'sb0000000000000000000001000000000000000000000100;
		11714: Delta = 46'sb1111111111111111111111000000000000000000000100;
		6899: Delta = 46'sb0000000000000000000000111111111111111111111100;
		11706: Delta = 46'sb1111111111111111111110111111111111111111111100;
		13810: Delta = 46'sb0000000000000000000010000000000000000000000100;
		4811: Delta = 46'sb1111111111111111111110000000000000000000000100;
		13802: Delta = 46'sb0000000000000000000001111111111111111111111100;
		4803: Delta = 46'sb1111111111111111111101111111111111111111111100;
		9003: Delta = 46'sb0000000000000000000100000000000000000000000100;
		9618: Delta = 46'sb1111111111111111111100000000000000000000000100;
		8995: Delta = 46'sb0000000000000000000011111111111111111111111100;
		9610: Delta = 46'sb1111111111111111111011111111111111111111111100;
		18002: Delta = 46'sb0000000000000000001000000000000000000000000100;
		619: Delta = 46'sb1111111111111111111000000000000000000000000100;
		17994: Delta = 46'sb0000000000000000000111111111111111111111111100;
		611: Delta = 46'sb1111111111111111110111111111111111111111111100;
		17387: Delta = 46'sb0000000000000000010000000000000000000000000100;
		1234: Delta = 46'sb1111111111111111110000000000000000000000000100;
		17379: Delta = 46'sb0000000000000000001111111111111111111111111100;
		1226: Delta = 46'sb1111111111111111101111111111111111111111111100;
		16157: Delta = 46'sb0000000000000000100000000000000000000000000100;
		2464: Delta = 46'sb1111111111111111100000000000000000000000000100;
		16149: Delta = 46'sb0000000000000000011111111111111111111111111100;
		2456: Delta = 46'sb1111111111111111011111111111111111111111111100;
		13697: Delta = 46'sb0000000000000001000000000000000000000000000100;
		4924: Delta = 46'sb1111111111111111000000000000000000000000000100;
		13689: Delta = 46'sb0000000000000000111111111111111111111111111100;
		4916: Delta = 46'sb1111111111111110111111111111111111111111111100;
		8777: Delta = 46'sb0000000000000010000000000000000000000000000100;
		9844: Delta = 46'sb1111111111111110000000000000000000000000000100;
		8769: Delta = 46'sb0000000000000001111111111111111111111111111100;
		9836: Delta = 46'sb1111111111111101111111111111111111111111111100;
		17550: Delta = 46'sb0000000000000100000000000000000000000000000100;
		1071: Delta = 46'sb1111111111111100000000000000000000000000000100;
		17542: Delta = 46'sb0000000000000011111111111111111111111111111100;
		1063: Delta = 46'sb1111111111111011111111111111111111111111111100;
		16483: Delta = 46'sb0000000000001000000000000000000000000000000100;
		2138: Delta = 46'sb1111111111111000000000000000000000000000000100;
		16475: Delta = 46'sb0000000000000111111111111111111111111111111100;
		2130: Delta = 46'sb1111111111110111111111111111111111111111111100;
		14349: Delta = 46'sb0000000000010000000000000000000000000000000100;
		4272: Delta = 46'sb1111111111110000000000000000000000000000000100;
		14341: Delta = 46'sb0000000000001111111111111111111111111111111100;
		4264: Delta = 46'sb1111111111101111111111111111111111111111111100;
		10081: Delta = 46'sb0000000000100000000000000000000000000000000100;
		8540: Delta = 46'sb1111111111100000000000000000000000000000000100;
		10073: Delta = 46'sb0000000000011111111111111111111111111111111100;
		8532: Delta = 46'sb1111111111011111111111111111111111111111111100;
		1545: Delta = 46'sb0000000001000000000000000000000000000000000100;
		17076: Delta = 46'sb1111111111000000000000000000000000000000000100;
		1537: Delta = 46'sb0000000000111111111111111111111111111111111100;
		17068: Delta = 46'sb1111111110111111111111111111111111111111111100;
		3086: Delta = 46'sb0000000010000000000000000000000000000000000100;
		15535: Delta = 46'sb1111111110000000000000000000000000000000000100;
		3078: Delta = 46'sb0000000001111111111111111111111111111111111100;
		15527: Delta = 46'sb1111111101111111111111111111111111111111111100;
		6168: Delta = 46'sb0000000100000000000000000000000000000000000100;
		12453: Delta = 46'sb1111111100000000000000000000000000000000000100;
		6160: Delta = 46'sb0000000011111111111111111111111111111111111100;
		12445: Delta = 46'sb1111111011111111111111111111111111111111111100;
		12332: Delta = 46'sb0000001000000000000000000000000000000000000100;
		6289: Delta = 46'sb1111111000000000000000000000000000000000000100;
		12324: Delta = 46'sb0000000111111111111111111111111111111111111100;
		6281: Delta = 46'sb1111110111111111111111111111111111111111111100;
		6047: Delta = 46'sb0000010000000000000000000000000000000000000100;
		12574: Delta = 46'sb1111110000000000000000000000000000000000000100;
		6039: Delta = 46'sb0000001111111111111111111111111111111111111100;
		12566: Delta = 46'sb1111101111111111111111111111111111111111111100;
		12090: Delta = 46'sb0000100000000000000000000000000000000000000100;
		6531: Delta = 46'sb1111100000000000000000000000000000000000000100;
		12082: Delta = 46'sb0000011111111111111111111111111111111111111100;
		6523: Delta = 46'sb1111011111111111111111111111111111111111111100;
		5563: Delta = 46'sb0001000000000000000000000000000000000000000100;
		13058: Delta = 46'sb1111000000000000000000000000000000000000000100;
		5555: Delta = 46'sb0000111111111111111111111111111111111111111100;
		13050: Delta = 46'sb1110111111111111111111111111111111111111111100;
		11122: Delta = 46'sb0010000000000000000000000000000000000000000100;
		7499: Delta = 46'sb1110000000000000000000000000000000000000000100;
		11114: Delta = 46'sb0001111111111111111111111111111111111111111100;
		7491: Delta = 46'sb1101111111111111111111111111111111111111111100;
		3627: Delta = 46'sb0100000000000000000000000000000000000000000100;
		14994: Delta = 46'sb1100000000000000000000000000000000000000000100;
		3619: Delta = 46'sb0011111111111111111111111111111111111111111100;
		14986: Delta = 46'sb1011111111111111111111111111111111111111111100;
		24: Delta = 46'sb0000000000000000000000000000000000000000011000;
		18589: Delta = 46'sb1111111111111111111111111111111111111111101000;
		40: Delta = 46'sb0000000000000000000000000000000000000000101000;
		18573: Delta = 46'sb1111111111111111111111111111111111111111011000;
		72: Delta = 46'sb0000000000000000000000000000000000000001001000;
		18557: Delta = 46'sb1111111111111111111111111111111111111111001000;
		56: Delta = 46'sb0000000000000000000000000000000000000000111000;
		18541: Delta = 46'sb1111111111111111111111111111111111111110111000;
		136: Delta = 46'sb0000000000000000000000000000000000000010001000;
		18493: Delta = 46'sb1111111111111111111111111111111111111110001000;
		120: Delta = 46'sb0000000000000000000000000000000000000001111000;
		18477: Delta = 46'sb1111111111111111111111111111111111111101111000;
		264: Delta = 46'sb0000000000000000000000000000000000000100001000;
		18365: Delta = 46'sb1111111111111111111111111111111111111100001000;
		248: Delta = 46'sb0000000000000000000000000000000000000011111000;
		18349: Delta = 46'sb1111111111111111111111111111111111111011111000;
		520: Delta = 46'sb0000000000000000000000000000000000001000001000;
		18109: Delta = 46'sb1111111111111111111111111111111111111000001000;
		504: Delta = 46'sb0000000000000000000000000000000000000111111000;
		18093: Delta = 46'sb1111111111111111111111111111111111110111111000;
		1032: Delta = 46'sb0000000000000000000000000000000000010000001000;
		17597: Delta = 46'sb1111111111111111111111111111111111110000001000;
		1016: Delta = 46'sb0000000000000000000000000000000000001111111000;
		17581: Delta = 46'sb1111111111111111111111111111111111101111111000;
		2056: Delta = 46'sb0000000000000000000000000000000000100000001000;
		16573: Delta = 46'sb1111111111111111111111111111111111100000001000;
		2040: Delta = 46'sb0000000000000000000000000000000000011111111000;
		16557: Delta = 46'sb1111111111111111111111111111111111011111111000;
		4104: Delta = 46'sb0000000000000000000000000000000001000000001000;
		14525: Delta = 46'sb1111111111111111111111111111111111000000001000;
		4088: Delta = 46'sb0000000000000000000000000000000000111111111000;
		14509: Delta = 46'sb1111111111111111111111111111111110111111111000;
		8200: Delta = 46'sb0000000000000000000000000000000010000000001000;
		10429: Delta = 46'sb1111111111111111111111111111111110000000001000;
		8184: Delta = 46'sb0000000000000000000000000000000001111111111000;
		10413: Delta = 46'sb1111111111111111111111111111111101111111111000;
		16392: Delta = 46'sb0000000000000000000000000000000100000000001000;
		2237: Delta = 46'sb1111111111111111111111111111111100000000001000;
		16376: Delta = 46'sb0000000000000000000000000000000011111111111000;
		2221: Delta = 46'sb1111111111111111111111111111111011111111111000;
		14163: Delta = 46'sb0000000000000000000000000000001000000000001000;
		4466: Delta = 46'sb1111111111111111111111111111111000000000001000;
		14147: Delta = 46'sb0000000000000000000000000000000111111111111000;
		4450: Delta = 46'sb1111111111111111111111111111110111111111111000;
		9705: Delta = 46'sb0000000000000000000000000000010000000000001000;
		8924: Delta = 46'sb1111111111111111111111111111110000000000001000;
		9689: Delta = 46'sb0000000000000000000000000000001111111111111000;
		8908: Delta = 46'sb1111111111111111111111111111101111111111111000;
		789: Delta = 46'sb0000000000000000000000000000100000000000001000;
		17840: Delta = 46'sb1111111111111111111111111111100000000000001000;
		773: Delta = 46'sb0000000000000000000000000000011111111111111000;
		17824: Delta = 46'sb1111111111111111111111111111011111111111111000;
		1570: Delta = 46'sb0000000000000000000000000001000000000000001000;
		17059: Delta = 46'sb1111111111111111111111111111000000000000001000;
		1554: Delta = 46'sb0000000000000000000000000000111111111111111000;
		17043: Delta = 46'sb1111111111111111111111111110111111111111111000;
		3132: Delta = 46'sb0000000000000000000000000010000000000000001000;
		15497: Delta = 46'sb1111111111111111111111111110000000000000001000;
		3116: Delta = 46'sb0000000000000000000000000001111111111111111000;
		15481: Delta = 46'sb1111111111111111111111111101111111111111111000;
		6256: Delta = 46'sb0000000000000000000000000100000000000000001000;
		12373: Delta = 46'sb1111111111111111111111111100000000000000001000;
		6240: Delta = 46'sb0000000000000000000000000011111111111111111000;
		12357: Delta = 46'sb1111111111111111111111111011111111111111111000;
		12504: Delta = 46'sb0000000000000000000000001000000000000000001000;
		6125: Delta = 46'sb1111111111111111111111111000000000000000001000;
		12488: Delta = 46'sb0000000000000000000000000111111111111111111000;
		6109: Delta = 46'sb1111111111111111111111110111111111111111111000;
		6387: Delta = 46'sb0000000000000000000000010000000000000000001000;
		12242: Delta = 46'sb1111111111111111111111110000000000000000001000;
		6371: Delta = 46'sb0000000000000000000000001111111111111111111000;
		12226: Delta = 46'sb1111111111111111111111101111111111111111111000;
		12766: Delta = 46'sb0000000000000000000000100000000000000000001000;
		5863: Delta = 46'sb1111111111111111111111100000000000000000001000;
		12750: Delta = 46'sb0000000000000000000000011111111111111111111000;
		5847: Delta = 46'sb1111111111111111111111011111111111111111111000;
		6911: Delta = 46'sb0000000000000000000001000000000000000000001000;
		11718: Delta = 46'sb1111111111111111111111000000000000000000001000;
		6895: Delta = 46'sb0000000000000000000000111111111111111111111000;
		11702: Delta = 46'sb1111111111111111111110111111111111111111111000;
		13814: Delta = 46'sb0000000000000000000010000000000000000000001000;
		4815: Delta = 46'sb1111111111111111111110000000000000000000001000;
		13798: Delta = 46'sb0000000000000000000001111111111111111111111000;
		4799: Delta = 46'sb1111111111111111111101111111111111111111111000;
		9007: Delta = 46'sb0000000000000000000100000000000000000000001000;
		9622: Delta = 46'sb1111111111111111111100000000000000000000001000;
		8991: Delta = 46'sb0000000000000000000011111111111111111111111000;
		9606: Delta = 46'sb1111111111111111111011111111111111111111111000;
		18006: Delta = 46'sb0000000000000000001000000000000000000000001000;
		623: Delta = 46'sb1111111111111111111000000000000000000000001000;
		17990: Delta = 46'sb0000000000000000000111111111111111111111111000;
		607: Delta = 46'sb1111111111111111110111111111111111111111111000;
		17391: Delta = 46'sb0000000000000000010000000000000000000000001000;
		1238: Delta = 46'sb1111111111111111110000000000000000000000001000;
		17375: Delta = 46'sb0000000000000000001111111111111111111111111000;
		1222: Delta = 46'sb1111111111111111101111111111111111111111111000;
		16161: Delta = 46'sb0000000000000000100000000000000000000000001000;
		2468: Delta = 46'sb1111111111111111100000000000000000000000001000;
		16145: Delta = 46'sb0000000000000000011111111111111111111111111000;
		2452: Delta = 46'sb1111111111111111011111111111111111111111111000;
		13701: Delta = 46'sb0000000000000001000000000000000000000000001000;
		4928: Delta = 46'sb1111111111111111000000000000000000000000001000;
		13685: Delta = 46'sb0000000000000000111111111111111111111111111000;
		4912: Delta = 46'sb1111111111111110111111111111111111111111111000;
		8781: Delta = 46'sb0000000000000010000000000000000000000000001000;
		9848: Delta = 46'sb1111111111111110000000000000000000000000001000;
		8765: Delta = 46'sb0000000000000001111111111111111111111111111000;
		9832: Delta = 46'sb1111111111111101111111111111111111111111111000;
		17554: Delta = 46'sb0000000000000100000000000000000000000000001000;
		1075: Delta = 46'sb1111111111111100000000000000000000000000001000;
		17538: Delta = 46'sb0000000000000011111111111111111111111111111000;
		1059: Delta = 46'sb1111111111111011111111111111111111111111111000;
		16487: Delta = 46'sb0000000000001000000000000000000000000000001000;
		2142: Delta = 46'sb1111111111111000000000000000000000000000001000;
		16471: Delta = 46'sb0000000000000111111111111111111111111111111000;
		2126: Delta = 46'sb1111111111110111111111111111111111111111111000;
		14353: Delta = 46'sb0000000000010000000000000000000000000000001000;
		4276: Delta = 46'sb1111111111110000000000000000000000000000001000;
		14337: Delta = 46'sb0000000000001111111111111111111111111111111000;
		4260: Delta = 46'sb1111111111101111111111111111111111111111111000;
		10085: Delta = 46'sb0000000000100000000000000000000000000000001000;
		8544: Delta = 46'sb1111111111100000000000000000000000000000001000;
		10069: Delta = 46'sb0000000000011111111111111111111111111111111000;
		8528: Delta = 46'sb1111111111011111111111111111111111111111111000;
		1549: Delta = 46'sb0000000001000000000000000000000000000000001000;
		17080: Delta = 46'sb1111111111000000000000000000000000000000001000;
		1533: Delta = 46'sb0000000000111111111111111111111111111111111000;
		17064: Delta = 46'sb1111111110111111111111111111111111111111111000;
		3090: Delta = 46'sb0000000010000000000000000000000000000000001000;
		15539: Delta = 46'sb1111111110000000000000000000000000000000001000;
		3074: Delta = 46'sb0000000001111111111111111111111111111111111000;
		15523: Delta = 46'sb1111111101111111111111111111111111111111111000;
		6172: Delta = 46'sb0000000100000000000000000000000000000000001000;
		12457: Delta = 46'sb1111111100000000000000000000000000000000001000;
		6156: Delta = 46'sb0000000011111111111111111111111111111111111000;
		12441: Delta = 46'sb1111111011111111111111111111111111111111111000;
		12336: Delta = 46'sb0000001000000000000000000000000000000000001000;
		6293: Delta = 46'sb1111111000000000000000000000000000000000001000;
		12320: Delta = 46'sb0000000111111111111111111111111111111111111000;
		6277: Delta = 46'sb1111110111111111111111111111111111111111111000;
		6051: Delta = 46'sb0000010000000000000000000000000000000000001000;
		12578: Delta = 46'sb1111110000000000000000000000000000000000001000;
		6035: Delta = 46'sb0000001111111111111111111111111111111111111000;
		12562: Delta = 46'sb1111101111111111111111111111111111111111111000;
		12094: Delta = 46'sb0000100000000000000000000000000000000000001000;
		6535: Delta = 46'sb1111100000000000000000000000000000000000001000;
		12078: Delta = 46'sb0000011111111111111111111111111111111111111000;
		6519: Delta = 46'sb1111011111111111111111111111111111111111111000;
		5567: Delta = 46'sb0001000000000000000000000000000000000000001000;
		13062: Delta = 46'sb1111000000000000000000000000000000000000001000;
		5551: Delta = 46'sb0000111111111111111111111111111111111111111000;
		13046: Delta = 46'sb1110111111111111111111111111111111111111111000;
		11126: Delta = 46'sb0010000000000000000000000000000000000000001000;
		7503: Delta = 46'sb1110000000000000000000000000000000000000001000;
		11110: Delta = 46'sb0001111111111111111111111111111111111111111000;
		7487: Delta = 46'sb1101111111111111111111111111111111111111111000;
		3631: Delta = 46'sb0100000000000000000000000000000000000000001000;
		14998: Delta = 46'sb1100000000000000000000000000000000000000001000;
		3615: Delta = 46'sb0011111111111111111111111111111111111111111000;
		14982: Delta = 46'sb1011111111111111111111111111111111111111111000;
		48: Delta = 46'sb0000000000000000000000000000000000000000110000;
		18565: Delta = 46'sb1111111111111111111111111111111111111111010000;
		80: Delta = 46'sb0000000000000000000000000000000000000001010000;
		18533: Delta = 46'sb1111111111111111111111111111111111111110110000;
		144: Delta = 46'sb0000000000000000000000000000000000000010010000;
		18501: Delta = 46'sb1111111111111111111111111111111111111110010000;
		112: Delta = 46'sb0000000000000000000000000000000000000001110000;
		18469: Delta = 46'sb1111111111111111111111111111111111111101110000;
		272: Delta = 46'sb0000000000000000000000000000000000000100010000;
		18373: Delta = 46'sb1111111111111111111111111111111111111100010000;
		240: Delta = 46'sb0000000000000000000000000000000000000011110000;
		18341: Delta = 46'sb1111111111111111111111111111111111111011110000;
		528: Delta = 46'sb0000000000000000000000000000000000001000010000;
		18117: Delta = 46'sb1111111111111111111111111111111111111000010000;
		496: Delta = 46'sb0000000000000000000000000000000000000111110000;
		18085: Delta = 46'sb1111111111111111111111111111111111110111110000;
		1040: Delta = 46'sb0000000000000000000000000000000000010000010000;
		17605: Delta = 46'sb1111111111111111111111111111111111110000010000;
		1008: Delta = 46'sb0000000000000000000000000000000000001111110000;
		17573: Delta = 46'sb1111111111111111111111111111111111101111110000;
		2064: Delta = 46'sb0000000000000000000000000000000000100000010000;
		16581: Delta = 46'sb1111111111111111111111111111111111100000010000;
		2032: Delta = 46'sb0000000000000000000000000000000000011111110000;
		16549: Delta = 46'sb1111111111111111111111111111111111011111110000;
		4112: Delta = 46'sb0000000000000000000000000000000001000000010000;
		14533: Delta = 46'sb1111111111111111111111111111111111000000010000;
		4080: Delta = 46'sb0000000000000000000000000000000000111111110000;
		14501: Delta = 46'sb1111111111111111111111111111111110111111110000;
		8208: Delta = 46'sb0000000000000000000000000000000010000000010000;
		10437: Delta = 46'sb1111111111111111111111111111111110000000010000;
		8176: Delta = 46'sb0000000000000000000000000000000001111111110000;
		10405: Delta = 46'sb1111111111111111111111111111111101111111110000;
		16400: Delta = 46'sb0000000000000000000000000000000100000000010000;
		2245: Delta = 46'sb1111111111111111111111111111111100000000010000;
		16368: Delta = 46'sb0000000000000000000000000000000011111111110000;
		2213: Delta = 46'sb1111111111111111111111111111111011111111110000;
		14171: Delta = 46'sb0000000000000000000000000000001000000000010000;
		4474: Delta = 46'sb1111111111111111111111111111111000000000010000;
		14139: Delta = 46'sb0000000000000000000000000000000111111111110000;
		4442: Delta = 46'sb1111111111111111111111111111110111111111110000;
		9713: Delta = 46'sb0000000000000000000000000000010000000000010000;
		8932: Delta = 46'sb1111111111111111111111111111110000000000010000;
		9681: Delta = 46'sb0000000000000000000000000000001111111111110000;
		8900: Delta = 46'sb1111111111111111111111111111101111111111110000;
		797: Delta = 46'sb0000000000000000000000000000100000000000010000;
		17848: Delta = 46'sb1111111111111111111111111111100000000000010000;
		765: Delta = 46'sb0000000000000000000000000000011111111111110000;
		17816: Delta = 46'sb1111111111111111111111111111011111111111110000;
		1578: Delta = 46'sb0000000000000000000000000001000000000000010000;
		17067: Delta = 46'sb1111111111111111111111111111000000000000010000;
		1546: Delta = 46'sb0000000000000000000000000000111111111111110000;
		17035: Delta = 46'sb1111111111111111111111111110111111111111110000;
		3140: Delta = 46'sb0000000000000000000000000010000000000000010000;
		15505: Delta = 46'sb1111111111111111111111111110000000000000010000;
		3108: Delta = 46'sb0000000000000000000000000001111111111111110000;
		15473: Delta = 46'sb1111111111111111111111111101111111111111110000;
		6264: Delta = 46'sb0000000000000000000000000100000000000000010000;
		12381: Delta = 46'sb1111111111111111111111111100000000000000010000;
		6232: Delta = 46'sb0000000000000000000000000011111111111111110000;
		12349: Delta = 46'sb1111111111111111111111111011111111111111110000;
		12512: Delta = 46'sb0000000000000000000000001000000000000000010000;
		6133: Delta = 46'sb1111111111111111111111111000000000000000010000;
		12480: Delta = 46'sb0000000000000000000000000111111111111111110000;
		6101: Delta = 46'sb1111111111111111111111110111111111111111110000;
		6395: Delta = 46'sb0000000000000000000000010000000000000000010000;
		12250: Delta = 46'sb1111111111111111111111110000000000000000010000;
		6363: Delta = 46'sb0000000000000000000000001111111111111111110000;
		12218: Delta = 46'sb1111111111111111111111101111111111111111110000;
		12774: Delta = 46'sb0000000000000000000000100000000000000000010000;
		5871: Delta = 46'sb1111111111111111111111100000000000000000010000;
		12742: Delta = 46'sb0000000000000000000000011111111111111111110000;
		5839: Delta = 46'sb1111111111111111111111011111111111111111110000;
		6919: Delta = 46'sb0000000000000000000001000000000000000000010000;
		11726: Delta = 46'sb1111111111111111111111000000000000000000010000;
		6887: Delta = 46'sb0000000000000000000000111111111111111111110000;
		11694: Delta = 46'sb1111111111111111111110111111111111111111110000;
		13822: Delta = 46'sb0000000000000000000010000000000000000000010000;
		4823: Delta = 46'sb1111111111111111111110000000000000000000010000;
		13790: Delta = 46'sb0000000000000000000001111111111111111111110000;
		4791: Delta = 46'sb1111111111111111111101111111111111111111110000;
		9015: Delta = 46'sb0000000000000000000100000000000000000000010000;
		9630: Delta = 46'sb1111111111111111111100000000000000000000010000;
		8983: Delta = 46'sb0000000000000000000011111111111111111111110000;
		9598: Delta = 46'sb1111111111111111111011111111111111111111110000;
		18014: Delta = 46'sb0000000000000000001000000000000000000000010000;
		631: Delta = 46'sb1111111111111111111000000000000000000000010000;
		17982: Delta = 46'sb0000000000000000000111111111111111111111110000;
		599: Delta = 46'sb1111111111111111110111111111111111111111110000;
		17399: Delta = 46'sb0000000000000000010000000000000000000000010000;
		1246: Delta = 46'sb1111111111111111110000000000000000000000010000;
		17367: Delta = 46'sb0000000000000000001111111111111111111111110000;
		1214: Delta = 46'sb1111111111111111101111111111111111111111110000;
		16169: Delta = 46'sb0000000000000000100000000000000000000000010000;
		2476: Delta = 46'sb1111111111111111100000000000000000000000010000;
		16137: Delta = 46'sb0000000000000000011111111111111111111111110000;
		2444: Delta = 46'sb1111111111111111011111111111111111111111110000;
		13709: Delta = 46'sb0000000000000001000000000000000000000000010000;
		4936: Delta = 46'sb1111111111111111000000000000000000000000010000;
		13677: Delta = 46'sb0000000000000000111111111111111111111111110000;
		4904: Delta = 46'sb1111111111111110111111111111111111111111110000;
		8789: Delta = 46'sb0000000000000010000000000000000000000000010000;
		9856: Delta = 46'sb1111111111111110000000000000000000000000010000;
		8757: Delta = 46'sb0000000000000001111111111111111111111111110000;
		9824: Delta = 46'sb1111111111111101111111111111111111111111110000;
		17562: Delta = 46'sb0000000000000100000000000000000000000000010000;
		1083: Delta = 46'sb1111111111111100000000000000000000000000010000;
		17530: Delta = 46'sb0000000000000011111111111111111111111111110000;
		1051: Delta = 46'sb1111111111111011111111111111111111111111110000;
		16495: Delta = 46'sb0000000000001000000000000000000000000000010000;
		2150: Delta = 46'sb1111111111111000000000000000000000000000010000;
		16463: Delta = 46'sb0000000000000111111111111111111111111111110000;
		2118: Delta = 46'sb1111111111110111111111111111111111111111110000;
		14361: Delta = 46'sb0000000000010000000000000000000000000000010000;
		4284: Delta = 46'sb1111111111110000000000000000000000000000010000;
		14329: Delta = 46'sb0000000000001111111111111111111111111111110000;
		4252: Delta = 46'sb1111111111101111111111111111111111111111110000;
		10093: Delta = 46'sb0000000000100000000000000000000000000000010000;
		8552: Delta = 46'sb1111111111100000000000000000000000000000010000;
		10061: Delta = 46'sb0000000000011111111111111111111111111111110000;
		8520: Delta = 46'sb1111111111011111111111111111111111111111110000;
		1557: Delta = 46'sb0000000001000000000000000000000000000000010000;
		17088: Delta = 46'sb1111111111000000000000000000000000000000010000;
		1525: Delta = 46'sb0000000000111111111111111111111111111111110000;
		17056: Delta = 46'sb1111111110111111111111111111111111111111110000;
		3098: Delta = 46'sb0000000010000000000000000000000000000000010000;
		15547: Delta = 46'sb1111111110000000000000000000000000000000010000;
		3066: Delta = 46'sb0000000001111111111111111111111111111111110000;
		15515: Delta = 46'sb1111111101111111111111111111111111111111110000;
		6180: Delta = 46'sb0000000100000000000000000000000000000000010000;
		12465: Delta = 46'sb1111111100000000000000000000000000000000010000;
		6148: Delta = 46'sb0000000011111111111111111111111111111111110000;
		12433: Delta = 46'sb1111111011111111111111111111111111111111110000;
		12344: Delta = 46'sb0000001000000000000000000000000000000000010000;
		6301: Delta = 46'sb1111111000000000000000000000000000000000010000;
		12312: Delta = 46'sb0000000111111111111111111111111111111111110000;
		6269: Delta = 46'sb1111110111111111111111111111111111111111110000;
		6059: Delta = 46'sb0000010000000000000000000000000000000000010000;
		12586: Delta = 46'sb1111110000000000000000000000000000000000010000;
		6027: Delta = 46'sb0000001111111111111111111111111111111111110000;
		12554: Delta = 46'sb1111101111111111111111111111111111111111110000;
		12102: Delta = 46'sb0000100000000000000000000000000000000000010000;
		6543: Delta = 46'sb1111100000000000000000000000000000000000010000;
		12070: Delta = 46'sb0000011111111111111111111111111111111111110000;
		6511: Delta = 46'sb1111011111111111111111111111111111111111110000;
		5575: Delta = 46'sb0001000000000000000000000000000000000000010000;
		13070: Delta = 46'sb1111000000000000000000000000000000000000010000;
		5543: Delta = 46'sb0000111111111111111111111111111111111111110000;
		13038: Delta = 46'sb1110111111111111111111111111111111111111110000;
		11134: Delta = 46'sb0010000000000000000000000000000000000000010000;
		7511: Delta = 46'sb1110000000000000000000000000000000000000010000;
		11102: Delta = 46'sb0001111111111111111111111111111111111111110000;
		7479: Delta = 46'sb1101111111111111111111111111111111111111110000;
		3639: Delta = 46'sb0100000000000000000000000000000000000000010000;
		15006: Delta = 46'sb1100000000000000000000000000000000000000010000;
		3607: Delta = 46'sb0011111111111111111111111111111111111111110000;
		14974: Delta = 46'sb1011111111111111111111111111111111111111110000;
		96: Delta = 46'sb0000000000000000000000000000000000000001100000;
		18517: Delta = 46'sb1111111111111111111111111111111111111110100000;
		160: Delta = 46'sb0000000000000000000000000000000000000010100000;
		18453: Delta = 46'sb1111111111111111111111111111111111111101100000;
		288: Delta = 46'sb0000000000000000000000000000000000000100100000;
		18389: Delta = 46'sb1111111111111111111111111111111111111100100000;
		224: Delta = 46'sb0000000000000000000000000000000000000011100000;
		18325: Delta = 46'sb1111111111111111111111111111111111111011100000;
		544: Delta = 46'sb0000000000000000000000000000000000001000100000;
		18133: Delta = 46'sb1111111111111111111111111111111111111000100000;
		480: Delta = 46'sb0000000000000000000000000000000000000111100000;
		18069: Delta = 46'sb1111111111111111111111111111111111110111100000;
		1056: Delta = 46'sb0000000000000000000000000000000000010000100000;
		17621: Delta = 46'sb1111111111111111111111111111111111110000100000;
		992: Delta = 46'sb0000000000000000000000000000000000001111100000;
		17557: Delta = 46'sb1111111111111111111111111111111111101111100000;
		2080: Delta = 46'sb0000000000000000000000000000000000100000100000;
		16597: Delta = 46'sb1111111111111111111111111111111111100000100000;
		2016: Delta = 46'sb0000000000000000000000000000000000011111100000;
		16533: Delta = 46'sb1111111111111111111111111111111111011111100000;
		4128: Delta = 46'sb0000000000000000000000000000000001000000100000;
		14549: Delta = 46'sb1111111111111111111111111111111111000000100000;
		4064: Delta = 46'sb0000000000000000000000000000000000111111100000;
		14485: Delta = 46'sb1111111111111111111111111111111110111111100000;
		8224: Delta = 46'sb0000000000000000000000000000000010000000100000;
		10453: Delta = 46'sb1111111111111111111111111111111110000000100000;
		8160: Delta = 46'sb0000000000000000000000000000000001111111100000;
		10389: Delta = 46'sb1111111111111111111111111111111101111111100000;
		16416: Delta = 46'sb0000000000000000000000000000000100000000100000;
		2261: Delta = 46'sb1111111111111111111111111111111100000000100000;
		16352: Delta = 46'sb0000000000000000000000000000000011111111100000;
		2197: Delta = 46'sb1111111111111111111111111111111011111111100000;
		14187: Delta = 46'sb0000000000000000000000000000001000000000100000;
		4490: Delta = 46'sb1111111111111111111111111111111000000000100000;
		14123: Delta = 46'sb0000000000000000000000000000000111111111100000;
		4426: Delta = 46'sb1111111111111111111111111111110111111111100000;
		9729: Delta = 46'sb0000000000000000000000000000010000000000100000;
		8948: Delta = 46'sb1111111111111111111111111111110000000000100000;
		9665: Delta = 46'sb0000000000000000000000000000001111111111100000;
		8884: Delta = 46'sb1111111111111111111111111111101111111111100000;
		813: Delta = 46'sb0000000000000000000000000000100000000000100000;
		17864: Delta = 46'sb1111111111111111111111111111100000000000100000;
		749: Delta = 46'sb0000000000000000000000000000011111111111100000;
		17800: Delta = 46'sb1111111111111111111111111111011111111111100000;
		1594: Delta = 46'sb0000000000000000000000000001000000000000100000;
		17083: Delta = 46'sb1111111111111111111111111111000000000000100000;
		1530: Delta = 46'sb0000000000000000000000000000111111111111100000;
		17019: Delta = 46'sb1111111111111111111111111110111111111111100000;
		3156: Delta = 46'sb0000000000000000000000000010000000000000100000;
		15521: Delta = 46'sb1111111111111111111111111110000000000000100000;
		3092: Delta = 46'sb0000000000000000000000000001111111111111100000;
		15457: Delta = 46'sb1111111111111111111111111101111111111111100000;
		6280: Delta = 46'sb0000000000000000000000000100000000000000100000;
		12397: Delta = 46'sb1111111111111111111111111100000000000000100000;
		6216: Delta = 46'sb0000000000000000000000000011111111111111100000;
		12333: Delta = 46'sb1111111111111111111111111011111111111111100000;
		12528: Delta = 46'sb0000000000000000000000001000000000000000100000;
		6149: Delta = 46'sb1111111111111111111111111000000000000000100000;
		12464: Delta = 46'sb0000000000000000000000000111111111111111100000;
		6085: Delta = 46'sb1111111111111111111111110111111111111111100000;
		6411: Delta = 46'sb0000000000000000000000010000000000000000100000;
		12266: Delta = 46'sb1111111111111111111111110000000000000000100000;
		6347: Delta = 46'sb0000000000000000000000001111111111111111100000;
		12202: Delta = 46'sb1111111111111111111111101111111111111111100000;
		12790: Delta = 46'sb0000000000000000000000100000000000000000100000;
		5887: Delta = 46'sb1111111111111111111111100000000000000000100000;
		12726: Delta = 46'sb0000000000000000000000011111111111111111100000;
		5823: Delta = 46'sb1111111111111111111111011111111111111111100000;
		6935: Delta = 46'sb0000000000000000000001000000000000000000100000;
		11742: Delta = 46'sb1111111111111111111111000000000000000000100000;
		6871: Delta = 46'sb0000000000000000000000111111111111111111100000;
		11678: Delta = 46'sb1111111111111111111110111111111111111111100000;
		13838: Delta = 46'sb0000000000000000000010000000000000000000100000;
		4839: Delta = 46'sb1111111111111111111110000000000000000000100000;
		13774: Delta = 46'sb0000000000000000000001111111111111111111100000;
		4775: Delta = 46'sb1111111111111111111101111111111111111111100000;
		9031: Delta = 46'sb0000000000000000000100000000000000000000100000;
		9646: Delta = 46'sb1111111111111111111100000000000000000000100000;
		8967: Delta = 46'sb0000000000000000000011111111111111111111100000;
		9582: Delta = 46'sb1111111111111111111011111111111111111111100000;
		18030: Delta = 46'sb0000000000000000001000000000000000000000100000;
		647: Delta = 46'sb1111111111111111111000000000000000000000100000;
		17966: Delta = 46'sb0000000000000000000111111111111111111111100000;
		583: Delta = 46'sb1111111111111111110111111111111111111111100000;
		17415: Delta = 46'sb0000000000000000010000000000000000000000100000;
		1262: Delta = 46'sb1111111111111111110000000000000000000000100000;
		17351: Delta = 46'sb0000000000000000001111111111111111111111100000;
		1198: Delta = 46'sb1111111111111111101111111111111111111111100000;
		16185: Delta = 46'sb0000000000000000100000000000000000000000100000;
		2492: Delta = 46'sb1111111111111111100000000000000000000000100000;
		16121: Delta = 46'sb0000000000000000011111111111111111111111100000;
		2428: Delta = 46'sb1111111111111111011111111111111111111111100000;
		13725: Delta = 46'sb0000000000000001000000000000000000000000100000;
		4952: Delta = 46'sb1111111111111111000000000000000000000000100000;
		13661: Delta = 46'sb0000000000000000111111111111111111111111100000;
		4888: Delta = 46'sb1111111111111110111111111111111111111111100000;
		8805: Delta = 46'sb0000000000000010000000000000000000000000100000;
		9872: Delta = 46'sb1111111111111110000000000000000000000000100000;
		8741: Delta = 46'sb0000000000000001111111111111111111111111100000;
		9808: Delta = 46'sb1111111111111101111111111111111111111111100000;
		17578: Delta = 46'sb0000000000000100000000000000000000000000100000;
		1099: Delta = 46'sb1111111111111100000000000000000000000000100000;
		17514: Delta = 46'sb0000000000000011111111111111111111111111100000;
		1035: Delta = 46'sb1111111111111011111111111111111111111111100000;
		16511: Delta = 46'sb0000000000001000000000000000000000000000100000;
		2166: Delta = 46'sb1111111111111000000000000000000000000000100000;
		16447: Delta = 46'sb0000000000000111111111111111111111111111100000;
		2102: Delta = 46'sb1111111111110111111111111111111111111111100000;
		14377: Delta = 46'sb0000000000010000000000000000000000000000100000;
		4300: Delta = 46'sb1111111111110000000000000000000000000000100000;
		14313: Delta = 46'sb0000000000001111111111111111111111111111100000;
		4236: Delta = 46'sb1111111111101111111111111111111111111111100000;
		10109: Delta = 46'sb0000000000100000000000000000000000000000100000;
		8568: Delta = 46'sb1111111111100000000000000000000000000000100000;
		10045: Delta = 46'sb0000000000011111111111111111111111111111100000;
		8504: Delta = 46'sb1111111111011111111111111111111111111111100000;
		1573: Delta = 46'sb0000000001000000000000000000000000000000100000;
		17104: Delta = 46'sb1111111111000000000000000000000000000000100000;
		1509: Delta = 46'sb0000000000111111111111111111111111111111100000;
		17040: Delta = 46'sb1111111110111111111111111111111111111111100000;
		3114: Delta = 46'sb0000000010000000000000000000000000000000100000;
		15563: Delta = 46'sb1111111110000000000000000000000000000000100000;
		3050: Delta = 46'sb0000000001111111111111111111111111111111100000;
		15499: Delta = 46'sb1111111101111111111111111111111111111111100000;
		6196: Delta = 46'sb0000000100000000000000000000000000000000100000;
		12481: Delta = 46'sb1111111100000000000000000000000000000000100000;
		6132: Delta = 46'sb0000000011111111111111111111111111111111100000;
		12417: Delta = 46'sb1111111011111111111111111111111111111111100000;
		12360: Delta = 46'sb0000001000000000000000000000000000000000100000;
		6317: Delta = 46'sb1111111000000000000000000000000000000000100000;
		12296: Delta = 46'sb0000000111111111111111111111111111111111100000;
		6253: Delta = 46'sb1111110111111111111111111111111111111111100000;
		6075: Delta = 46'sb0000010000000000000000000000000000000000100000;
		12602: Delta = 46'sb1111110000000000000000000000000000000000100000;
		6011: Delta = 46'sb0000001111111111111111111111111111111111100000;
		12538: Delta = 46'sb1111101111111111111111111111111111111111100000;
		12118: Delta = 46'sb0000100000000000000000000000000000000000100000;
		6559: Delta = 46'sb1111100000000000000000000000000000000000100000;
		12054: Delta = 46'sb0000011111111111111111111111111111111111100000;
		6495: Delta = 46'sb1111011111111111111111111111111111111111100000;
		5591: Delta = 46'sb0001000000000000000000000000000000000000100000;
		13086: Delta = 46'sb1111000000000000000000000000000000000000100000;
		5527: Delta = 46'sb0000111111111111111111111111111111111111100000;
		13022: Delta = 46'sb1110111111111111111111111111111111111111100000;
		11150: Delta = 46'sb0010000000000000000000000000000000000000100000;
		7527: Delta = 46'sb1110000000000000000000000000000000000000100000;
		11086: Delta = 46'sb0001111111111111111111111111111111111111100000;
		7463: Delta = 46'sb1101111111111111111111111111111111111111100000;
		3655: Delta = 46'sb0100000000000000000000000000000000000000100000;
		15022: Delta = 46'sb1100000000000000000000000000000000000000100000;
		3591: Delta = 46'sb0011111111111111111111111111111111111111100000;
		14958: Delta = 46'sb1011111111111111111111111111111111111111100000;
		192: Delta = 46'sb0000000000000000000000000000000000000011000000;
		18421: Delta = 46'sb1111111111111111111111111111111111111101000000;
		320: Delta = 46'sb0000000000000000000000000000000000000101000000;
		18293: Delta = 46'sb1111111111111111111111111111111111111011000000;
		576: Delta = 46'sb0000000000000000000000000000000000001001000000;
		18165: Delta = 46'sb1111111111111111111111111111111111111001000000;
		448: Delta = 46'sb0000000000000000000000000000000000000111000000;
		18037: Delta = 46'sb1111111111111111111111111111111111110111000000;
		1088: Delta = 46'sb0000000000000000000000000000000000010001000000;
		17653: Delta = 46'sb1111111111111111111111111111111111110001000000;
		960: Delta = 46'sb0000000000000000000000000000000000001111000000;
		17525: Delta = 46'sb1111111111111111111111111111111111101111000000;
		2112: Delta = 46'sb0000000000000000000000000000000000100001000000;
		16629: Delta = 46'sb1111111111111111111111111111111111100001000000;
		1984: Delta = 46'sb0000000000000000000000000000000000011111000000;
		16501: Delta = 46'sb1111111111111111111111111111111111011111000000;
		4160: Delta = 46'sb0000000000000000000000000000000001000001000000;
		14581: Delta = 46'sb1111111111111111111111111111111111000001000000;
		4032: Delta = 46'sb0000000000000000000000000000000000111111000000;
		14453: Delta = 46'sb1111111111111111111111111111111110111111000000;
		8256: Delta = 46'sb0000000000000000000000000000000010000001000000;
		10485: Delta = 46'sb1111111111111111111111111111111110000001000000;
		8128: Delta = 46'sb0000000000000000000000000000000001111111000000;
		10357: Delta = 46'sb1111111111111111111111111111111101111111000000;
		16448: Delta = 46'sb0000000000000000000000000000000100000001000000;
		2293: Delta = 46'sb1111111111111111111111111111111100000001000000;
		16320: Delta = 46'sb0000000000000000000000000000000011111111000000;
		2165: Delta = 46'sb1111111111111111111111111111111011111111000000;
		14219: Delta = 46'sb0000000000000000000000000000001000000001000000;
		4522: Delta = 46'sb1111111111111111111111111111111000000001000000;
		14091: Delta = 46'sb0000000000000000000000000000000111111111000000;
		4394: Delta = 46'sb1111111111111111111111111111110111111111000000;
		9761: Delta = 46'sb0000000000000000000000000000010000000001000000;
		8980: Delta = 46'sb1111111111111111111111111111110000000001000000;
		9633: Delta = 46'sb0000000000000000000000000000001111111111000000;
		8852: Delta = 46'sb1111111111111111111111111111101111111111000000;
		845: Delta = 46'sb0000000000000000000000000000100000000001000000;
		17896: Delta = 46'sb1111111111111111111111111111100000000001000000;
		717: Delta = 46'sb0000000000000000000000000000011111111111000000;
		17768: Delta = 46'sb1111111111111111111111111111011111111111000000;
		1626: Delta = 46'sb0000000000000000000000000001000000000001000000;
		17115: Delta = 46'sb1111111111111111111111111111000000000001000000;
		1498: Delta = 46'sb0000000000000000000000000000111111111111000000;
		16987: Delta = 46'sb1111111111111111111111111110111111111111000000;
		3188: Delta = 46'sb0000000000000000000000000010000000000001000000;
		15553: Delta = 46'sb1111111111111111111111111110000000000001000000;
		3060: Delta = 46'sb0000000000000000000000000001111111111111000000;
		15425: Delta = 46'sb1111111111111111111111111101111111111111000000;
		6312: Delta = 46'sb0000000000000000000000000100000000000001000000;
		12429: Delta = 46'sb1111111111111111111111111100000000000001000000;
		6184: Delta = 46'sb0000000000000000000000000011111111111111000000;
		12301: Delta = 46'sb1111111111111111111111111011111111111111000000;
		12560: Delta = 46'sb0000000000000000000000001000000000000001000000;
		6181: Delta = 46'sb1111111111111111111111111000000000000001000000;
		12432: Delta = 46'sb0000000000000000000000000111111111111111000000;
		6053: Delta = 46'sb1111111111111111111111110111111111111111000000;
		6443: Delta = 46'sb0000000000000000000000010000000000000001000000;
		12298: Delta = 46'sb1111111111111111111111110000000000000001000000;
		6315: Delta = 46'sb0000000000000000000000001111111111111111000000;
		12170: Delta = 46'sb1111111111111111111111101111111111111111000000;
		12822: Delta = 46'sb0000000000000000000000100000000000000001000000;
		5919: Delta = 46'sb1111111111111111111111100000000000000001000000;
		12694: Delta = 46'sb0000000000000000000000011111111111111111000000;
		5791: Delta = 46'sb1111111111111111111111011111111111111111000000;
		6967: Delta = 46'sb0000000000000000000001000000000000000001000000;
		11774: Delta = 46'sb1111111111111111111111000000000000000001000000;
		6839: Delta = 46'sb0000000000000000000000111111111111111111000000;
		11646: Delta = 46'sb1111111111111111111110111111111111111111000000;
		13870: Delta = 46'sb0000000000000000000010000000000000000001000000;
		4871: Delta = 46'sb1111111111111111111110000000000000000001000000;
		13742: Delta = 46'sb0000000000000000000001111111111111111111000000;
		4743: Delta = 46'sb1111111111111111111101111111111111111111000000;
		9063: Delta = 46'sb0000000000000000000100000000000000000001000000;
		9678: Delta = 46'sb1111111111111111111100000000000000000001000000;
		8935: Delta = 46'sb0000000000000000000011111111111111111111000000;
		9550: Delta = 46'sb1111111111111111111011111111111111111111000000;
		18062: Delta = 46'sb0000000000000000001000000000000000000001000000;
		679: Delta = 46'sb1111111111111111111000000000000000000001000000;
		17934: Delta = 46'sb0000000000000000000111111111111111111111000000;
		551: Delta = 46'sb1111111111111111110111111111111111111111000000;
		17447: Delta = 46'sb0000000000000000010000000000000000000001000000;
		1294: Delta = 46'sb1111111111111111110000000000000000000001000000;
		17319: Delta = 46'sb0000000000000000001111111111111111111111000000;
		1166: Delta = 46'sb1111111111111111101111111111111111111111000000;
		16217: Delta = 46'sb0000000000000000100000000000000000000001000000;
		2524: Delta = 46'sb1111111111111111100000000000000000000001000000;
		16089: Delta = 46'sb0000000000000000011111111111111111111111000000;
		2396: Delta = 46'sb1111111111111111011111111111111111111111000000;
		13757: Delta = 46'sb0000000000000001000000000000000000000001000000;
		4984: Delta = 46'sb1111111111111111000000000000000000000001000000;
		13629: Delta = 46'sb0000000000000000111111111111111111111111000000;
		4856: Delta = 46'sb1111111111111110111111111111111111111111000000;
		8837: Delta = 46'sb0000000000000010000000000000000000000001000000;
		9904: Delta = 46'sb1111111111111110000000000000000000000001000000;
		8709: Delta = 46'sb0000000000000001111111111111111111111111000000;
		9776: Delta = 46'sb1111111111111101111111111111111111111111000000;
		17610: Delta = 46'sb0000000000000100000000000000000000000001000000;
		1131: Delta = 46'sb1111111111111100000000000000000000000001000000;
		17482: Delta = 46'sb0000000000000011111111111111111111111111000000;
		1003: Delta = 46'sb1111111111111011111111111111111111111111000000;
		16543: Delta = 46'sb0000000000001000000000000000000000000001000000;
		2198: Delta = 46'sb1111111111111000000000000000000000000001000000;
		16415: Delta = 46'sb0000000000000111111111111111111111111111000000;
		2070: Delta = 46'sb1111111111110111111111111111111111111111000000;
		14409: Delta = 46'sb0000000000010000000000000000000000000001000000;
		4332: Delta = 46'sb1111111111110000000000000000000000000001000000;
		14281: Delta = 46'sb0000000000001111111111111111111111111111000000;
		4204: Delta = 46'sb1111111111101111111111111111111111111111000000;
		10141: Delta = 46'sb0000000000100000000000000000000000000001000000;
		8600: Delta = 46'sb1111111111100000000000000000000000000001000000;
		10013: Delta = 46'sb0000000000011111111111111111111111111111000000;
		8472: Delta = 46'sb1111111111011111111111111111111111111111000000;
		1605: Delta = 46'sb0000000001000000000000000000000000000001000000;
		17136: Delta = 46'sb1111111111000000000000000000000000000001000000;
		1477: Delta = 46'sb0000000000111111111111111111111111111111000000;
		17008: Delta = 46'sb1111111110111111111111111111111111111111000000;
		3146: Delta = 46'sb0000000010000000000000000000000000000001000000;
		15595: Delta = 46'sb1111111110000000000000000000000000000001000000;
		3018: Delta = 46'sb0000000001111111111111111111111111111111000000;
		15467: Delta = 46'sb1111111101111111111111111111111111111111000000;
		6228: Delta = 46'sb0000000100000000000000000000000000000001000000;
		12513: Delta = 46'sb1111111100000000000000000000000000000001000000;
		6100: Delta = 46'sb0000000011111111111111111111111111111111000000;
		12385: Delta = 46'sb1111111011111111111111111111111111111111000000;
		12392: Delta = 46'sb0000001000000000000000000000000000000001000000;
		6349: Delta = 46'sb1111111000000000000000000000000000000001000000;
		12264: Delta = 46'sb0000000111111111111111111111111111111111000000;
		6221: Delta = 46'sb1111110111111111111111111111111111111111000000;
		6107: Delta = 46'sb0000010000000000000000000000000000000001000000;
		12634: Delta = 46'sb1111110000000000000000000000000000000001000000;
		5979: Delta = 46'sb0000001111111111111111111111111111111111000000;
		12506: Delta = 46'sb1111101111111111111111111111111111111111000000;
		12150: Delta = 46'sb0000100000000000000000000000000000000001000000;
		6591: Delta = 46'sb1111100000000000000000000000000000000001000000;
		12022: Delta = 46'sb0000011111111111111111111111111111111111000000;
		6463: Delta = 46'sb1111011111111111111111111111111111111111000000;
		5623: Delta = 46'sb0001000000000000000000000000000000000001000000;
		13118: Delta = 46'sb1111000000000000000000000000000000000001000000;
		5495: Delta = 46'sb0000111111111111111111111111111111111111000000;
		12990: Delta = 46'sb1110111111111111111111111111111111111111000000;
		11182: Delta = 46'sb0010000000000000000000000000000000000001000000;
		7559: Delta = 46'sb1110000000000000000000000000000000000001000000;
		11054: Delta = 46'sb0001111111111111111111111111111111111111000000;
		7431: Delta = 46'sb1101111111111111111111111111111111111111000000;
		3687: Delta = 46'sb0100000000000000000000000000000000000001000000;
		15054: Delta = 46'sb1100000000000000000000000000000000000001000000;
		3559: Delta = 46'sb0011111111111111111111111111111111111111000000;
		14926: Delta = 46'sb1011111111111111111111111111111111111111000000;
		384: Delta = 46'sb0000000000000000000000000000000000000110000000;
		18229: Delta = 46'sb1111111111111111111111111111111111111010000000;
		640: Delta = 46'sb0000000000000000000000000000000000001010000000;
		17973: Delta = 46'sb1111111111111111111111111111111111110110000000;
		1152: Delta = 46'sb0000000000000000000000000000000000010010000000;
		17717: Delta = 46'sb1111111111111111111111111111111111110010000000;
		896: Delta = 46'sb0000000000000000000000000000000000001110000000;
		17461: Delta = 46'sb1111111111111111111111111111111111101110000000;
		2176: Delta = 46'sb0000000000000000000000000000000000100010000000;
		16693: Delta = 46'sb1111111111111111111111111111111111100010000000;
		1920: Delta = 46'sb0000000000000000000000000000000000011110000000;
		16437: Delta = 46'sb1111111111111111111111111111111111011110000000;
		4224: Delta = 46'sb0000000000000000000000000000000001000010000000;
		14645: Delta = 46'sb1111111111111111111111111111111111000010000000;
		3968: Delta = 46'sb0000000000000000000000000000000000111110000000;
		14389: Delta = 46'sb1111111111111111111111111111111110111110000000;
		8320: Delta = 46'sb0000000000000000000000000000000010000010000000;
		10549: Delta = 46'sb1111111111111111111111111111111110000010000000;
		8064: Delta = 46'sb0000000000000000000000000000000001111110000000;
		10293: Delta = 46'sb1111111111111111111111111111111101111110000000;
		16512: Delta = 46'sb0000000000000000000000000000000100000010000000;
		2357: Delta = 46'sb1111111111111111111111111111111100000010000000;
		16256: Delta = 46'sb0000000000000000000000000000000011111110000000;
		2101: Delta = 46'sb1111111111111111111111111111111011111110000000;
		14283: Delta = 46'sb0000000000000000000000000000001000000010000000;
		4586: Delta = 46'sb1111111111111111111111111111111000000010000000;
		14027: Delta = 46'sb0000000000000000000000000000000111111110000000;
		4330: Delta = 46'sb1111111111111111111111111111110111111110000000;
		9825: Delta = 46'sb0000000000000000000000000000010000000010000000;
		9044: Delta = 46'sb1111111111111111111111111111110000000010000000;
		9569: Delta = 46'sb0000000000000000000000000000001111111110000000;
		8788: Delta = 46'sb1111111111111111111111111111101111111110000000;
		909: Delta = 46'sb0000000000000000000000000000100000000010000000;
		17960: Delta = 46'sb1111111111111111111111111111100000000010000000;
		653: Delta = 46'sb0000000000000000000000000000011111111110000000;
		17704: Delta = 46'sb1111111111111111111111111111011111111110000000;
		1690: Delta = 46'sb0000000000000000000000000001000000000010000000;
		17179: Delta = 46'sb1111111111111111111111111111000000000010000000;
		1434: Delta = 46'sb0000000000000000000000000000111111111110000000;
		16923: Delta = 46'sb1111111111111111111111111110111111111110000000;
		3252: Delta = 46'sb0000000000000000000000000010000000000010000000;
		15617: Delta = 46'sb1111111111111111111111111110000000000010000000;
		2996: Delta = 46'sb0000000000000000000000000001111111111110000000;
		15361: Delta = 46'sb1111111111111111111111111101111111111110000000;
		6376: Delta = 46'sb0000000000000000000000000100000000000010000000;
		12493: Delta = 46'sb1111111111111111111111111100000000000010000000;
		6120: Delta = 46'sb0000000000000000000000000011111111111110000000;
		12237: Delta = 46'sb1111111111111111111111111011111111111110000000;
		12624: Delta = 46'sb0000000000000000000000001000000000000010000000;
		6245: Delta = 46'sb1111111111111111111111111000000000000010000000;
		12368: Delta = 46'sb0000000000000000000000000111111111111110000000;
		5989: Delta = 46'sb1111111111111111111111110111111111111110000000;
		6507: Delta = 46'sb0000000000000000000000010000000000000010000000;
		12362: Delta = 46'sb1111111111111111111111110000000000000010000000;
		6251: Delta = 46'sb0000000000000000000000001111111111111110000000;
		12106: Delta = 46'sb1111111111111111111111101111111111111110000000;
		12886: Delta = 46'sb0000000000000000000000100000000000000010000000;
		5983: Delta = 46'sb1111111111111111111111100000000000000010000000;
		12630: Delta = 46'sb0000000000000000000000011111111111111110000000;
		5727: Delta = 46'sb1111111111111111111111011111111111111110000000;
		7031: Delta = 46'sb0000000000000000000001000000000000000010000000;
		11838: Delta = 46'sb1111111111111111111111000000000000000010000000;
		6775: Delta = 46'sb0000000000000000000000111111111111111110000000;
		11582: Delta = 46'sb1111111111111111111110111111111111111110000000;
		13934: Delta = 46'sb0000000000000000000010000000000000000010000000;
		4935: Delta = 46'sb1111111111111111111110000000000000000010000000;
		13678: Delta = 46'sb0000000000000000000001111111111111111110000000;
		4679: Delta = 46'sb1111111111111111111101111111111111111110000000;
		9127: Delta = 46'sb0000000000000000000100000000000000000010000000;
		9742: Delta = 46'sb1111111111111111111100000000000000000010000000;
		8871: Delta = 46'sb0000000000000000000011111111111111111110000000;
		9486: Delta = 46'sb1111111111111111111011111111111111111110000000;
		18126: Delta = 46'sb0000000000000000001000000000000000000010000000;
		743: Delta = 46'sb1111111111111111111000000000000000000010000000;
		17870: Delta = 46'sb0000000000000000000111111111111111111110000000;
		487: Delta = 46'sb1111111111111111110111111111111111111110000000;
		17511: Delta = 46'sb0000000000000000010000000000000000000010000000;
		1358: Delta = 46'sb1111111111111111110000000000000000000010000000;
		17255: Delta = 46'sb0000000000000000001111111111111111111110000000;
		1102: Delta = 46'sb1111111111111111101111111111111111111110000000;
		16281: Delta = 46'sb0000000000000000100000000000000000000010000000;
		2588: Delta = 46'sb1111111111111111100000000000000000000010000000;
		16025: Delta = 46'sb0000000000000000011111111111111111111110000000;
		2332: Delta = 46'sb1111111111111111011111111111111111111110000000;
		13821: Delta = 46'sb0000000000000001000000000000000000000010000000;
		5048: Delta = 46'sb1111111111111111000000000000000000000010000000;
		13565: Delta = 46'sb0000000000000000111111111111111111111110000000;
		4792: Delta = 46'sb1111111111111110111111111111111111111110000000;
		8901: Delta = 46'sb0000000000000010000000000000000000000010000000;
		9968: Delta = 46'sb1111111111111110000000000000000000000010000000;
		8645: Delta = 46'sb0000000000000001111111111111111111111110000000;
		9712: Delta = 46'sb1111111111111101111111111111111111111110000000;
		17674: Delta = 46'sb0000000000000100000000000000000000000010000000;
		1195: Delta = 46'sb1111111111111100000000000000000000000010000000;
		17418: Delta = 46'sb0000000000000011111111111111111111111110000000;
		939: Delta = 46'sb1111111111111011111111111111111111111110000000;
		16607: Delta = 46'sb0000000000001000000000000000000000000010000000;
		2262: Delta = 46'sb1111111111111000000000000000000000000010000000;
		16351: Delta = 46'sb0000000000000111111111111111111111111110000000;
		2006: Delta = 46'sb1111111111110111111111111111111111111110000000;
		14473: Delta = 46'sb0000000000010000000000000000000000000010000000;
		4396: Delta = 46'sb1111111111110000000000000000000000000010000000;
		14217: Delta = 46'sb0000000000001111111111111111111111111110000000;
		4140: Delta = 46'sb1111111111101111111111111111111111111110000000;
		10205: Delta = 46'sb0000000000100000000000000000000000000010000000;
		8664: Delta = 46'sb1111111111100000000000000000000000000010000000;
		9949: Delta = 46'sb0000000000011111111111111111111111111110000000;
		8408: Delta = 46'sb1111111111011111111111111111111111111110000000;
		1669: Delta = 46'sb0000000001000000000000000000000000000010000000;
		17200: Delta = 46'sb1111111111000000000000000000000000000010000000;
		1413: Delta = 46'sb0000000000111111111111111111111111111110000000;
		16944: Delta = 46'sb1111111110111111111111111111111111111110000000;
		3210: Delta = 46'sb0000000010000000000000000000000000000010000000;
		15659: Delta = 46'sb1111111110000000000000000000000000000010000000;
		2954: Delta = 46'sb0000000001111111111111111111111111111110000000;
		15403: Delta = 46'sb1111111101111111111111111111111111111110000000;
		6292: Delta = 46'sb0000000100000000000000000000000000000010000000;
		12577: Delta = 46'sb1111111100000000000000000000000000000010000000;
		6036: Delta = 46'sb0000000011111111111111111111111111111110000000;
		12321: Delta = 46'sb1111111011111111111111111111111111111110000000;
		12456: Delta = 46'sb0000001000000000000000000000000000000010000000;
		6413: Delta = 46'sb1111111000000000000000000000000000000010000000;
		12200: Delta = 46'sb0000000111111111111111111111111111111110000000;
		6157: Delta = 46'sb1111110111111111111111111111111111111110000000;
		6171: Delta = 46'sb0000010000000000000000000000000000000010000000;
		12698: Delta = 46'sb1111110000000000000000000000000000000010000000;
		5915: Delta = 46'sb0000001111111111111111111111111111111110000000;
		12442: Delta = 46'sb1111101111111111111111111111111111111110000000;
		12214: Delta = 46'sb0000100000000000000000000000000000000010000000;
		6655: Delta = 46'sb1111100000000000000000000000000000000010000000;
		11958: Delta = 46'sb0000011111111111111111111111111111111110000000;
		6399: Delta = 46'sb1111011111111111111111111111111111111110000000;
		5687: Delta = 46'sb0001000000000000000000000000000000000010000000;
		13182: Delta = 46'sb1111000000000000000000000000000000000010000000;
		5431: Delta = 46'sb0000111111111111111111111111111111111110000000;
		12926: Delta = 46'sb1110111111111111111111111111111111111110000000;
		11246: Delta = 46'sb0010000000000000000000000000000000000010000000;
		7623: Delta = 46'sb1110000000000000000000000000000000000010000000;
		10990: Delta = 46'sb0001111111111111111111111111111111111110000000;
		7367: Delta = 46'sb1101111111111111111111111111111111111110000000;
		3751: Delta = 46'sb0100000000000000000000000000000000000010000000;
		15118: Delta = 46'sb1100000000000000000000000000000000000010000000;
		3495: Delta = 46'sb0011111111111111111111111111111111111110000000;
		14862: Delta = 46'sb1011111111111111111111111111111111111110000000;
		768: Delta = 46'sb0000000000000000000000000000000000001100000000;
		17845: Delta = 46'sb1111111111111111111111111111111111110100000000;
		1280: Delta = 46'sb0000000000000000000000000000000000010100000000;
		17333: Delta = 46'sb1111111111111111111111111111111111101100000000;
		2304: Delta = 46'sb0000000000000000000000000000000000100100000000;
		16821: Delta = 46'sb1111111111111111111111111111111111100100000000;
		1792: Delta = 46'sb0000000000000000000000000000000000011100000000;
		16309: Delta = 46'sb1111111111111111111111111111111111011100000000;
		4352: Delta = 46'sb0000000000000000000000000000000001000100000000;
		14773: Delta = 46'sb1111111111111111111111111111111111000100000000;
		3840: Delta = 46'sb0000000000000000000000000000000000111100000000;
		14261: Delta = 46'sb1111111111111111111111111111111110111100000000;
		8448: Delta = 46'sb0000000000000000000000000000000010000100000000;
		10677: Delta = 46'sb1111111111111111111111111111111110000100000000;
		7936: Delta = 46'sb0000000000000000000000000000000001111100000000;
		10165: Delta = 46'sb1111111111111111111111111111111101111100000000;
		16640: Delta = 46'sb0000000000000000000000000000000100000100000000;
		2485: Delta = 46'sb1111111111111111111111111111111100000100000000;
		16128: Delta = 46'sb0000000000000000000000000000000011111100000000;
		1973: Delta = 46'sb1111111111111111111111111111111011111100000000;
		14411: Delta = 46'sb0000000000000000000000000000001000000100000000;
		4714: Delta = 46'sb1111111111111111111111111111111000000100000000;
		13899: Delta = 46'sb0000000000000000000000000000000111111100000000;
		4202: Delta = 46'sb1111111111111111111111111111110111111100000000;
		9953: Delta = 46'sb0000000000000000000000000000010000000100000000;
		9172: Delta = 46'sb1111111111111111111111111111110000000100000000;
		9441: Delta = 46'sb0000000000000000000000000000001111111100000000;
		8660: Delta = 46'sb1111111111111111111111111111101111111100000000;
		1037: Delta = 46'sb0000000000000000000000000000100000000100000000;
		18088: Delta = 46'sb1111111111111111111111111111100000000100000000;
		525: Delta = 46'sb0000000000000000000000000000011111111100000000;
		17576: Delta = 46'sb1111111111111111111111111111011111111100000000;
		1818: Delta = 46'sb0000000000000000000000000001000000000100000000;
		17307: Delta = 46'sb1111111111111111111111111111000000000100000000;
		1306: Delta = 46'sb0000000000000000000000000000111111111100000000;
		16795: Delta = 46'sb1111111111111111111111111110111111111100000000;
		3380: Delta = 46'sb0000000000000000000000000010000000000100000000;
		15745: Delta = 46'sb1111111111111111111111111110000000000100000000;
		2868: Delta = 46'sb0000000000000000000000000001111111111100000000;
		15233: Delta = 46'sb1111111111111111111111111101111111111100000000;
		6504: Delta = 46'sb0000000000000000000000000100000000000100000000;
		12621: Delta = 46'sb1111111111111111111111111100000000000100000000;
		5992: Delta = 46'sb0000000000000000000000000011111111111100000000;
		12109: Delta = 46'sb1111111111111111111111111011111111111100000000;
		12752: Delta = 46'sb0000000000000000000000001000000000000100000000;
		6373: Delta = 46'sb1111111111111111111111111000000000000100000000;
		12240: Delta = 46'sb0000000000000000000000000111111111111100000000;
		5861: Delta = 46'sb1111111111111111111111110111111111111100000000;
		6635: Delta = 46'sb0000000000000000000000010000000000000100000000;
		12490: Delta = 46'sb1111111111111111111111110000000000000100000000;
		6123: Delta = 46'sb0000000000000000000000001111111111111100000000;
		11978: Delta = 46'sb1111111111111111111111101111111111111100000000;
		13014: Delta = 46'sb0000000000000000000000100000000000000100000000;
		6111: Delta = 46'sb1111111111111111111111100000000000000100000000;
		12502: Delta = 46'sb0000000000000000000000011111111111111100000000;
		5599: Delta = 46'sb1111111111111111111111011111111111111100000000;
		7159: Delta = 46'sb0000000000000000000001000000000000000100000000;
		11966: Delta = 46'sb1111111111111111111111000000000000000100000000;
		6647: Delta = 46'sb0000000000000000000000111111111111111100000000;
		11454: Delta = 46'sb1111111111111111111110111111111111111100000000;
		14062: Delta = 46'sb0000000000000000000010000000000000000100000000;
		5063: Delta = 46'sb1111111111111111111110000000000000000100000000;
		13550: Delta = 46'sb0000000000000000000001111111111111111100000000;
		4551: Delta = 46'sb1111111111111111111101111111111111111100000000;
		9255: Delta = 46'sb0000000000000000000100000000000000000100000000;
		9870: Delta = 46'sb1111111111111111111100000000000000000100000000;
		8743: Delta = 46'sb0000000000000000000011111111111111111100000000;
		9358: Delta = 46'sb1111111111111111111011111111111111111100000000;
		18254: Delta = 46'sb0000000000000000001000000000000000000100000000;
		871: Delta = 46'sb1111111111111111111000000000000000000100000000;
		17742: Delta = 46'sb0000000000000000000111111111111111111100000000;
		359: Delta = 46'sb1111111111111111110111111111111111111100000000;
		17639: Delta = 46'sb0000000000000000010000000000000000000100000000;
		1486: Delta = 46'sb1111111111111111110000000000000000000100000000;
		17127: Delta = 46'sb0000000000000000001111111111111111111100000000;
		974: Delta = 46'sb1111111111111111101111111111111111111100000000;
		16409: Delta = 46'sb0000000000000000100000000000000000000100000000;
		2716: Delta = 46'sb1111111111111111100000000000000000000100000000;
		15897: Delta = 46'sb0000000000000000011111111111111111111100000000;
		2204: Delta = 46'sb1111111111111111011111111111111111111100000000;
		13949: Delta = 46'sb0000000000000001000000000000000000000100000000;
		5176: Delta = 46'sb1111111111111111000000000000000000000100000000;
		13437: Delta = 46'sb0000000000000000111111111111111111111100000000;
		4664: Delta = 46'sb1111111111111110111111111111111111111100000000;
		9029: Delta = 46'sb0000000000000010000000000000000000000100000000;
		10096: Delta = 46'sb1111111111111110000000000000000000000100000000;
		8517: Delta = 46'sb0000000000000001111111111111111111111100000000;
		9584: Delta = 46'sb1111111111111101111111111111111111111100000000;
		17802: Delta = 46'sb0000000000000100000000000000000000000100000000;
		1323: Delta = 46'sb1111111111111100000000000000000000000100000000;
		17290: Delta = 46'sb0000000000000011111111111111111111111100000000;
		811: Delta = 46'sb1111111111111011111111111111111111111100000000;
		16735: Delta = 46'sb0000000000001000000000000000000000000100000000;
		2390: Delta = 46'sb1111111111111000000000000000000000000100000000;
		16223: Delta = 46'sb0000000000000111111111111111111111111100000000;
		1878: Delta = 46'sb1111111111110111111111111111111111111100000000;
		14601: Delta = 46'sb0000000000010000000000000000000000000100000000;
		4524: Delta = 46'sb1111111111110000000000000000000000000100000000;
		14089: Delta = 46'sb0000000000001111111111111111111111111100000000;
		4012: Delta = 46'sb1111111111101111111111111111111111111100000000;
		10333: Delta = 46'sb0000000000100000000000000000000000000100000000;
		8792: Delta = 46'sb1111111111100000000000000000000000000100000000;
		9821: Delta = 46'sb0000000000011111111111111111111111111100000000;
		8280: Delta = 46'sb1111111111011111111111111111111111111100000000;
		1797: Delta = 46'sb0000000001000000000000000000000000000100000000;
		17328: Delta = 46'sb1111111111000000000000000000000000000100000000;
		1285: Delta = 46'sb0000000000111111111111111111111111111100000000;
		16816: Delta = 46'sb1111111110111111111111111111111111111100000000;
		3338: Delta = 46'sb0000000010000000000000000000000000000100000000;
		15787: Delta = 46'sb1111111110000000000000000000000000000100000000;
		2826: Delta = 46'sb0000000001111111111111111111111111111100000000;
		15275: Delta = 46'sb1111111101111111111111111111111111111100000000;
		6420: Delta = 46'sb0000000100000000000000000000000000000100000000;
		12705: Delta = 46'sb1111111100000000000000000000000000000100000000;
		5908: Delta = 46'sb0000000011111111111111111111111111111100000000;
		12193: Delta = 46'sb1111111011111111111111111111111111111100000000;
		12584: Delta = 46'sb0000001000000000000000000000000000000100000000;
		6541: Delta = 46'sb1111111000000000000000000000000000000100000000;
		12072: Delta = 46'sb0000000111111111111111111111111111111100000000;
		6029: Delta = 46'sb1111110111111111111111111111111111111100000000;
		6299: Delta = 46'sb0000010000000000000000000000000000000100000000;
		12826: Delta = 46'sb1111110000000000000000000000000000000100000000;
		5787: Delta = 46'sb0000001111111111111111111111111111111100000000;
		12314: Delta = 46'sb1111101111111111111111111111111111111100000000;
		12342: Delta = 46'sb0000100000000000000000000000000000000100000000;
		6783: Delta = 46'sb1111100000000000000000000000000000000100000000;
		11830: Delta = 46'sb0000011111111111111111111111111111111100000000;
		6271: Delta = 46'sb1111011111111111111111111111111111111100000000;
		5815: Delta = 46'sb0001000000000000000000000000000000000100000000;
		13310: Delta = 46'sb1111000000000000000000000000000000000100000000;
		5303: Delta = 46'sb0000111111111111111111111111111111111100000000;
		12798: Delta = 46'sb1110111111111111111111111111111111111100000000;
		11374: Delta = 46'sb0010000000000000000000000000000000000100000000;
		7751: Delta = 46'sb1110000000000000000000000000000000000100000000;
		10862: Delta = 46'sb0001111111111111111111111111111111111100000000;
		7239: Delta = 46'sb1101111111111111111111111111111111111100000000;
		3879: Delta = 46'sb0100000000000000000000000000000000000100000000;
		15246: Delta = 46'sb1100000000000000000000000000000000000100000000;
		3367: Delta = 46'sb0011111111111111111111111111111111111100000000;
		14734: Delta = 46'sb1011111111111111111111111111111111111100000000;
		1536: Delta = 46'sb0000000000000000000000000000000000011000000000;
		17077: Delta = 46'sb1111111111111111111111111111111111101000000000;
		2560: Delta = 46'sb0000000000000000000000000000000000101000000000;
		16053: Delta = 46'sb1111111111111111111111111111111111011000000000;
		4608: Delta = 46'sb0000000000000000000000000000000001001000000000;
		15029: Delta = 46'sb1111111111111111111111111111111111001000000000;
		3584: Delta = 46'sb0000000000000000000000000000000000111000000000;
		14005: Delta = 46'sb1111111111111111111111111111111110111000000000;
		8704: Delta = 46'sb0000000000000000000000000000000010001000000000;
		10933: Delta = 46'sb1111111111111111111111111111111110001000000000;
		7680: Delta = 46'sb0000000000000000000000000000000001111000000000;
		9909: Delta = 46'sb1111111111111111111111111111111101111000000000;
		16896: Delta = 46'sb0000000000000000000000000000000100001000000000;
		2741: Delta = 46'sb1111111111111111111111111111111100001000000000;
		15872: Delta = 46'sb0000000000000000000000000000000011111000000000;
		1717: Delta = 46'sb1111111111111111111111111111111011111000000000;
		14667: Delta = 46'sb0000000000000000000000000000001000001000000000;
		4970: Delta = 46'sb1111111111111111111111111111111000001000000000;
		13643: Delta = 46'sb0000000000000000000000000000000111111000000000;
		3946: Delta = 46'sb1111111111111111111111111111110111111000000000;
		10209: Delta = 46'sb0000000000000000000000000000010000001000000000;
		9428: Delta = 46'sb1111111111111111111111111111110000001000000000;
		9185: Delta = 46'sb0000000000000000000000000000001111111000000000;
		8404: Delta = 46'sb1111111111111111111111111111101111111000000000;
		1293: Delta = 46'sb0000000000000000000000000000100000001000000000;
		18344: Delta = 46'sb1111111111111111111111111111100000001000000000;
		269: Delta = 46'sb0000000000000000000000000000011111111000000000;
		17320: Delta = 46'sb1111111111111111111111111111011111111000000000;
		2074: Delta = 46'sb0000000000000000000000000001000000001000000000;
		17563: Delta = 46'sb1111111111111111111111111111000000001000000000;
		1050: Delta = 46'sb0000000000000000000000000000111111111000000000;
		16539: Delta = 46'sb1111111111111111111111111110111111111000000000;
		3636: Delta = 46'sb0000000000000000000000000010000000001000000000;
		16001: Delta = 46'sb1111111111111111111111111110000000001000000000;
		2612: Delta = 46'sb0000000000000000000000000001111111111000000000;
		14977: Delta = 46'sb1111111111111111111111111101111111111000000000;
		6760: Delta = 46'sb0000000000000000000000000100000000001000000000;
		12877: Delta = 46'sb1111111111111111111111111100000000001000000000;
		5736: Delta = 46'sb0000000000000000000000000011111111111000000000;
		11853: Delta = 46'sb1111111111111111111111111011111111111000000000;
		13008: Delta = 46'sb0000000000000000000000001000000000001000000000;
		6629: Delta = 46'sb1111111111111111111111111000000000001000000000;
		11984: Delta = 46'sb0000000000000000000000000111111111111000000000;
		5605: Delta = 46'sb1111111111111111111111110111111111111000000000;
		6891: Delta = 46'sb0000000000000000000000010000000000001000000000;
		12746: Delta = 46'sb1111111111111111111111110000000000001000000000;
		5867: Delta = 46'sb0000000000000000000000001111111111111000000000;
		11722: Delta = 46'sb1111111111111111111111101111111111111000000000;
		13270: Delta = 46'sb0000000000000000000000100000000000001000000000;
		6367: Delta = 46'sb1111111111111111111111100000000000001000000000;
		12246: Delta = 46'sb0000000000000000000000011111111111111000000000;
		5343: Delta = 46'sb1111111111111111111111011111111111111000000000;
		7415: Delta = 46'sb0000000000000000000001000000000000001000000000;
		12222: Delta = 46'sb1111111111111111111111000000000000001000000000;
		6391: Delta = 46'sb0000000000000000000000111111111111111000000000;
		11198: Delta = 46'sb1111111111111111111110111111111111111000000000;
		14318: Delta = 46'sb0000000000000000000010000000000000001000000000;
		5319: Delta = 46'sb1111111111111111111110000000000000001000000000;
		13294: Delta = 46'sb0000000000000000000001111111111111111000000000;
		4295: Delta = 46'sb1111111111111111111101111111111111111000000000;
		9511: Delta = 46'sb0000000000000000000100000000000000001000000000;
		10126: Delta = 46'sb1111111111111111111100000000000000001000000000;
		8487: Delta = 46'sb0000000000000000000011111111111111111000000000;
		9102: Delta = 46'sb1111111111111111111011111111111111111000000000;
		18510: Delta = 46'sb0000000000000000001000000000000000001000000000;
		1127: Delta = 46'sb1111111111111111111000000000000000001000000000;
		17486: Delta = 46'sb0000000000000000000111111111111111111000000000;
		103: Delta = 46'sb1111111111111111110111111111111111111000000000;
		17895: Delta = 46'sb0000000000000000010000000000000000001000000000;
		1742: Delta = 46'sb1111111111111111110000000000000000001000000000;
		16871: Delta = 46'sb0000000000000000001111111111111111111000000000;
		718: Delta = 46'sb1111111111111111101111111111111111111000000000;
		16665: Delta = 46'sb0000000000000000100000000000000000001000000000;
		2972: Delta = 46'sb1111111111111111100000000000000000001000000000;
		15641: Delta = 46'sb0000000000000000011111111111111111111000000000;
		1948: Delta = 46'sb1111111111111111011111111111111111111000000000;
		14205: Delta = 46'sb0000000000000001000000000000000000001000000000;
		5432: Delta = 46'sb1111111111111111000000000000000000001000000000;
		13181: Delta = 46'sb0000000000000000111111111111111111111000000000;
		4408: Delta = 46'sb1111111111111110111111111111111111111000000000;
		9285: Delta = 46'sb0000000000000010000000000000000000001000000000;
		10352: Delta = 46'sb1111111111111110000000000000000000001000000000;
		8261: Delta = 46'sb0000000000000001111111111111111111111000000000;
		9328: Delta = 46'sb1111111111111101111111111111111111111000000000;
		18058: Delta = 46'sb0000000000000100000000000000000000001000000000;
		1579: Delta = 46'sb1111111111111100000000000000000000001000000000;
		17034: Delta = 46'sb0000000000000011111111111111111111111000000000;
		555: Delta = 46'sb1111111111111011111111111111111111111000000000;
		16991: Delta = 46'sb0000000000001000000000000000000000001000000000;
		2646: Delta = 46'sb1111111111111000000000000000000000001000000000;
		15967: Delta = 46'sb0000000000000111111111111111111111111000000000;
		1622: Delta = 46'sb1111111111110111111111111111111111111000000000;
		14857: Delta = 46'sb0000000000010000000000000000000000001000000000;
		4780: Delta = 46'sb1111111111110000000000000000000000001000000000;
		13833: Delta = 46'sb0000000000001111111111111111111111111000000000;
		3756: Delta = 46'sb1111111111101111111111111111111111111000000000;
		10589: Delta = 46'sb0000000000100000000000000000000000001000000000;
		9048: Delta = 46'sb1111111111100000000000000000000000001000000000;
		9565: Delta = 46'sb0000000000011111111111111111111111111000000000;
		8024: Delta = 46'sb1111111111011111111111111111111111111000000000;
		2053: Delta = 46'sb0000000001000000000000000000000000001000000000;
		17584: Delta = 46'sb1111111111000000000000000000000000001000000000;
		1029: Delta = 46'sb0000000000111111111111111111111111111000000000;
		16560: Delta = 46'sb1111111110111111111111111111111111111000000000;
		3594: Delta = 46'sb0000000010000000000000000000000000001000000000;
		16043: Delta = 46'sb1111111110000000000000000000000000001000000000;
		2570: Delta = 46'sb0000000001111111111111111111111111111000000000;
		15019: Delta = 46'sb1111111101111111111111111111111111111000000000;
		6676: Delta = 46'sb0000000100000000000000000000000000001000000000;
		12961: Delta = 46'sb1111111100000000000000000000000000001000000000;
		5652: Delta = 46'sb0000000011111111111111111111111111111000000000;
		11937: Delta = 46'sb1111111011111111111111111111111111111000000000;
		12840: Delta = 46'sb0000001000000000000000000000000000001000000000;
		6797: Delta = 46'sb1111111000000000000000000000000000001000000000;
		11816: Delta = 46'sb0000000111111111111111111111111111111000000000;
		5773: Delta = 46'sb1111110111111111111111111111111111111000000000;
		6555: Delta = 46'sb0000010000000000000000000000000000001000000000;
		13082: Delta = 46'sb1111110000000000000000000000000000001000000000;
		5531: Delta = 46'sb0000001111111111111111111111111111111000000000;
		12058: Delta = 46'sb1111101111111111111111111111111111111000000000;
		12598: Delta = 46'sb0000100000000000000000000000000000001000000000;
		7039: Delta = 46'sb1111100000000000000000000000000000001000000000;
		11574: Delta = 46'sb0000011111111111111111111111111111111000000000;
		6015: Delta = 46'sb1111011111111111111111111111111111111000000000;
		6071: Delta = 46'sb0001000000000000000000000000000000001000000000;
		13566: Delta = 46'sb1111000000000000000000000000000000001000000000;
		5047: Delta = 46'sb0000111111111111111111111111111111111000000000;
		12542: Delta = 46'sb1110111111111111111111111111111111111000000000;
		11630: Delta = 46'sb0010000000000000000000000000000000001000000000;
		8007: Delta = 46'sb1110000000000000000000000000000000001000000000;
		10606: Delta = 46'sb0001111111111111111111111111111111111000000000;
		6983: Delta = 46'sb1101111111111111111111111111111111111000000000;
		4135: Delta = 46'sb0100000000000000000000000000000000001000000000;
		15502: Delta = 46'sb1100000000000000000000000000000000001000000000;
		3111: Delta = 46'sb0011111111111111111111111111111111111000000000;
		14478: Delta = 46'sb1011111111111111111111111111111111111000000000;
		3072: Delta = 46'sb0000000000000000000000000000000000110000000000;
		15541: Delta = 46'sb1111111111111111111111111111111111010000000000;
		5120: Delta = 46'sb0000000000000000000000000000000001010000000000;
		13493: Delta = 46'sb1111111111111111111111111111111110110000000000;
		9216: Delta = 46'sb0000000000000000000000000000000010010000000000;
		11445: Delta = 46'sb1111111111111111111111111111111110010000000000;
		7168: Delta = 46'sb0000000000000000000000000000000001110000000000;
		9397: Delta = 46'sb1111111111111111111111111111111101110000000000;
		17408: Delta = 46'sb0000000000000000000000000000000100010000000000;
		3253: Delta = 46'sb1111111111111111111111111111111100010000000000;
		15360: Delta = 46'sb0000000000000000000000000000000011110000000000;
		1205: Delta = 46'sb1111111111111111111111111111111011110000000000;
		15179: Delta = 46'sb0000000000000000000000000000001000010000000000;
		5482: Delta = 46'sb1111111111111111111111111111111000010000000000;
		13131: Delta = 46'sb0000000000000000000000000000000111110000000000;
		3434: Delta = 46'sb1111111111111111111111111111110111110000000000;
		10721: Delta = 46'sb0000000000000000000000000000010000010000000000;
		9940: Delta = 46'sb1111111111111111111111111111110000010000000000;
		8673: Delta = 46'sb0000000000000000000000000000001111110000000000;
		7892: Delta = 46'sb1111111111111111111111111111101111110000000000;
		1805: Delta = 46'sb0000000000000000000000000000100000010000000000;
		243: Delta = 46'sb1111111111111111111111111111100000010000000000;
		18370: Delta = 46'sb0000000000000000000000000000011111110000000000;
		16808: Delta = 46'sb1111111111111111111111111111011111110000000000;
		2586: Delta = 46'sb0000000000000000000000000001000000010000000000;
		18075: Delta = 46'sb1111111111111111111111111111000000010000000000;
		538: Delta = 46'sb0000000000000000000000000000111111110000000000;
		16027: Delta = 46'sb1111111111111111111111111110111111110000000000;
		4148: Delta = 46'sb0000000000000000000000000010000000010000000000;
		16513: Delta = 46'sb1111111111111111111111111110000000010000000000;
		2100: Delta = 46'sb0000000000000000000000000001111111110000000000;
		14465: Delta = 46'sb1111111111111111111111111101111111110000000000;
		7272: Delta = 46'sb0000000000000000000000000100000000010000000000;
		13389: Delta = 46'sb1111111111111111111111111100000000010000000000;
		5224: Delta = 46'sb0000000000000000000000000011111111110000000000;
		11341: Delta = 46'sb1111111111111111111111111011111111110000000000;
		13520: Delta = 46'sb0000000000000000000000001000000000010000000000;
		7141: Delta = 46'sb1111111111111111111111111000000000010000000000;
		11472: Delta = 46'sb0000000000000000000000000111111111110000000000;
		5093: Delta = 46'sb1111111111111111111111110111111111110000000000;
		7403: Delta = 46'sb0000000000000000000000010000000000010000000000;
		13258: Delta = 46'sb1111111111111111111111110000000000010000000000;
		5355: Delta = 46'sb0000000000000000000000001111111111110000000000;
		11210: Delta = 46'sb1111111111111111111111101111111111110000000000;
		13782: Delta = 46'sb0000000000000000000000100000000000010000000000;
		6879: Delta = 46'sb1111111111111111111111100000000000010000000000;
		11734: Delta = 46'sb0000000000000000000000011111111111110000000000;
		4831: Delta = 46'sb1111111111111111111111011111111111110000000000;
		7927: Delta = 46'sb0000000000000000000001000000000000010000000000;
		12734: Delta = 46'sb1111111111111111111111000000000000010000000000;
		5879: Delta = 46'sb0000000000000000000000111111111111110000000000;
		10686: Delta = 46'sb1111111111111111111110111111111111110000000000;
		14830: Delta = 46'sb0000000000000000000010000000000000010000000000;
		5831: Delta = 46'sb1111111111111111111110000000000000010000000000;
		12782: Delta = 46'sb0000000000000000000001111111111111110000000000;
		3783: Delta = 46'sb1111111111111111111101111111111111110000000000;
		10023: Delta = 46'sb0000000000000000000100000000000000010000000000;
		10638: Delta = 46'sb1111111111111111111100000000000000010000000000;
		7975: Delta = 46'sb0000000000000000000011111111111111110000000000;
		8590: Delta = 46'sb1111111111111111111011111111111111110000000000;
		409: Delta = 46'sb0000000000000000001000000000000000010000000000;
		1639: Delta = 46'sb1111111111111111111000000000000000010000000000;
		16974: Delta = 46'sb0000000000000000000111111111111111110000000000;
		18204: Delta = 46'sb1111111111111111110111111111111111110000000000;
		18407: Delta = 46'sb0000000000000000010000000000000000010000000000;
		2254: Delta = 46'sb1111111111111111110000000000000000010000000000;
		16359: Delta = 46'sb0000000000000000001111111111111111110000000000;
		206: Delta = 46'sb1111111111111111101111111111111111110000000000;
		17177: Delta = 46'sb0000000000000000100000000000000000010000000000;
		3484: Delta = 46'sb1111111111111111100000000000000000010000000000;
		15129: Delta = 46'sb0000000000000000011111111111111111110000000000;
		1436: Delta = 46'sb1111111111111111011111111111111111110000000000;
		14717: Delta = 46'sb0000000000000001000000000000000000010000000000;
		5944: Delta = 46'sb1111111111111111000000000000000000010000000000;
		12669: Delta = 46'sb0000000000000000111111111111111111110000000000;
		3896: Delta = 46'sb1111111111111110111111111111111111110000000000;
		9797: Delta = 46'sb0000000000000010000000000000000000010000000000;
		10864: Delta = 46'sb1111111111111110000000000000000000010000000000;
		7749: Delta = 46'sb0000000000000001111111111111111111110000000000;
		8816: Delta = 46'sb1111111111111101111111111111111111110000000000;
		18570: Delta = 46'sb0000000000000100000000000000000000010000000000;
		2091: Delta = 46'sb1111111111111100000000000000000000010000000000;
		16522: Delta = 46'sb0000000000000011111111111111111111110000000000;
		43: Delta = 46'sb1111111111111011111111111111111111110000000000;
		17503: Delta = 46'sb0000000000001000000000000000000000010000000000;
		3158: Delta = 46'sb1111111111111000000000000000000000010000000000;
		15455: Delta = 46'sb0000000000000111111111111111111111110000000000;
		1110: Delta = 46'sb1111111111110111111111111111111111110000000000;
		15369: Delta = 46'sb0000000000010000000000000000000000010000000000;
		5292: Delta = 46'sb1111111111110000000000000000000000010000000000;
		13321: Delta = 46'sb0000000000001111111111111111111111110000000000;
		3244: Delta = 46'sb1111111111101111111111111111111111110000000000;
		11101: Delta = 46'sb0000000000100000000000000000000000010000000000;
		9560: Delta = 46'sb1111111111100000000000000000000000010000000000;
		9053: Delta = 46'sb0000000000011111111111111111111111110000000000;
		7512: Delta = 46'sb1111111111011111111111111111111111110000000000;
		2565: Delta = 46'sb0000000001000000000000000000000000010000000000;
		18096: Delta = 46'sb1111111111000000000000000000000000010000000000;
		517: Delta = 46'sb0000000000111111111111111111111111110000000000;
		16048: Delta = 46'sb1111111110111111111111111111111111110000000000;
		4106: Delta = 46'sb0000000010000000000000000000000000010000000000;
		16555: Delta = 46'sb1111111110000000000000000000000000010000000000;
		2058: Delta = 46'sb0000000001111111111111111111111111110000000000;
		14507: Delta = 46'sb1111111101111111111111111111111111110000000000;
		7188: Delta = 46'sb0000000100000000000000000000000000010000000000;
		13473: Delta = 46'sb1111111100000000000000000000000000010000000000;
		5140: Delta = 46'sb0000000011111111111111111111111111110000000000;
		11425: Delta = 46'sb1111111011111111111111111111111111110000000000;
		13352: Delta = 46'sb0000001000000000000000000000000000010000000000;
		7309: Delta = 46'sb1111111000000000000000000000000000010000000000;
		11304: Delta = 46'sb0000000111111111111111111111111111110000000000;
		5261: Delta = 46'sb1111110111111111111111111111111111110000000000;
		7067: Delta = 46'sb0000010000000000000000000000000000010000000000;
		13594: Delta = 46'sb1111110000000000000000000000000000010000000000;
		5019: Delta = 46'sb0000001111111111111111111111111111110000000000;
		11546: Delta = 46'sb1111101111111111111111111111111111110000000000;
		13110: Delta = 46'sb0000100000000000000000000000000000010000000000;
		7551: Delta = 46'sb1111100000000000000000000000000000010000000000;
		11062: Delta = 46'sb0000011111111111111111111111111111110000000000;
		5503: Delta = 46'sb1111011111111111111111111111111111110000000000;
		6583: Delta = 46'sb0001000000000000000000000000000000010000000000;
		14078: Delta = 46'sb1111000000000000000000000000000000010000000000;
		4535: Delta = 46'sb0000111111111111111111111111111111110000000000;
		12030: Delta = 46'sb1110111111111111111111111111111111110000000000;
		12142: Delta = 46'sb0010000000000000000000000000000000010000000000;
		8519: Delta = 46'sb1110000000000000000000000000000000010000000000;
		10094: Delta = 46'sb0001111111111111111111111111111111110000000000;
		6471: Delta = 46'sb1101111111111111111111111111111111110000000000;
		4647: Delta = 46'sb0100000000000000000000000000000000010000000000;
		16014: Delta = 46'sb1100000000000000000000000000000000010000000000;
		2599: Delta = 46'sb0011111111111111111111111111111111110000000000;
		13966: Delta = 46'sb1011111111111111111111111111111111110000000000;
		6144: Delta = 46'sb0000000000000000000000000000000001100000000000;
		12469: Delta = 46'sb1111111111111111111111111111111110100000000000;
		10240: Delta = 46'sb0000000000000000000000000000000010100000000000;
		8373: Delta = 46'sb1111111111111111111111111111111101100000000000;
		18432: Delta = 46'sb0000000000000000000000000000000100100000000000;
		4277: Delta = 46'sb1111111111111111111111111111111100100000000000;
		14336: Delta = 46'sb0000000000000000000000000000000011100000000000;
		181: Delta = 46'sb1111111111111111111111111111111011100000000000;
		16203: Delta = 46'sb0000000000000000000000000000001000100000000000;
		6506: Delta = 46'sb1111111111111111111111111111111000100000000000;
		12107: Delta = 46'sb0000000000000000000000000000000111100000000000;
		2410: Delta = 46'sb1111111111111111111111111111110111100000000000;
		11745: Delta = 46'sb0000000000000000000000000000010000100000000000;
		10964: Delta = 46'sb1111111111111111111111111111110000100000000000;
		7649: Delta = 46'sb0000000000000000000000000000001111100000000000;
		6868: Delta = 46'sb1111111111111111111111111111101111100000000000;
		2829: Delta = 46'sb0000000000000000000000000000100000100000000000;
		1267: Delta = 46'sb1111111111111111111111111111100000100000000000;
		17346: Delta = 46'sb0000000000000000000000000000011111100000000000;
		15784: Delta = 46'sb1111111111111111111111111111011111100000000000;
		3610: Delta = 46'sb0000000000000000000000000001000000100000000000;
		486: Delta = 46'sb1111111111111111111111111111000000100000000000;
		18127: Delta = 46'sb0000000000000000000000000000111111100000000000;
		15003: Delta = 46'sb1111111111111111111111111110111111100000000000;
		5172: Delta = 46'sb0000000000000000000000000010000000100000000000;
		17537: Delta = 46'sb1111111111111111111111111110000000100000000000;
		1076: Delta = 46'sb0000000000000000000000000001111111100000000000;
		13441: Delta = 46'sb1111111111111111111111111101111111100000000000;
		8296: Delta = 46'sb0000000000000000000000000100000000100000000000;
		14413: Delta = 46'sb1111111111111111111111111100000000100000000000;
		4200: Delta = 46'sb0000000000000000000000000011111111100000000000;
		10317: Delta = 46'sb1111111111111111111111111011111111100000000000;
		14544: Delta = 46'sb0000000000000000000000001000000000100000000000;
		8165: Delta = 46'sb1111111111111111111111111000000000100000000000;
		10448: Delta = 46'sb0000000000000000000000000111111111100000000000;
		4069: Delta = 46'sb1111111111111111111111110111111111100000000000;
		8427: Delta = 46'sb0000000000000000000000010000000000100000000000;
		14282: Delta = 46'sb1111111111111111111111110000000000100000000000;
		4331: Delta = 46'sb0000000000000000000000001111111111100000000000;
		10186: Delta = 46'sb1111111111111111111111101111111111100000000000;
		14806: Delta = 46'sb0000000000000000000000100000000000100000000000;
		7903: Delta = 46'sb1111111111111111111111100000000000100000000000;
		10710: Delta = 46'sb0000000000000000000000011111111111100000000000;
		3807: Delta = 46'sb1111111111111111111111011111111111100000000000;
		8951: Delta = 46'sb0000000000000000000001000000000000100000000000;
		13758: Delta = 46'sb1111111111111111111111000000000000100000000000;
		4855: Delta = 46'sb0000000000000000000000111111111111100000000000;
		9662: Delta = 46'sb1111111111111111111110111111111111100000000000;
		15854: Delta = 46'sb0000000000000000000010000000000000100000000000;
		6855: Delta = 46'sb1111111111111111111110000000000000100000000000;
		11758: Delta = 46'sb0000000000000000000001111111111111100000000000;
		2759: Delta = 46'sb1111111111111111111101111111111111100000000000;
		11047: Delta = 46'sb0000000000000000000100000000000000100000000000;
		11662: Delta = 46'sb1111111111111111111100000000000000100000000000;
		6951: Delta = 46'sb0000000000000000000011111111111111100000000000;
		7566: Delta = 46'sb1111111111111111111011111111111111100000000000;
		1433: Delta = 46'sb0000000000000000001000000000000000100000000000;
		2663: Delta = 46'sb1111111111111111111000000000000000100000000000;
		15950: Delta = 46'sb0000000000000000000111111111111111100000000000;
		17180: Delta = 46'sb1111111111111111110111111111111111100000000000;
		818: Delta = 46'sb0000000000000000010000000000000000100000000000;
		3278: Delta = 46'sb1111111111111111110000000000000000100000000000;
		15335: Delta = 46'sb0000000000000000001111111111111111100000000000;
		17795: Delta = 46'sb1111111111111111101111111111111111100000000000;
		18201: Delta = 46'sb0000000000000000100000000000000000100000000000;
		4508: Delta = 46'sb1111111111111111100000000000000000100000000000;
		14105: Delta = 46'sb0000000000000000011111111111111111100000000000;
		412: Delta = 46'sb1111111111111111011111111111111111100000000000;
		15741: Delta = 46'sb0000000000000001000000000000000000100000000000;
		6968: Delta = 46'sb1111111111111111000000000000000000100000000000;
		11645: Delta = 46'sb0000000000000000111111111111111111100000000000;
		2872: Delta = 46'sb1111111111111110111111111111111111100000000000;
		10821: Delta = 46'sb0000000000000010000000000000000000100000000000;
		11888: Delta = 46'sb1111111111111110000000000000000000100000000000;
		6725: Delta = 46'sb0000000000000001111111111111111111100000000000;
		7792: Delta = 46'sb1111111111111101111111111111111111100000000000;
		981: Delta = 46'sb0000000000000100000000000000000000100000000000;
		3115: Delta = 46'sb1111111111111100000000000000000000100000000000;
		15498: Delta = 46'sb0000000000000011111111111111111111100000000000;
		17632: Delta = 46'sb1111111111111011111111111111111111100000000000;
		18527: Delta = 46'sb0000000000001000000000000000000000100000000000;
		4182: Delta = 46'sb1111111111111000000000000000000000100000000000;
		14431: Delta = 46'sb0000000000000111111111111111111111100000000000;
		86: Delta = 46'sb1111111111110111111111111111111111100000000000;
		16393: Delta = 46'sb0000000000010000000000000000000000100000000000;
		6316: Delta = 46'sb1111111111110000000000000000000000100000000000;
		12297: Delta = 46'sb0000000000001111111111111111111111100000000000;
		2220: Delta = 46'sb1111111111101111111111111111111111100000000000;
		12125: Delta = 46'sb0000000000100000000000000000000000100000000000;
		10584: Delta = 46'sb1111111111100000000000000000000000100000000000;
		8029: Delta = 46'sb0000000000011111111111111111111111100000000000;
		6488: Delta = 46'sb1111111111011111111111111111111111100000000000;
		3589: Delta = 46'sb0000000001000000000000000000000000100000000000;
		507: Delta = 46'sb1111111111000000000000000000000000100000000000;
		18106: Delta = 46'sb0000000000111111111111111111111111100000000000;
		15024: Delta = 46'sb1111111110111111111111111111111111100000000000;
		5130: Delta = 46'sb0000000010000000000000000000000000100000000000;
		17579: Delta = 46'sb1111111110000000000000000000000000100000000000;
		1034: Delta = 46'sb0000000001111111111111111111111111100000000000;
		13483: Delta = 46'sb1111111101111111111111111111111111100000000000;
		8212: Delta = 46'sb0000000100000000000000000000000000100000000000;
		14497: Delta = 46'sb1111111100000000000000000000000000100000000000;
		4116: Delta = 46'sb0000000011111111111111111111111111100000000000;
		10401: Delta = 46'sb1111111011111111111111111111111111100000000000;
		14376: Delta = 46'sb0000001000000000000000000000000000100000000000;
		8333: Delta = 46'sb1111111000000000000000000000000000100000000000;
		10280: Delta = 46'sb0000000111111111111111111111111111100000000000;
		4237: Delta = 46'sb1111110111111111111111111111111111100000000000;
		8091: Delta = 46'sb0000010000000000000000000000000000100000000000;
		14618: Delta = 46'sb1111110000000000000000000000000000100000000000;
		3995: Delta = 46'sb0000001111111111111111111111111111100000000000;
		10522: Delta = 46'sb1111101111111111111111111111111111100000000000;
		14134: Delta = 46'sb0000100000000000000000000000000000100000000000;
		8575: Delta = 46'sb1111100000000000000000000000000000100000000000;
		10038: Delta = 46'sb0000011111111111111111111111111111100000000000;
		4479: Delta = 46'sb1111011111111111111111111111111111100000000000;
		7607: Delta = 46'sb0001000000000000000000000000000000100000000000;
		15102: Delta = 46'sb1111000000000000000000000000000000100000000000;
		3511: Delta = 46'sb0000111111111111111111111111111111100000000000;
		11006: Delta = 46'sb1110111111111111111111111111111111100000000000;
		13166: Delta = 46'sb0010000000000000000000000000000000100000000000;
		9543: Delta = 46'sb1110000000000000000000000000000000100000000000;
		9070: Delta = 46'sb0001111111111111111111111111111111100000000000;
		5447: Delta = 46'sb1101111111111111111111111111111111100000000000;
		5671: Delta = 46'sb0100000000000000000000000000000000100000000000;
		17038: Delta = 46'sb1100000000000000000000000000000000100000000000;
		1575: Delta = 46'sb0011111111111111111111111111111111100000000000;
		12942: Delta = 46'sb1011111111111111111111111111111111100000000000;
		12288: Delta = 46'sb0000000000000000000000000000000011000000000000;
		6325: Delta = 46'sb1111111111111111111111111111111101000000000000;
		1867: Delta = 46'sb0000000000000000000000000000000101000000000000;
		16746: Delta = 46'sb1111111111111111111111111111111011000000000000;
		18251: Delta = 46'sb0000000000000000000000000000001001000000000000;
		8554: Delta = 46'sb1111111111111111111111111111111001000000000000;
		10059: Delta = 46'sb0000000000000000000000000000000111000000000000;
		362: Delta = 46'sb1111111111111111111111111111110111000000000000;
		13793: Delta = 46'sb0000000000000000000000000000010001000000000000;
		13012: Delta = 46'sb1111111111111111111111111111110001000000000000;
		5601: Delta = 46'sb0000000000000000000000000000001111000000000000;
		4820: Delta = 46'sb1111111111111111111111111111101111000000000000;
		4877: Delta = 46'sb0000000000000000000000000000100001000000000000;
		3315: Delta = 46'sb1111111111111111111111111111100001000000000000;
		15298: Delta = 46'sb0000000000000000000000000000011111000000000000;
		13736: Delta = 46'sb1111111111111111111111111111011111000000000000;
		5658: Delta = 46'sb0000000000000000000000000001000001000000000000;
		2534: Delta = 46'sb1111111111111111111111111111000001000000000000;
		16079: Delta = 46'sb0000000000000000000000000000111111000000000000;
		12955: Delta = 46'sb1111111111111111111111111110111111000000000000;
		7220: Delta = 46'sb0000000000000000000000000010000001000000000000;
		972: Delta = 46'sb1111111111111111111111111110000001000000000000;
		17641: Delta = 46'sb0000000000000000000000000001111111000000000000;
		11393: Delta = 46'sb1111111111111111111111111101111111000000000000;
		10344: Delta = 46'sb0000000000000000000000000100000001000000000000;
		16461: Delta = 46'sb1111111111111111111111111100000001000000000000;
		2152: Delta = 46'sb0000000000000000000000000011111111000000000000;
		8269: Delta = 46'sb1111111111111111111111111011111111000000000000;
		16592: Delta = 46'sb0000000000000000000000001000000001000000000000;
		10213: Delta = 46'sb1111111111111111111111111000000001000000000000;
		8400: Delta = 46'sb0000000000000000000000000111111111000000000000;
		2021: Delta = 46'sb1111111111111111111111110111111111000000000000;
		10475: Delta = 46'sb0000000000000000000000010000000001000000000000;
		16330: Delta = 46'sb1111111111111111111111110000000001000000000000;
		2283: Delta = 46'sb0000000000000000000000001111111111000000000000;
		8138: Delta = 46'sb1111111111111111111111101111111111000000000000;
		16854: Delta = 46'sb0000000000000000000000100000000001000000000000;
		9951: Delta = 46'sb1111111111111111111111100000000001000000000000;
		8662: Delta = 46'sb0000000000000000000000011111111111000000000000;
		1759: Delta = 46'sb1111111111111111111111011111111111000000000000;
		10999: Delta = 46'sb0000000000000000000001000000000001000000000000;
		15806: Delta = 46'sb1111111111111111111111000000000001000000000000;
		2807: Delta = 46'sb0000000000000000000000111111111111000000000000;
		7614: Delta = 46'sb1111111111111111111110111111111111000000000000;
		17902: Delta = 46'sb0000000000000000000010000000000001000000000000;
		8903: Delta = 46'sb1111111111111111111110000000000001000000000000;
		9710: Delta = 46'sb0000000000000000000001111111111111000000000000;
		711: Delta = 46'sb1111111111111111111101111111111111000000000000;
		13095: Delta = 46'sb0000000000000000000100000000000001000000000000;
		13710: Delta = 46'sb1111111111111111111100000000000001000000000000;
		4903: Delta = 46'sb0000000000000000000011111111111111000000000000;
		5518: Delta = 46'sb1111111111111111111011111111111111000000000000;
		3481: Delta = 46'sb0000000000000000001000000000000001000000000000;
		4711: Delta = 46'sb1111111111111111111000000000000001000000000000;
		13902: Delta = 46'sb0000000000000000000111111111111111000000000000;
		15132: Delta = 46'sb1111111111111111110111111111111111000000000000;
		2866: Delta = 46'sb0000000000000000010000000000000001000000000000;
		5326: Delta = 46'sb1111111111111111110000000000000001000000000000;
		13287: Delta = 46'sb0000000000000000001111111111111111000000000000;
		15747: Delta = 46'sb1111111111111111101111111111111111000000000000;
		1636: Delta = 46'sb0000000000000000100000000000000001000000000000;
		6556: Delta = 46'sb1111111111111111100000000000000001000000000000;
		12057: Delta = 46'sb0000000000000000011111111111111111000000000000;
		16977: Delta = 46'sb1111111111111111011111111111111111000000000000;
		17789: Delta = 46'sb0000000000000001000000000000000001000000000000;
		9016: Delta = 46'sb1111111111111111000000000000000001000000000000;
		9597: Delta = 46'sb0000000000000000111111111111111111000000000000;
		824: Delta = 46'sb1111111111111110111111111111111111000000000000;
		12869: Delta = 46'sb0000000000000010000000000000000001000000000000;
		13936: Delta = 46'sb1111111111111110000000000000000001000000000000;
		4677: Delta = 46'sb0000000000000001111111111111111111000000000000;
		5744: Delta = 46'sb1111111111111101111111111111111111000000000000;
		3029: Delta = 46'sb0000000000000100000000000000000001000000000000;
		5163: Delta = 46'sb1111111111111100000000000000000001000000000000;
		13450: Delta = 46'sb0000000000000011111111111111111111000000000000;
		15584: Delta = 46'sb1111111111111011111111111111111111000000000000;
		1962: Delta = 46'sb0000000000001000000000000000000001000000000000;
		6230: Delta = 46'sb1111111111111000000000000000000001000000000000;
		12383: Delta = 46'sb0000000000000111111111111111111111000000000000;
		16651: Delta = 46'sb1111111111110111111111111111111111000000000000;
		18441: Delta = 46'sb0000000000010000000000000000000001000000000000;
		8364: Delta = 46'sb1111111111110000000000000000000001000000000000;
		10249: Delta = 46'sb0000000000001111111111111111111111000000000000;
		172: Delta = 46'sb1111111111101111111111111111111111000000000000;
		14173: Delta = 46'sb0000000000100000000000000000000001000000000000;
		12632: Delta = 46'sb1111111111100000000000000000000001000000000000;
		5981: Delta = 46'sb0000000000011111111111111111111111000000000000;
		4440: Delta = 46'sb1111111111011111111111111111111111000000000000;
		5637: Delta = 46'sb0000000001000000000000000000000001000000000000;
		2555: Delta = 46'sb1111111111000000000000000000000001000000000000;
		16058: Delta = 46'sb0000000000111111111111111111111111000000000000;
		12976: Delta = 46'sb1111111110111111111111111111111111000000000000;
		7178: Delta = 46'sb0000000010000000000000000000000001000000000000;
		1014: Delta = 46'sb1111111110000000000000000000000001000000000000;
		17599: Delta = 46'sb0000000001111111111111111111111111000000000000;
		11435: Delta = 46'sb1111111101111111111111111111111111000000000000;
		10260: Delta = 46'sb0000000100000000000000000000000001000000000000;
		16545: Delta = 46'sb1111111100000000000000000000000001000000000000;
		2068: Delta = 46'sb0000000011111111111111111111111111000000000000;
		8353: Delta = 46'sb1111111011111111111111111111111111000000000000;
		16424: Delta = 46'sb0000001000000000000000000000000001000000000000;
		10381: Delta = 46'sb1111111000000000000000000000000001000000000000;
		8232: Delta = 46'sb0000000111111111111111111111111111000000000000;
		2189: Delta = 46'sb1111110111111111111111111111111111000000000000;
		10139: Delta = 46'sb0000010000000000000000000000000001000000000000;
		16666: Delta = 46'sb1111110000000000000000000000000001000000000000;
		1947: Delta = 46'sb0000001111111111111111111111111111000000000000;
		8474: Delta = 46'sb1111101111111111111111111111111111000000000000;
		16182: Delta = 46'sb0000100000000000000000000000000001000000000000;
		10623: Delta = 46'sb1111100000000000000000000000000001000000000000;
		7990: Delta = 46'sb0000011111111111111111111111111111000000000000;
		2431: Delta = 46'sb1111011111111111111111111111111111000000000000;
		9655: Delta = 46'sb0001000000000000000000000000000001000000000000;
		17150: Delta = 46'sb1111000000000000000000000000000001000000000000;
		1463: Delta = 46'sb0000111111111111111111111111111111000000000000;
		8958: Delta = 46'sb1110111111111111111111111111111111000000000000;
		15214: Delta = 46'sb0010000000000000000000000000000001000000000000;
		11591: Delta = 46'sb1110000000000000000000000000000001000000000000;
		7022: Delta = 46'sb0001111111111111111111111111111111000000000000;
		3399: Delta = 46'sb1101111111111111111111111111111111000000000000;
		7719: Delta = 46'sb0100000000000000000000000000000001000000000000;
		473: Delta = 46'sb1100000000000000000000000000000001000000000000;
		18140: Delta = 46'sb0011111111111111111111111111111111000000000000;
		10894: Delta = 46'sb1011111111111111111111111111111111000000000000;
		5963: Delta = 46'sb0000000000000000000000000000000110000000000000;
		12650: Delta = 46'sb1111111111111111111111111111111010000000000000;
		3734: Delta = 46'sb0000000000000000000000000000001010000000000000;
		14879: Delta = 46'sb1111111111111111111111111111110110000000000000;
		17889: Delta = 46'sb0000000000000000000000000000010010000000000000;
		17108: Delta = 46'sb1111111111111111111111111111110010000000000000;
		1505: Delta = 46'sb0000000000000000000000000000001110000000000000;
		724: Delta = 46'sb1111111111111111111111111111101110000000000000;
		8973: Delta = 46'sb0000000000000000000000000000100010000000000000;
		7411: Delta = 46'sb1111111111111111111111111111100010000000000000;
		11202: Delta = 46'sb0000000000000000000000000000011110000000000000;
		9640: Delta = 46'sb1111111111111111111111111111011110000000000000;
		9754: Delta = 46'sb0000000000000000000000000001000010000000000000;
		6630: Delta = 46'sb1111111111111111111111111111000010000000000000;
		11983: Delta = 46'sb0000000000000000000000000000111110000000000000;
		8859: Delta = 46'sb1111111111111111111111111110111110000000000000;
		11316: Delta = 46'sb0000000000000000000000000010000010000000000000;
		5068: Delta = 46'sb1111111111111111111111111110000010000000000000;
		13545: Delta = 46'sb0000000000000000000000000001111110000000000000;
		7297: Delta = 46'sb1111111111111111111111111101111110000000000000;
		14440: Delta = 46'sb0000000000000000000000000100000010000000000000;
		1944: Delta = 46'sb1111111111111111111111111100000010000000000000;
		16669: Delta = 46'sb0000000000000000000000000011111110000000000000;
		4173: Delta = 46'sb1111111111111111111111111011111110000000000000;
		2075: Delta = 46'sb0000000000000000000000001000000010000000000000;
		14309: Delta = 46'sb1111111111111111111111111000000010000000000000;
		4304: Delta = 46'sb0000000000000000000000000111111110000000000000;
		16538: Delta = 46'sb1111111111111111111111110111111110000000000000;
		14571: Delta = 46'sb0000000000000000000000010000000010000000000000;
		1813: Delta = 46'sb1111111111111111111111110000000010000000000000;
		16800: Delta = 46'sb0000000000000000000000001111111110000000000000;
		4042: Delta = 46'sb1111111111111111111111101111111110000000000000;
		2337: Delta = 46'sb0000000000000000000000100000000010000000000000;
		14047: Delta = 46'sb1111111111111111111111100000000010000000000000;
		4566: Delta = 46'sb0000000000000000000000011111111110000000000000;
		16276: Delta = 46'sb1111111111111111111111011111111110000000000000;
		15095: Delta = 46'sb0000000000000000000001000000000010000000000000;
		1289: Delta = 46'sb1111111111111111111111000000000010000000000000;
		17324: Delta = 46'sb0000000000000000000000111111111110000000000000;
		3518: Delta = 46'sb1111111111111111111110111111111110000000000000;
		3385: Delta = 46'sb0000000000000000000010000000000010000000000000;
		12999: Delta = 46'sb1111111111111111111110000000000010000000000000;
		5614: Delta = 46'sb0000000000000000000001111111111110000000000000;
		15228: Delta = 46'sb1111111111111111111101111111111110000000000000;
		17191: Delta = 46'sb0000000000000000000100000000000010000000000000;
		17806: Delta = 46'sb1111111111111111111100000000000010000000000000;
		807: Delta = 46'sb0000000000000000000011111111111110000000000000;
		1422: Delta = 46'sb1111111111111111111011111111111110000000000000;
		7577: Delta = 46'sb0000000000000000001000000000000010000000000000;
		8807: Delta = 46'sb1111111111111111111000000000000010000000000000;
		9806: Delta = 46'sb0000000000000000000111111111111110000000000000;
		11036: Delta = 46'sb1111111111111111110111111111111110000000000000;
		6962: Delta = 46'sb0000000000000000010000000000000010000000000000;
		9422: Delta = 46'sb1111111111111111110000000000000010000000000000;
		9191: Delta = 46'sb0000000000000000001111111111111110000000000000;
		11651: Delta = 46'sb1111111111111111101111111111111110000000000000;
		5732: Delta = 46'sb0000000000000000100000000000000010000000000000;
		10652: Delta = 46'sb1111111111111111100000000000000010000000000000;
		7961: Delta = 46'sb0000000000000000011111111111111110000000000000;
		12881: Delta = 46'sb1111111111111111011111111111111110000000000000;
		3272: Delta = 46'sb0000000000000001000000000000000010000000000000;
		13112: Delta = 46'sb1111111111111111000000000000000010000000000000;
		5501: Delta = 46'sb0000000000000000111111111111111110000000000000;
		15341: Delta = 46'sb1111111111111110111111111111111110000000000000;
		16965: Delta = 46'sb0000000000000010000000000000000010000000000000;
		18032: Delta = 46'sb1111111111111110000000000000000010000000000000;
		581: Delta = 46'sb0000000000000001111111111111111110000000000000;
		1648: Delta = 46'sb1111111111111101111111111111111110000000000000;
		7125: Delta = 46'sb0000000000000100000000000000000010000000000000;
		9259: Delta = 46'sb1111111111111100000000000000000010000000000000;
		9354: Delta = 46'sb0000000000000011111111111111111110000000000000;
		11488: Delta = 46'sb1111111111111011111111111111111110000000000000;
		6058: Delta = 46'sb0000000000001000000000000000000010000000000000;
		10326: Delta = 46'sb1111111111111000000000000000000010000000000000;
		8287: Delta = 46'sb0000000000000111111111111111111110000000000000;
		12555: Delta = 46'sb1111111111110111111111111111111110000000000000;
		3924: Delta = 46'sb0000000000010000000000000000000010000000000000;
		12460: Delta = 46'sb1111111111110000000000000000000010000000000000;
		6153: Delta = 46'sb0000000000001111111111111111111110000000000000;
		14689: Delta = 46'sb1111111111101111111111111111111110000000000000;
		18269: Delta = 46'sb0000000000100000000000000000000010000000000000;
		16728: Delta = 46'sb1111111111100000000000000000000010000000000000;
		1885: Delta = 46'sb0000000000011111111111111111111110000000000000;
		344: Delta = 46'sb1111111111011111111111111111111110000000000000;
		9733: Delta = 46'sb0000000001000000000000000000000010000000000000;
		6651: Delta = 46'sb1111111111000000000000000000000010000000000000;
		11962: Delta = 46'sb0000000000111111111111111111111110000000000000;
		8880: Delta = 46'sb1111111110111111111111111111111110000000000000;
		11274: Delta = 46'sb0000000010000000000000000000000010000000000000;
		5110: Delta = 46'sb1111111110000000000000000000000010000000000000;
		13503: Delta = 46'sb0000000001111111111111111111111110000000000000;
		7339: Delta = 46'sb1111111101111111111111111111111110000000000000;
		14356: Delta = 46'sb0000000100000000000000000000000010000000000000;
		2028: Delta = 46'sb1111111100000000000000000000000010000000000000;
		16585: Delta = 46'sb0000000011111111111111111111111110000000000000;
		4257: Delta = 46'sb1111111011111111111111111111111110000000000000;
		1907: Delta = 46'sb0000001000000000000000000000000010000000000000;
		14477: Delta = 46'sb1111111000000000000000000000000010000000000000;
		4136: Delta = 46'sb0000000111111111111111111111111110000000000000;
		16706: Delta = 46'sb1111110111111111111111111111111110000000000000;
		14235: Delta = 46'sb0000010000000000000000000000000010000000000000;
		2149: Delta = 46'sb1111110000000000000000000000000010000000000000;
		16464: Delta = 46'sb0000001111111111111111111111111110000000000000;
		4378: Delta = 46'sb1111101111111111111111111111111110000000000000;
		1665: Delta = 46'sb0000100000000000000000000000000010000000000000;
		14719: Delta = 46'sb1111100000000000000000000000000010000000000000;
		3894: Delta = 46'sb0000011111111111111111111111111110000000000000;
		16948: Delta = 46'sb1111011111111111111111111111111110000000000000;
		13751: Delta = 46'sb0001000000000000000000000000000010000000000000;
		2633: Delta = 46'sb1111000000000000000000000000000010000000000000;
		15980: Delta = 46'sb0000111111111111111111111111111110000000000000;
		4862: Delta = 46'sb1110111111111111111111111111111110000000000000;
		697: Delta = 46'sb0010000000000000000000000000000010000000000000;
		15687: Delta = 46'sb1110000000000000000000000000000010000000000000;
		2926: Delta = 46'sb0001111111111111111111111111111110000000000000;
		17916: Delta = 46'sb1101111111111111111111111111111110000000000000;
		11815: Delta = 46'sb0100000000000000000000000000000010000000000000;
		4569: Delta = 46'sb1100000000000000000000000000000010000000000000;
		14044: Delta = 46'sb0011111111111111111111111111111110000000000000;
		6798: Delta = 46'sb1011111111111111111111111111111110000000000000;
		11926: Delta = 46'sb0000000000000000000000000000001100000000000000;
		6687: Delta = 46'sb1111111111111111111111111111110100000000000000;
		7468: Delta = 46'sb0000000000000000000000000000010100000000000000;
		11145: Delta = 46'sb1111111111111111111111111111101100000000000000;
		17165: Delta = 46'sb0000000000000000000000000000100100000000000000;
		15603: Delta = 46'sb1111111111111111111111111111100100000000000000;
		3010: Delta = 46'sb0000000000000000000000000000011100000000000000;
		1448: Delta = 46'sb1111111111111111111111111111011100000000000000;
		17946: Delta = 46'sb0000000000000000000000000001000100000000000000;
		14822: Delta = 46'sb1111111111111111111111111111000100000000000000;
		3791: Delta = 46'sb0000000000000000000000000000111100000000000000;
		667: Delta = 46'sb1111111111111111111111111110111100000000000000;
		895: Delta = 46'sb0000000000000000000000000010000100000000000000;
		13260: Delta = 46'sb1111111111111111111111111110000100000000000000;
		5353: Delta = 46'sb0000000000000000000000000001111100000000000000;
		17718: Delta = 46'sb1111111111111111111111111101111100000000000000;
		4019: Delta = 46'sb0000000000000000000000000100000100000000000000;
		10136: Delta = 46'sb1111111111111111111111111100000100000000000000;
		8477: Delta = 46'sb0000000000000000000000000011111100000000000000;
		14594: Delta = 46'sb1111111111111111111111111011111100000000000000;
		10267: Delta = 46'sb0000000000000000000000001000000100000000000000;
		3888: Delta = 46'sb1111111111111111111111111000000100000000000000;
		14725: Delta = 46'sb0000000000000000000000000111111100000000000000;
		8346: Delta = 46'sb1111111111111111111111110111111100000000000000;
		4150: Delta = 46'sb0000000000000000000000010000000100000000000000;
		10005: Delta = 46'sb1111111111111111111111110000000100000000000000;
		8608: Delta = 46'sb0000000000000000000000001111111100000000000000;
		14463: Delta = 46'sb1111111111111111111111101111111100000000000000;
		10529: Delta = 46'sb0000000000000000000000100000000100000000000000;
		3626: Delta = 46'sb1111111111111111111111100000000100000000000000;
		14987: Delta = 46'sb0000000000000000000000011111111100000000000000;
		8084: Delta = 46'sb1111111111111111111111011111111100000000000000;
		4674: Delta = 46'sb0000000000000000000001000000000100000000000000;
		9481: Delta = 46'sb1111111111111111111111000000000100000000000000;
		9132: Delta = 46'sb0000000000000000000000111111111100000000000000;
		13939: Delta = 46'sb1111111111111111111110111111111100000000000000;
		11577: Delta = 46'sb0000000000000000000010000000000100000000000000;
		2578: Delta = 46'sb1111111111111111111110000000000100000000000000;
		16035: Delta = 46'sb0000000000000000000001111111111100000000000000;
		7036: Delta = 46'sb1111111111111111111101111111111100000000000000;
		6770: Delta = 46'sb0000000000000000000100000000000100000000000000;
		7385: Delta = 46'sb1111111111111111111100000000000100000000000000;
		11228: Delta = 46'sb0000000000000000000011111111111100000000000000;
		11843: Delta = 46'sb1111111111111111111011111111111100000000000000;
		15769: Delta = 46'sb0000000000000000001000000000000100000000000000;
		16999: Delta = 46'sb1111111111111111111000000000000100000000000000;
		1614: Delta = 46'sb0000000000000000000111111111111100000000000000;
		2844: Delta = 46'sb1111111111111111110111111111111100000000000000;
		15154: Delta = 46'sb0000000000000000010000000000000100000000000000;
		17614: Delta = 46'sb1111111111111111110000000000000100000000000000;
		999: Delta = 46'sb0000000000000000001111111111111100000000000000;
		3459: Delta = 46'sb1111111111111111101111111111111100000000000000;
		13924: Delta = 46'sb0000000000000000100000000000000100000000000000;
		231: Delta = 46'sb1111111111111111100000000000000100000000000000;
		18382: Delta = 46'sb0000000000000000011111111111111100000000000000;
		4689: Delta = 46'sb1111111111111111011111111111111100000000000000;
		11464: Delta = 46'sb0000000000000001000000000000000100000000000000;
		2691: Delta = 46'sb1111111111111111000000000000000100000000000000;
		15922: Delta = 46'sb0000000000000000111111111111111100000000000000;
		7149: Delta = 46'sb1111111111111110111111111111111100000000000000;
		6544: Delta = 46'sb0000000000000010000000000000000100000000000000;
		7611: Delta = 46'sb1111111111111110000000000000000100000000000000;
		11002: Delta = 46'sb0000000000000001111111111111111100000000000000;
		12069: Delta = 46'sb1111111111111101111111111111111100000000000000;
		15317: Delta = 46'sb0000000000000100000000000000000100000000000000;
		17451: Delta = 46'sb1111111111111100000000000000000100000000000000;
		1162: Delta = 46'sb0000000000000011111111111111111100000000000000;
		3296: Delta = 46'sb1111111111111011111111111111111100000000000000;
		14250: Delta = 46'sb0000000000001000000000000000000100000000000000;
		18518: Delta = 46'sb1111111111111000000000000000000100000000000000;
		95: Delta = 46'sb0000000000000111111111111111111100000000000000;
		4363: Delta = 46'sb1111111111110111111111111111111100000000000000;
		12116: Delta = 46'sb0000000000010000000000000000000100000000000000;
		2039: Delta = 46'sb1111111111110000000000000000000100000000000000;
		16574: Delta = 46'sb0000000000001111111111111111111100000000000000;
		6497: Delta = 46'sb1111111111101111111111111111111100000000000000;
		7848: Delta = 46'sb0000000000100000000000000000000100000000000000;
		6307: Delta = 46'sb1111111111100000000000000000000100000000000000;
		12306: Delta = 46'sb0000000000011111111111111111111100000000000000;
		10765: Delta = 46'sb1111111111011111111111111111111100000000000000;
		17925: Delta = 46'sb0000000001000000000000000000000100000000000000;
		14843: Delta = 46'sb1111111111000000000000000000000100000000000000;
		3770: Delta = 46'sb0000000000111111111111111111111100000000000000;
		688: Delta = 46'sb1111111110111111111111111111111100000000000000;
		853: Delta = 46'sb0000000010000000000000000000000100000000000000;
		13302: Delta = 46'sb1111111110000000000000000000000100000000000000;
		5311: Delta = 46'sb0000000001111111111111111111111100000000000000;
		17760: Delta = 46'sb1111111101111111111111111111111100000000000000;
		3935: Delta = 46'sb0000000100000000000000000000000100000000000000;
		10220: Delta = 46'sb1111111100000000000000000000000100000000000000;
		8393: Delta = 46'sb0000000011111111111111111111111100000000000000;
		14678: Delta = 46'sb1111111011111111111111111111111100000000000000;
		10099: Delta = 46'sb0000001000000000000000000000000100000000000000;
		4056: Delta = 46'sb1111111000000000000000000000000100000000000000;
		14557: Delta = 46'sb0000000111111111111111111111111100000000000000;
		8514: Delta = 46'sb1111110111111111111111111111111100000000000000;
		3814: Delta = 46'sb0000010000000000000000000000000100000000000000;
		10341: Delta = 46'sb1111110000000000000000000000000100000000000000;
		8272: Delta = 46'sb0000001111111111111111111111111100000000000000;
		14799: Delta = 46'sb1111101111111111111111111111111100000000000000;
		9857: Delta = 46'sb0000100000000000000000000000000100000000000000;
		4298: Delta = 46'sb1111100000000000000000000000000100000000000000;
		14315: Delta = 46'sb0000011111111111111111111111111100000000000000;
		8756: Delta = 46'sb1111011111111111111111111111111100000000000000;
		3330: Delta = 46'sb0001000000000000000000000000000100000000000000;
		10825: Delta = 46'sb1111000000000000000000000000000100000000000000;
		7788: Delta = 46'sb0000111111111111111111111111111100000000000000;
		15283: Delta = 46'sb1110111111111111111111111111111100000000000000;
		8889: Delta = 46'sb0010000000000000000000000000000100000000000000;
		5266: Delta = 46'sb1110000000000000000000000000000100000000000000;
		13347: Delta = 46'sb0001111111111111111111111111111100000000000000;
		9724: Delta = 46'sb1101111111111111111111111111111100000000000000;
		1394: Delta = 46'sb0100000000000000000000000000000100000000000000;
		12761: Delta = 46'sb1100000000000000000000000000000100000000000000;
		5852: Delta = 46'sb0011111111111111111111111111111100000000000000;
		17219: Delta = 46'sb1011111111111111111111111111111100000000000000;
		5239: Delta = 46'sb0000000000000000000000000000011000000000000000;
		13374: Delta = 46'sb1111111111111111111111111111101000000000000000;
		14936: Delta = 46'sb0000000000000000000000000000101000000000000000;
		3677: Delta = 46'sb1111111111111111111111111111011000000000000000;
		15717: Delta = 46'sb0000000000000000000000000001001000000000000000;
		12593: Delta = 46'sb1111111111111111111111111111001000000000000000;
		6020: Delta = 46'sb0000000000000000000000000000111000000000000000;
		2896: Delta = 46'sb1111111111111111111111111110111000000000000000;
		17279: Delta = 46'sb0000000000000000000000000010001000000000000000;
		11031: Delta = 46'sb1111111111111111111111111110001000000000000000;
		7582: Delta = 46'sb0000000000000000000000000001111000000000000000;
		1334: Delta = 46'sb1111111111111111111111111101111000000000000000;
		1790: Delta = 46'sb0000000000000000000000000100001000000000000000;
		7907: Delta = 46'sb1111111111111111111111111100001000000000000000;
		10706: Delta = 46'sb0000000000000000000000000011111000000000000000;
		16823: Delta = 46'sb1111111111111111111111111011111000000000000000;
		8038: Delta = 46'sb0000000000000000000000001000001000000000000000;
		1659: Delta = 46'sb1111111111111111111111111000001000000000000000;
		16954: Delta = 46'sb0000000000000000000000000111111000000000000000;
		10575: Delta = 46'sb1111111111111111111111110111111000000000000000;
		1921: Delta = 46'sb0000000000000000000000010000001000000000000000;
		7776: Delta = 46'sb1111111111111111111111110000001000000000000000;
		10837: Delta = 46'sb0000000000000000000000001111111000000000000000;
		16692: Delta = 46'sb1111111111111111111111101111111000000000000000;
		8300: Delta = 46'sb0000000000000000000000100000001000000000000000;
		1397: Delta = 46'sb1111111111111111111111100000001000000000000000;
		17216: Delta = 46'sb0000000000000000000000011111111000000000000000;
		10313: Delta = 46'sb1111111111111111111111011111111000000000000000;
		2445: Delta = 46'sb0000000000000000000001000000001000000000000000;
		7252: Delta = 46'sb1111111111111111111111000000001000000000000000;
		11361: Delta = 46'sb0000000000000000000000111111111000000000000000;
		16168: Delta = 46'sb1111111111111111111110111111111000000000000000;
		9348: Delta = 46'sb0000000000000000000010000000001000000000000000;
		349: Delta = 46'sb1111111111111111111110000000001000000000000000;
		18264: Delta = 46'sb0000000000000000000001111111111000000000000000;
		9265: Delta = 46'sb1111111111111111111101111111111000000000000000;
		4541: Delta = 46'sb0000000000000000000100000000001000000000000000;
		5156: Delta = 46'sb1111111111111111111100000000001000000000000000;
		13457: Delta = 46'sb0000000000000000000011111111111000000000000000;
		14072: Delta = 46'sb1111111111111111111011111111111000000000000000;
		13540: Delta = 46'sb0000000000000000001000000000001000000000000000;
		14770: Delta = 46'sb1111111111111111111000000000001000000000000000;
		3843: Delta = 46'sb0000000000000000000111111111111000000000000000;
		5073: Delta = 46'sb1111111111111111110111111111111000000000000000;
		12925: Delta = 46'sb0000000000000000010000000000001000000000000000;
		15385: Delta = 46'sb1111111111111111110000000000001000000000000000;
		3228: Delta = 46'sb0000000000000000001111111111111000000000000000;
		5688: Delta = 46'sb1111111111111111101111111111111000000000000000;
		11695: Delta = 46'sb0000000000000000100000000000001000000000000000;
		16615: Delta = 46'sb1111111111111111100000000000001000000000000000;
		1998: Delta = 46'sb0000000000000000011111111111111000000000000000;
		6918: Delta = 46'sb1111111111111111011111111111111000000000000000;
		9235: Delta = 46'sb0000000000000001000000000000001000000000000000;
		462: Delta = 46'sb1111111111111111000000000000001000000000000000;
		18151: Delta = 46'sb0000000000000000111111111111111000000000000000;
		9378: Delta = 46'sb1111111111111110111111111111111000000000000000;
		4315: Delta = 46'sb0000000000000010000000000000001000000000000000;
		5382: Delta = 46'sb1111111111111110000000000000001000000000000000;
		13231: Delta = 46'sb0000000000000001111111111111111000000000000000;
		14298: Delta = 46'sb1111111111111101111111111111111000000000000000;
		13088: Delta = 46'sb0000000000000100000000000000001000000000000000;
		15222: Delta = 46'sb1111111111111100000000000000001000000000000000;
		3391: Delta = 46'sb0000000000000011111111111111111000000000000000;
		5525: Delta = 46'sb1111111111111011111111111111111000000000000000;
		12021: Delta = 46'sb0000000000001000000000000000001000000000000000;
		16289: Delta = 46'sb1111111111111000000000000000001000000000000000;
		2324: Delta = 46'sb0000000000000111111111111111111000000000000000;
		6592: Delta = 46'sb1111111111110111111111111111111000000000000000;
		9887: Delta = 46'sb0000000000010000000000000000001000000000000000;
		18423: Delta = 46'sb1111111111110000000000000000001000000000000000;
		190: Delta = 46'sb0000000000001111111111111111111000000000000000;
		8726: Delta = 46'sb1111111111101111111111111111111000000000000000;
		5619: Delta = 46'sb0000000000100000000000000000001000000000000000;
		4078: Delta = 46'sb1111111111100000000000000000001000000000000000;
		14535: Delta = 46'sb0000000000011111111111111111111000000000000000;
		12994: Delta = 46'sb1111111111011111111111111111111000000000000000;
		15696: Delta = 46'sb0000000001000000000000000000001000000000000000;
		12614: Delta = 46'sb1111111111000000000000000000001000000000000000;
		5999: Delta = 46'sb0000000000111111111111111111111000000000000000;
		2917: Delta = 46'sb1111111110111111111111111111111000000000000000;
		17237: Delta = 46'sb0000000010000000000000000000001000000000000000;
		11073: Delta = 46'sb1111111110000000000000000000001000000000000000;
		7540: Delta = 46'sb0000000001111111111111111111111000000000000000;
		1376: Delta = 46'sb1111111101111111111111111111111000000000000000;
		1706: Delta = 46'sb0000000100000000000000000000001000000000000000;
		7991: Delta = 46'sb1111111100000000000000000000001000000000000000;
		10622: Delta = 46'sb0000000011111111111111111111111000000000000000;
		16907: Delta = 46'sb1111111011111111111111111111111000000000000000;
		7870: Delta = 46'sb0000001000000000000000000000001000000000000000;
		1827: Delta = 46'sb1111111000000000000000000000001000000000000000;
		16786: Delta = 46'sb0000000111111111111111111111111000000000000000;
		10743: Delta = 46'sb1111110111111111111111111111111000000000000000;
		1585: Delta = 46'sb0000010000000000000000000000001000000000000000;
		8112: Delta = 46'sb1111110000000000000000000000001000000000000000;
		10501: Delta = 46'sb0000001111111111111111111111111000000000000000;
		17028: Delta = 46'sb1111101111111111111111111111111000000000000000;
		7628: Delta = 46'sb0000100000000000000000000000001000000000000000;
		2069: Delta = 46'sb1111100000000000000000000000001000000000000000;
		16544: Delta = 46'sb0000011111111111111111111111111000000000000000;
		10985: Delta = 46'sb1111011111111111111111111111111000000000000000;
		1101: Delta = 46'sb0001000000000000000000000000001000000000000000;
		8596: Delta = 46'sb1111000000000000000000000000001000000000000000;
		10017: Delta = 46'sb0000111111111111111111111111111000000000000000;
		17512: Delta = 46'sb1110111111111111111111111111111000000000000000;
		6660: Delta = 46'sb0010000000000000000000000000001000000000000000;
		3037: Delta = 46'sb1110000000000000000000000000001000000000000000;
		15576: Delta = 46'sb0001111111111111111111111111111000000000000000;
		11953: Delta = 46'sb1101111111111111111111111111111000000000000000;
		17778: Delta = 46'sb0100000000000000000000000000001000000000000000;
		10532: Delta = 46'sb1100000000000000000000000000001000000000000000;
		8081: Delta = 46'sb0011111111111111111111111111111000000000000000;
		835: Delta = 46'sb1011111111111111111111111111111000000000000000;
		10478: Delta = 46'sb0000000000000000000000000000110000000000000000;
		8135: Delta = 46'sb1111111111111111111111111111010000000000000000;
		11259: Delta = 46'sb0000000000000000000000000001010000000000000000;
		7354: Delta = 46'sb1111111111111111111111111110110000000000000000;
		12821: Delta = 46'sb0000000000000000000000000010010000000000000000;
		6573: Delta = 46'sb1111111111111111111111111110010000000000000000;
		12040: Delta = 46'sb0000000000000000000000000001110000000000000000;
		5792: Delta = 46'sb1111111111111111111111111101110000000000000000;
		15945: Delta = 46'sb0000000000000000000000000100010000000000000000;
		3449: Delta = 46'sb1111111111111111111111111100010000000000000000;
		15164: Delta = 46'sb0000000000000000000000000011110000000000000000;
		2668: Delta = 46'sb1111111111111111111111111011110000000000000000;
		3580: Delta = 46'sb0000000000000000000000001000010000000000000000;
		15814: Delta = 46'sb1111111111111111111111111000010000000000000000;
		2799: Delta = 46'sb0000000000000000000000000111110000000000000000;
		15033: Delta = 46'sb1111111111111111111111110111110000000000000000;
		16076: Delta = 46'sb0000000000000000000000010000010000000000000000;
		3318: Delta = 46'sb1111111111111111111111110000010000000000000000;
		15295: Delta = 46'sb0000000000000000000000001111110000000000000000;
		2537: Delta = 46'sb1111111111111111111111101111110000000000000000;
		3842: Delta = 46'sb0000000000000000000000100000010000000000000000;
		15552: Delta = 46'sb1111111111111111111111100000010000000000000000;
		3061: Delta = 46'sb0000000000000000000000011111110000000000000000;
		14771: Delta = 46'sb1111111111111111111111011111110000000000000000;
		16600: Delta = 46'sb0000000000000000000001000000010000000000000000;
		2794: Delta = 46'sb1111111111111111111111000000010000000000000000;
		15819: Delta = 46'sb0000000000000000000000111111110000000000000000;
		2013: Delta = 46'sb1111111111111111111110111111110000000000000000;
		4890: Delta = 46'sb0000000000000000000010000000010000000000000000;
		14504: Delta = 46'sb1111111111111111111110000000010000000000000000;
		4109: Delta = 46'sb0000000000000000000001111111110000000000000000;
		13723: Delta = 46'sb1111111111111111111101111111110000000000000000;
		83: Delta = 46'sb0000000000000000000100000000010000000000000000;
		698: Delta = 46'sb1111111111111111111100000000010000000000000000;
		17915: Delta = 46'sb0000000000000000000011111111110000000000000000;
		18530: Delta = 46'sb1111111111111111111011111111110000000000000000;
		9082: Delta = 46'sb0000000000000000001000000000010000000000000000;
		10312: Delta = 46'sb1111111111111111111000000000010000000000000000;
		8301: Delta = 46'sb0000000000000000000111111111110000000000000000;
		9531: Delta = 46'sb1111111111111111110111111111110000000000000000;
		8467: Delta = 46'sb0000000000000000010000000000010000000000000000;
		10927: Delta = 46'sb1111111111111111110000000000010000000000000000;
		7686: Delta = 46'sb0000000000000000001111111111110000000000000000;
		10146: Delta = 46'sb1111111111111111101111111111110000000000000000;
		7237: Delta = 46'sb0000000000000000100000000000010000000000000000;
		12157: Delta = 46'sb1111111111111111100000000000010000000000000000;
		6456: Delta = 46'sb0000000000000000011111111111110000000000000000;
		11376: Delta = 46'sb1111111111111111011111111111110000000000000000;
		4777: Delta = 46'sb0000000000000001000000000000010000000000000000;
		14617: Delta = 46'sb1111111111111111000000000000010000000000000000;
		3996: Delta = 46'sb0000000000000000111111111111110000000000000000;
		13836: Delta = 46'sb1111111111111110111111111111110000000000000000;
		18470: Delta = 46'sb0000000000000010000000000000010000000000000000;
		924: Delta = 46'sb1111111111111110000000000000010000000000000000;
		17689: Delta = 46'sb0000000000000001111111111111110000000000000000;
		143: Delta = 46'sb1111111111111101111111111111110000000000000000;
		8630: Delta = 46'sb0000000000000100000000000000010000000000000000;
		10764: Delta = 46'sb1111111111111100000000000000010000000000000000;
		7849: Delta = 46'sb0000000000000011111111111111110000000000000000;
		9983: Delta = 46'sb1111111111111011111111111111110000000000000000;
		7563: Delta = 46'sb0000000000001000000000000000010000000000000000;
		11831: Delta = 46'sb1111111111111000000000000000010000000000000000;
		6782: Delta = 46'sb0000000000000111111111111111110000000000000000;
		11050: Delta = 46'sb1111111111110111111111111111110000000000000000;
		5429: Delta = 46'sb0000000000010000000000000000010000000000000000;
		13965: Delta = 46'sb1111111111110000000000000000010000000000000000;
		4648: Delta = 46'sb0000000000001111111111111111110000000000000000;
		13184: Delta = 46'sb1111111111101111111111111111110000000000000000;
		1161: Delta = 46'sb0000000000100000000000000000010000000000000000;
		18233: Delta = 46'sb1111111111100000000000000000010000000000000000;
		380: Delta = 46'sb0000000000011111111111111111110000000000000000;
		17452: Delta = 46'sb1111111111011111111111111111110000000000000000;
		11238: Delta = 46'sb0000000001000000000000000000010000000000000000;
		8156: Delta = 46'sb1111111111000000000000000000010000000000000000;
		10457: Delta = 46'sb0000000000111111111111111111110000000000000000;
		7375: Delta = 46'sb1111111110111111111111111111110000000000000000;
		12779: Delta = 46'sb0000000010000000000000000000010000000000000000;
		6615: Delta = 46'sb1111111110000000000000000000010000000000000000;
		11998: Delta = 46'sb0000000001111111111111111111110000000000000000;
		5834: Delta = 46'sb1111111101111111111111111111110000000000000000;
		15861: Delta = 46'sb0000000100000000000000000000010000000000000000;
		3533: Delta = 46'sb1111111100000000000000000000010000000000000000;
		15080: Delta = 46'sb0000000011111111111111111111110000000000000000;
		2752: Delta = 46'sb1111111011111111111111111111110000000000000000;
		3412: Delta = 46'sb0000001000000000000000000000010000000000000000;
		15982: Delta = 46'sb1111111000000000000000000000010000000000000000;
		2631: Delta = 46'sb0000000111111111111111111111110000000000000000;
		15201: Delta = 46'sb1111110111111111111111111111110000000000000000;
		15740: Delta = 46'sb0000010000000000000000000000010000000000000000;
		3654: Delta = 46'sb1111110000000000000000000000010000000000000000;
		14959: Delta = 46'sb0000001111111111111111111111110000000000000000;
		2873: Delta = 46'sb1111101111111111111111111111110000000000000000;
		3170: Delta = 46'sb0000100000000000000000000000010000000000000000;
		16224: Delta = 46'sb1111100000000000000000000000010000000000000000;
		2389: Delta = 46'sb0000011111111111111111111111110000000000000000;
		15443: Delta = 46'sb1111011111111111111111111111110000000000000000;
		15256: Delta = 46'sb0001000000000000000000000000010000000000000000;
		4138: Delta = 46'sb1111000000000000000000000000010000000000000000;
		14475: Delta = 46'sb0000111111111111111111111111110000000000000000;
		3357: Delta = 46'sb1110111111111111111111111111110000000000000000;
		2202: Delta = 46'sb0010000000000000000000000000010000000000000000;
		17192: Delta = 46'sb1110000000000000000000000000010000000000000000;
		1421: Delta = 46'sb0001111111111111111111111111110000000000000000;
		16411: Delta = 46'sb1101111111111111111111111111110000000000000000;
		13320: Delta = 46'sb0100000000000000000000000000010000000000000000;
		6074: Delta = 46'sb1100000000000000000000000000010000000000000000;
		12539: Delta = 46'sb0011111111111111111111111111110000000000000000;
		5293: Delta = 46'sb1011111111111111111111111111110000000000000000;
		2343: Delta = 46'sb0000000000000000000000000001100000000000000000;
		16270: Delta = 46'sb1111111111111111111111111110100000000000000000;
		3905: Delta = 46'sb0000000000000000000000000010100000000000000000;
		14708: Delta = 46'sb1111111111111111111111111101100000000000000000;
		7029: Delta = 46'sb0000000000000000000000000100100000000000000000;
		13146: Delta = 46'sb1111111111111111111111111100100000000000000000;
		5467: Delta = 46'sb0000000000000000000000000011100000000000000000;
		11584: Delta = 46'sb1111111111111111111111111011100000000000000000;
		13277: Delta = 46'sb0000000000000000000000001000100000000000000000;
		6898: Delta = 46'sb1111111111111111111111111000100000000000000000;
		11715: Delta = 46'sb0000000000000000000000000111100000000000000000;
		5336: Delta = 46'sb1111111111111111111111110111100000000000000000;
		7160: Delta = 46'sb0000000000000000000000010000100000000000000000;
		13015: Delta = 46'sb1111111111111111111111110000100000000000000000;
		5598: Delta = 46'sb0000000000000000000000001111100000000000000000;
		11453: Delta = 46'sb1111111111111111111111101111100000000000000000;
		13539: Delta = 46'sb0000000000000000000000100000100000000000000000;
		6636: Delta = 46'sb1111111111111111111111100000100000000000000000;
		11977: Delta = 46'sb0000000000000000000000011111100000000000000000;
		5074: Delta = 46'sb1111111111111111111111011111100000000000000000;
		7684: Delta = 46'sb0000000000000000000001000000100000000000000000;
		12491: Delta = 46'sb1111111111111111111111000000100000000000000000;
		6122: Delta = 46'sb0000000000000000000000111111100000000000000000;
		10929: Delta = 46'sb1111111111111111111110111111100000000000000000;
		14587: Delta = 46'sb0000000000000000000010000000100000000000000000;
		5588: Delta = 46'sb1111111111111111111110000000100000000000000000;
		13025: Delta = 46'sb0000000000000000000001111111100000000000000000;
		4026: Delta = 46'sb1111111111111111111101111111100000000000000000;
		9780: Delta = 46'sb0000000000000000000100000000100000000000000000;
		10395: Delta = 46'sb1111111111111111111100000000100000000000000000;
		8218: Delta = 46'sb0000000000000000000011111111100000000000000000;
		8833: Delta = 46'sb1111111111111111111011111111100000000000000000;
		166: Delta = 46'sb0000000000000000001000000000100000000000000000;
		1396: Delta = 46'sb1111111111111111111000000000100000000000000000;
		17217: Delta = 46'sb0000000000000000000111111111100000000000000000;
		18447: Delta = 46'sb1111111111111111110111111111100000000000000000;
		18164: Delta = 46'sb0000000000000000010000000000100000000000000000;
		2011: Delta = 46'sb1111111111111111110000000000100000000000000000;
		16602: Delta = 46'sb0000000000000000001111111111100000000000000000;
		449: Delta = 46'sb1111111111111111101111111111100000000000000000;
		16934: Delta = 46'sb0000000000000000100000000000100000000000000000;
		3241: Delta = 46'sb1111111111111111100000000000100000000000000000;
		15372: Delta = 46'sb0000000000000000011111111111100000000000000000;
		1679: Delta = 46'sb1111111111111111011111111111100000000000000000;
		14474: Delta = 46'sb0000000000000001000000000000100000000000000000;
		5701: Delta = 46'sb1111111111111111000000000000100000000000000000;
		12912: Delta = 46'sb0000000000000000111111111111100000000000000000;
		4139: Delta = 46'sb1111111111111110111111111111100000000000000000;
		9554: Delta = 46'sb0000000000000010000000000000100000000000000000;
		10621: Delta = 46'sb1111111111111110000000000000100000000000000000;
		7992: Delta = 46'sb0000000000000001111111111111100000000000000000;
		9059: Delta = 46'sb1111111111111101111111111111100000000000000000;
		18327: Delta = 46'sb0000000000000100000000000000100000000000000000;
		1848: Delta = 46'sb1111111111111100000000000000100000000000000000;
		16765: Delta = 46'sb0000000000000011111111111111100000000000000000;
		286: Delta = 46'sb1111111111111011111111111111100000000000000000;
		17260: Delta = 46'sb0000000000001000000000000000100000000000000000;
		2915: Delta = 46'sb1111111111111000000000000000100000000000000000;
		15698: Delta = 46'sb0000000000000111111111111111100000000000000000;
		1353: Delta = 46'sb1111111111110111111111111111100000000000000000;
		15126: Delta = 46'sb0000000000010000000000000000100000000000000000;
		5049: Delta = 46'sb1111111111110000000000000000100000000000000000;
		13564: Delta = 46'sb0000000000001111111111111111100000000000000000;
		3487: Delta = 46'sb1111111111101111111111111111100000000000000000;
		10858: Delta = 46'sb0000000000100000000000000000100000000000000000;
		9317: Delta = 46'sb1111111111100000000000000000100000000000000000;
		9296: Delta = 46'sb0000000000011111111111111111100000000000000000;
		7755: Delta = 46'sb1111111111011111111111111111100000000000000000;
		2322: Delta = 46'sb0000000001000000000000000000100000000000000000;
		17853: Delta = 46'sb1111111111000000000000000000100000000000000000;
		760: Delta = 46'sb0000000000111111111111111111100000000000000000;
		16291: Delta = 46'sb1111111110111111111111111111100000000000000000;
		3863: Delta = 46'sb0000000010000000000000000000100000000000000000;
		16312: Delta = 46'sb1111111110000000000000000000100000000000000000;
		2301: Delta = 46'sb0000000001111111111111111111100000000000000000;
		14750: Delta = 46'sb1111111101111111111111111111100000000000000000;
		6945: Delta = 46'sb0000000100000000000000000000100000000000000000;
		13230: Delta = 46'sb1111111100000000000000000000100000000000000000;
		5383: Delta = 46'sb0000000011111111111111111111100000000000000000;
		11668: Delta = 46'sb1111111011111111111111111111100000000000000000;
		13109: Delta = 46'sb0000001000000000000000000000100000000000000000;
		7066: Delta = 46'sb1111111000000000000000000000100000000000000000;
		11547: Delta = 46'sb0000000111111111111111111111100000000000000000;
		5504: Delta = 46'sb1111110111111111111111111111100000000000000000;
		6824: Delta = 46'sb0000010000000000000000000000100000000000000000;
		13351: Delta = 46'sb1111110000000000000000000000100000000000000000;
		5262: Delta = 46'sb0000001111111111111111111111100000000000000000;
		11789: Delta = 46'sb1111101111111111111111111111100000000000000000;
		12867: Delta = 46'sb0000100000000000000000000000100000000000000000;
		7308: Delta = 46'sb1111100000000000000000000000100000000000000000;
		11305: Delta = 46'sb0000011111111111111111111111100000000000000000;
		5746: Delta = 46'sb1111011111111111111111111111100000000000000000;
		6340: Delta = 46'sb0001000000000000000000000000100000000000000000;
		13835: Delta = 46'sb1111000000000000000000000000100000000000000000;
		4778: Delta = 46'sb0000111111111111111111111111100000000000000000;
		12273: Delta = 46'sb1110111111111111111111111111100000000000000000;
		11899: Delta = 46'sb0010000000000000000000000000100000000000000000;
		8276: Delta = 46'sb1110000000000000000000000000100000000000000000;
		10337: Delta = 46'sb0001111111111111111111111111100000000000000000;
		6714: Delta = 46'sb1101111111111111111111111111100000000000000000;
		4404: Delta = 46'sb0100000000000000000000000000100000000000000000;
		15771: Delta = 46'sb1100000000000000000000000000100000000000000000;
		2842: Delta = 46'sb0011111111111111111111111111100000000000000000;
		14209: Delta = 46'sb1011111111111111111111111111100000000000000000;
		4686: Delta = 46'sb0000000000000000000000000011000000000000000000;
		13927: Delta = 46'sb1111111111111111111111111101000000000000000000;
		7810: Delta = 46'sb0000000000000000000000000101000000000000000000;
		10803: Delta = 46'sb1111111111111111111111111011000000000000000000;
		14058: Delta = 46'sb0000000000000000000000001001000000000000000000;
		7679: Delta = 46'sb1111111111111111111111111001000000000000000000;
		10934: Delta = 46'sb0000000000000000000000000111000000000000000000;
		4555: Delta = 46'sb1111111111111111111111110111000000000000000000;
		7941: Delta = 46'sb0000000000000000000000010001000000000000000000;
		13796: Delta = 46'sb1111111111111111111111110001000000000000000000;
		4817: Delta = 46'sb0000000000000000000000001111000000000000000000;
		10672: Delta = 46'sb1111111111111111111111101111000000000000000000;
		14320: Delta = 46'sb0000000000000000000000100001000000000000000000;
		7417: Delta = 46'sb1111111111111111111111100001000000000000000000;
		11196: Delta = 46'sb0000000000000000000000011111000000000000000000;
		4293: Delta = 46'sb1111111111111111111111011111000000000000000000;
		8465: Delta = 46'sb0000000000000000000001000001000000000000000000;
		13272: Delta = 46'sb1111111111111111111111000001000000000000000000;
		5341: Delta = 46'sb0000000000000000000000111111000000000000000000;
		10148: Delta = 46'sb1111111111111111111110111111000000000000000000;
		15368: Delta = 46'sb0000000000000000000010000001000000000000000000;
		6369: Delta = 46'sb1111111111111111111110000001000000000000000000;
		12244: Delta = 46'sb0000000000000000000001111111000000000000000000;
		3245: Delta = 46'sb1111111111111111111101111111000000000000000000;
		10561: Delta = 46'sb0000000000000000000100000001000000000000000000;
		11176: Delta = 46'sb1111111111111111111100000001000000000000000000;
		7437: Delta = 46'sb0000000000000000000011111111000000000000000000;
		8052: Delta = 46'sb1111111111111111111011111111000000000000000000;
		947: Delta = 46'sb0000000000000000001000000001000000000000000000;
		2177: Delta = 46'sb1111111111111111111000000001000000000000000000;
		16436: Delta = 46'sb0000000000000000000111111111000000000000000000;
		17666: Delta = 46'sb1111111111111111110111111111000000000000000000;
		332: Delta = 46'sb0000000000000000010000000001000000000000000000;
		2792: Delta = 46'sb1111111111111111110000000001000000000000000000;
		15821: Delta = 46'sb0000000000000000001111111111000000000000000000;
		18281: Delta = 46'sb1111111111111111101111111111000000000000000000;
		17715: Delta = 46'sb0000000000000000100000000001000000000000000000;
		4022: Delta = 46'sb1111111111111111100000000001000000000000000000;
		14591: Delta = 46'sb0000000000000000011111111111000000000000000000;
		898: Delta = 46'sb1111111111111111011111111111000000000000000000;
		15255: Delta = 46'sb0000000000000001000000000001000000000000000000;
		6482: Delta = 46'sb1111111111111111000000000001000000000000000000;
		12131: Delta = 46'sb0000000000000000111111111111000000000000000000;
		3358: Delta = 46'sb1111111111111110111111111111000000000000000000;
		10335: Delta = 46'sb0000000000000010000000000001000000000000000000;
		11402: Delta = 46'sb1111111111111110000000000001000000000000000000;
		7211: Delta = 46'sb0000000000000001111111111111000000000000000000;
		8278: Delta = 46'sb1111111111111101111111111111000000000000000000;
		495: Delta = 46'sb0000000000000100000000000001000000000000000000;
		2629: Delta = 46'sb1111111111111100000000000001000000000000000000;
		15984: Delta = 46'sb0000000000000011111111111111000000000000000000;
		18118: Delta = 46'sb1111111111111011111111111111000000000000000000;
		18041: Delta = 46'sb0000000000001000000000000001000000000000000000;
		3696: Delta = 46'sb1111111111111000000000000001000000000000000000;
		14917: Delta = 46'sb0000000000000111111111111111000000000000000000;
		572: Delta = 46'sb1111111111110111111111111111000000000000000000;
		15907: Delta = 46'sb0000000000010000000000000001000000000000000000;
		5830: Delta = 46'sb1111111111110000000000000001000000000000000000;
		12783: Delta = 46'sb0000000000001111111111111111000000000000000000;
		2706: Delta = 46'sb1111111111101111111111111111000000000000000000;
		11639: Delta = 46'sb0000000000100000000000000001000000000000000000;
		10098: Delta = 46'sb1111111111100000000000000001000000000000000000;
		8515: Delta = 46'sb0000000000011111111111111111000000000000000000;
		6974: Delta = 46'sb1111111111011111111111111111000000000000000000;
		3103: Delta = 46'sb0000000001000000000000000001000000000000000000;
		21: Delta = 46'sb1111111111000000000000000001000000000000000000;
		18592: Delta = 46'sb0000000000111111111111111111000000000000000000;
		15510: Delta = 46'sb1111111110111111111111111111000000000000000000;
		4644: Delta = 46'sb0000000010000000000000000001000000000000000000;
		17093: Delta = 46'sb1111111110000000000000000001000000000000000000;
		1520: Delta = 46'sb0000000001111111111111111111000000000000000000;
		13969: Delta = 46'sb1111111101111111111111111111000000000000000000;
		7726: Delta = 46'sb0000000100000000000000000001000000000000000000;
		14011: Delta = 46'sb1111111100000000000000000001000000000000000000;
		4602: Delta = 46'sb0000000011111111111111111111000000000000000000;
		10887: Delta = 46'sb1111111011111111111111111111000000000000000000;
		13890: Delta = 46'sb0000001000000000000000000001000000000000000000;
		7847: Delta = 46'sb1111111000000000000000000001000000000000000000;
		10766: Delta = 46'sb0000000111111111111111111111000000000000000000;
		4723: Delta = 46'sb1111110111111111111111111111000000000000000000;
		7605: Delta = 46'sb0000010000000000000000000001000000000000000000;
		14132: Delta = 46'sb1111110000000000000000000001000000000000000000;
		4481: Delta = 46'sb0000001111111111111111111111000000000000000000;
		11008: Delta = 46'sb1111101111111111111111111111000000000000000000;
		13648: Delta = 46'sb0000100000000000000000000001000000000000000000;
		8089: Delta = 46'sb1111100000000000000000000001000000000000000000;
		10524: Delta = 46'sb0000011111111111111111111111000000000000000000;
		4965: Delta = 46'sb1111011111111111111111111111000000000000000000;
		7121: Delta = 46'sb0001000000000000000000000001000000000000000000;
		14616: Delta = 46'sb1111000000000000000000000001000000000000000000;
		3997: Delta = 46'sb0000111111111111111111111111000000000000000000;
		11492: Delta = 46'sb1110111111111111111111111111000000000000000000;
		12680: Delta = 46'sb0010000000000000000000000001000000000000000000;
		9057: Delta = 46'sb1110000000000000000000000001000000000000000000;
		9556: Delta = 46'sb0001111111111111111111111111000000000000000000;
		5933: Delta = 46'sb1101111111111111111111111111000000000000000000;
		5185: Delta = 46'sb0100000000000000000000000001000000000000000000;
		16552: Delta = 46'sb1100000000000000000000000001000000000000000000;
		2061: Delta = 46'sb0011111111111111111111111111000000000000000000;
		13428: Delta = 46'sb1011111111111111111111111111000000000000000000;
		9372: Delta = 46'sb0000000000000000000000000110000000000000000000;
		9241: Delta = 46'sb1111111111111111111111111010000000000000000000;
		15620: Delta = 46'sb0000000000000000000000001010000000000000000000;
		2993: Delta = 46'sb1111111111111111111111110110000000000000000000;
		9503: Delta = 46'sb0000000000000000000000010010000000000000000000;
		15358: Delta = 46'sb1111111111111111111111110010000000000000000000;
		3255: Delta = 46'sb0000000000000000000000001110000000000000000000;
		9110: Delta = 46'sb1111111111111111111111101110000000000000000000;
		15882: Delta = 46'sb0000000000000000000000100010000000000000000000;
		8979: Delta = 46'sb1111111111111111111111100010000000000000000000;
		9634: Delta = 46'sb0000000000000000000000011110000000000000000000;
		2731: Delta = 46'sb1111111111111111111111011110000000000000000000;
		10027: Delta = 46'sb0000000000000000000001000010000000000000000000;
		14834: Delta = 46'sb1111111111111111111111000010000000000000000000;
		3779: Delta = 46'sb0000000000000000000000111110000000000000000000;
		8586: Delta = 46'sb1111111111111111111110111110000000000000000000;
		16930: Delta = 46'sb0000000000000000000010000010000000000000000000;
		7931: Delta = 46'sb1111111111111111111110000010000000000000000000;
		10682: Delta = 46'sb0000000000000000000001111110000000000000000000;
		1683: Delta = 46'sb1111111111111111111101111110000000000000000000;
		12123: Delta = 46'sb0000000000000000000100000010000000000000000000;
		12738: Delta = 46'sb1111111111111111111100000010000000000000000000;
		5875: Delta = 46'sb0000000000000000000011111110000000000000000000;
		6490: Delta = 46'sb1111111111111111111011111110000000000000000000;
		2509: Delta = 46'sb0000000000000000001000000010000000000000000000;
		3739: Delta = 46'sb1111111111111111111000000010000000000000000000;
		14874: Delta = 46'sb0000000000000000000111111110000000000000000000;
		16104: Delta = 46'sb1111111111111111110111111110000000000000000000;
		1894: Delta = 46'sb0000000000000000010000000010000000000000000000;
		4354: Delta = 46'sb1111111111111111110000000010000000000000000000;
		14259: Delta = 46'sb0000000000000000001111111110000000000000000000;
		16719: Delta = 46'sb1111111111111111101111111110000000000000000000;
		664: Delta = 46'sb0000000000000000100000000010000000000000000000;
		5584: Delta = 46'sb1111111111111111100000000010000000000000000000;
		13029: Delta = 46'sb0000000000000000011111111110000000000000000000;
		17949: Delta = 46'sb1111111111111111011111111110000000000000000000;
		16817: Delta = 46'sb0000000000000001000000000010000000000000000000;
		8044: Delta = 46'sb1111111111111111000000000010000000000000000000;
		10569: Delta = 46'sb0000000000000000111111111110000000000000000000;
		1796: Delta = 46'sb1111111111111110111111111110000000000000000000;
		11897: Delta = 46'sb0000000000000010000000000010000000000000000000;
		12964: Delta = 46'sb1111111111111110000000000010000000000000000000;
		5649: Delta = 46'sb0000000000000001111111111110000000000000000000;
		6716: Delta = 46'sb1111111111111101111111111110000000000000000000;
		2057: Delta = 46'sb0000000000000100000000000010000000000000000000;
		4191: Delta = 46'sb1111111111111100000000000010000000000000000000;
		14422: Delta = 46'sb0000000000000011111111111110000000000000000000;
		16556: Delta = 46'sb1111111111111011111111111110000000000000000000;
		990: Delta = 46'sb0000000000001000000000000010000000000000000000;
		5258: Delta = 46'sb1111111111111000000000000010000000000000000000;
		13355: Delta = 46'sb0000000000000111111111111110000000000000000000;
		17623: Delta = 46'sb1111111111110111111111111110000000000000000000;
		17469: Delta = 46'sb0000000000010000000000000010000000000000000000;
		7392: Delta = 46'sb1111111111110000000000000010000000000000000000;
		11221: Delta = 46'sb0000000000001111111111111110000000000000000000;
		1144: Delta = 46'sb1111111111101111111111111110000000000000000000;
		13201: Delta = 46'sb0000000000100000000000000010000000000000000000;
		11660: Delta = 46'sb1111111111100000000000000010000000000000000000;
		6953: Delta = 46'sb0000000000011111111111111110000000000000000000;
		5412: Delta = 46'sb1111111111011111111111111110000000000000000000;
		4665: Delta = 46'sb0000000001000000000000000010000000000000000000;
		1583: Delta = 46'sb1111111111000000000000000010000000000000000000;
		17030: Delta = 46'sb0000000000111111111111111110000000000000000000;
		13948: Delta = 46'sb1111111110111111111111111110000000000000000000;
		6206: Delta = 46'sb0000000010000000000000000010000000000000000000;
		42: Delta = 46'sb1111111110000000000000000010000000000000000000;
		18571: Delta = 46'sb0000000001111111111111111110000000000000000000;
		12407: Delta = 46'sb1111111101111111111111111110000000000000000000;
		9288: Delta = 46'sb0000000100000000000000000010000000000000000000;
		15573: Delta = 46'sb1111111100000000000000000010000000000000000000;
		3040: Delta = 46'sb0000000011111111111111111110000000000000000000;
		9325: Delta = 46'sb1111111011111111111111111110000000000000000000;
		15452: Delta = 46'sb0000001000000000000000000010000000000000000000;
		9409: Delta = 46'sb1111111000000000000000000010000000000000000000;
		9204: Delta = 46'sb0000000111111111111111111110000000000000000000;
		3161: Delta = 46'sb1111110111111111111111111110000000000000000000;
		9167: Delta = 46'sb0000010000000000000000000010000000000000000000;
		15694: Delta = 46'sb1111110000000000000000000010000000000000000000;
		2919: Delta = 46'sb0000001111111111111111111110000000000000000000;
		9446: Delta = 46'sb1111101111111111111111111110000000000000000000;
		15210: Delta = 46'sb0000100000000000000000000010000000000000000000;
		9651: Delta = 46'sb1111100000000000000000000010000000000000000000;
		8962: Delta = 46'sb0000011111111111111111111110000000000000000000;
		3403: Delta = 46'sb1111011111111111111111111110000000000000000000;
		8683: Delta = 46'sb0001000000000000000000000010000000000000000000;
		16178: Delta = 46'sb1111000000000000000000000010000000000000000000;
		2435: Delta = 46'sb0000111111111111111111111110000000000000000000;
		9930: Delta = 46'sb1110111111111111111111111110000000000000000000;
		14242: Delta = 46'sb0010000000000000000000000010000000000000000000;
		10619: Delta = 46'sb1110000000000000000000000010000000000000000000;
		7994: Delta = 46'sb0001111111111111111111111110000000000000000000;
		4371: Delta = 46'sb1101111111111111111111111110000000000000000000;
		6747: Delta = 46'sb0100000000000000000000000010000000000000000000;
		18114: Delta = 46'sb1100000000000000000000000010000000000000000000;
		499: Delta = 46'sb0011111111111111111111111110000000000000000000;
		11866: Delta = 46'sb1011111111111111111111111110000000000000000000;
		131: Delta = 46'sb0000000000000000000000001100000000000000000000;
		18482: Delta = 46'sb1111111111111111111111110100000000000000000000;
		12627: Delta = 46'sb0000000000000000000000010100000000000000000000;
		5986: Delta = 46'sb1111111111111111111111101100000000000000000000;
		393: Delta = 46'sb0000000000000000000000100100000000000000000000;
		12103: Delta = 46'sb1111111111111111111111100100000000000000000000;
		6510: Delta = 46'sb0000000000000000000000011100000000000000000000;
		18220: Delta = 46'sb1111111111111111111111011100000000000000000000;
		13151: Delta = 46'sb0000000000000000000001000100000000000000000000;
		17958: Delta = 46'sb1111111111111111111111000100000000000000000000;
		655: Delta = 46'sb0000000000000000000000111100000000000000000000;
		5462: Delta = 46'sb1111111111111111111110111100000000000000000000;
		1441: Delta = 46'sb0000000000000000000010000100000000000000000000;
		11055: Delta = 46'sb1111111111111111111110000100000000000000000000;
		7558: Delta = 46'sb0000000000000000000001111100000000000000000000;
		17172: Delta = 46'sb1111111111111111111101111100000000000000000000;
		15247: Delta = 46'sb0000000000000000000100000100000000000000000000;
		15862: Delta = 46'sb1111111111111111111100000100000000000000000000;
		2751: Delta = 46'sb0000000000000000000011111100000000000000000000;
		3366: Delta = 46'sb1111111111111111111011111100000000000000000000;
		5633: Delta = 46'sb0000000000000000001000000100000000000000000000;
		6863: Delta = 46'sb1111111111111111111000000100000000000000000000;
		11750: Delta = 46'sb0000000000000000000111111100000000000000000000;
		12980: Delta = 46'sb1111111111111111110111111100000000000000000000;
		5018: Delta = 46'sb0000000000000000010000000100000000000000000000;
		7478: Delta = 46'sb1111111111111111110000000100000000000000000000;
		11135: Delta = 46'sb0000000000000000001111111100000000000000000000;
		13595: Delta = 46'sb1111111111111111101111111100000000000000000000;
		3788: Delta = 46'sb0000000000000000100000000100000000000000000000;
		8708: Delta = 46'sb1111111111111111100000000100000000000000000000;
		9905: Delta = 46'sb0000000000000000011111111100000000000000000000;
		14825: Delta = 46'sb1111111111111111011111111100000000000000000000;
		1328: Delta = 46'sb0000000000000001000000000100000000000000000000;
		11168: Delta = 46'sb1111111111111111000000000100000000000000000000;
		7445: Delta = 46'sb0000000000000000111111111100000000000000000000;
		17285: Delta = 46'sb1111111111111110111111111100000000000000000000;
		15021: Delta = 46'sb0000000000000010000000000100000000000000000000;
		16088: Delta = 46'sb1111111111111110000000000100000000000000000000;
		2525: Delta = 46'sb0000000000000001111111111100000000000000000000;
		3592: Delta = 46'sb1111111111111101111111111100000000000000000000;
		5181: Delta = 46'sb0000000000000100000000000100000000000000000000;
		7315: Delta = 46'sb1111111111111100000000000100000000000000000000;
		11298: Delta = 46'sb0000000000000011111111111100000000000000000000;
		13432: Delta = 46'sb1111111111111011111111111100000000000000000000;
		4114: Delta = 46'sb0000000000001000000000000100000000000000000000;
		8382: Delta = 46'sb1111111111111000000000000100000000000000000000;
		10231: Delta = 46'sb0000000000000111111111111100000000000000000000;
		14499: Delta = 46'sb1111111111110111111111111100000000000000000000;
		1980: Delta = 46'sb0000000000010000000000000100000000000000000000;
		10516: Delta = 46'sb1111111111110000000000000100000000000000000000;
		8097: Delta = 46'sb0000000000001111111111111100000000000000000000;
		16633: Delta = 46'sb1111111111101111111111111100000000000000000000;
		16325: Delta = 46'sb0000000000100000000000000100000000000000000000;
		14784: Delta = 46'sb1111111111100000000000000100000000000000000000;
		3829: Delta = 46'sb0000000000011111111111111100000000000000000000;
		2288: Delta = 46'sb1111111111011111111111111100000000000000000000;
		7789: Delta = 46'sb0000000001000000000000000100000000000000000000;
		4707: Delta = 46'sb1111111111000000000000000100000000000000000000;
		13906: Delta = 46'sb0000000000111111111111111100000000000000000000;
		10824: Delta = 46'sb1111111110111111111111111100000000000000000000;
		9330: Delta = 46'sb0000000010000000000000000100000000000000000000;
		3166: Delta = 46'sb1111111110000000000000000100000000000000000000;
		15447: Delta = 46'sb0000000001111111111111111100000000000000000000;
		9283: Delta = 46'sb1111111101111111111111111100000000000000000000;
		12412: Delta = 46'sb0000000100000000000000000100000000000000000000;
		84: Delta = 46'sb1111111100000000000000000100000000000000000000;
		18529: Delta = 46'sb0000000011111111111111111100000000000000000000;
		6201: Delta = 46'sb1111111011111111111111111100000000000000000000;
		18576: Delta = 46'sb0000001000000000000000000100000000000000000000;
		12533: Delta = 46'sb1111111000000000000000000100000000000000000000;
		6080: Delta = 46'sb0000000111111111111111111100000000000000000000;
		37: Delta = 46'sb1111110111111111111111111100000000000000000000;
		12291: Delta = 46'sb0000010000000000000000000100000000000000000000;
		205: Delta = 46'sb1111110000000000000000000100000000000000000000;
		18408: Delta = 46'sb0000001111111111111111111100000000000000000000;
		6322: Delta = 46'sb1111101111111111111111111100000000000000000000;
		18334: Delta = 46'sb0000100000000000000000000100000000000000000000;
		12775: Delta = 46'sb1111100000000000000000000100000000000000000000;
		5838: Delta = 46'sb0000011111111111111111111100000000000000000000;
		279: Delta = 46'sb1111011111111111111111111100000000000000000000;
		11807: Delta = 46'sb0001000000000000000000000100000000000000000000;
		689: Delta = 46'sb1111000000000000000000000100000000000000000000;
		17924: Delta = 46'sb0000111111111111111111111100000000000000000000;
		6806: Delta = 46'sb1110111111111111111111111100000000000000000000;
		17366: Delta = 46'sb0010000000000000000000000100000000000000000000;
		13743: Delta = 46'sb1110000000000000000000000100000000000000000000;
		4870: Delta = 46'sb0001111111111111111111111100000000000000000000;
		1247: Delta = 46'sb1101111111111111111111111100000000000000000000;
		9871: Delta = 46'sb0100000000000000000000000100000000000000000000;
		2625: Delta = 46'sb1100000000000000000000000100000000000000000000;
		15988: Delta = 46'sb0011111111111111111111111100000000000000000000;
		8742: Delta = 46'sb1011111111111111111111111100000000000000000000;
		262: Delta = 46'sb0000000000000000000000011000000000000000000000;
		18351: Delta = 46'sb1111111111111111111111101000000000000000000000;
		6641: Delta = 46'sb0000000000000000000000101000000000000000000000;
		11972: Delta = 46'sb1111111111111111111111011000000000000000000000;
		786: Delta = 46'sb0000000000000000000001001000000000000000000000;
		5593: Delta = 46'sb1111111111111111111111001000000000000000000000;
		13020: Delta = 46'sb0000000000000000000000111000000000000000000000;
		17827: Delta = 46'sb1111111111111111111110111000000000000000000000;
		7689: Delta = 46'sb0000000000000000000010001000000000000000000000;
		17303: Delta = 46'sb1111111111111111111110001000000000000000000000;
		1310: Delta = 46'sb0000000000000000000001111000000000000000000000;
		10924: Delta = 46'sb1111111111111111111101111000000000000000000000;
		2882: Delta = 46'sb0000000000000000000100001000000000000000000000;
		3497: Delta = 46'sb1111111111111111111100001000000000000000000000;
		15116: Delta = 46'sb0000000000000000000011111000000000000000000000;
		15731: Delta = 46'sb1111111111111111111011111000000000000000000000;
		11881: Delta = 46'sb0000000000000000001000001000000000000000000000;
		13111: Delta = 46'sb1111111111111111111000001000000000000000000000;
		5502: Delta = 46'sb0000000000000000000111111000000000000000000000;
		6732: Delta = 46'sb1111111111111111110111111000000000000000000000;
		11266: Delta = 46'sb0000000000000000010000001000000000000000000000;
		13726: Delta = 46'sb1111111111111111110000001000000000000000000000;
		4887: Delta = 46'sb0000000000000000001111111000000000000000000000;
		7347: Delta = 46'sb1111111111111111101111111000000000000000000000;
		10036: Delta = 46'sb0000000000000000100000001000000000000000000000;
		14956: Delta = 46'sb1111111111111111100000001000000000000000000000;
		3657: Delta = 46'sb0000000000000000011111111000000000000000000000;
		8577: Delta = 46'sb1111111111111111011111111000000000000000000000;
		7576: Delta = 46'sb0000000000000001000000001000000000000000000000;
		17416: Delta = 46'sb1111111111111111000000001000000000000000000000;
		1197: Delta = 46'sb0000000000000000111111111000000000000000000000;
		11037: Delta = 46'sb1111111111111110111111111000000000000000000000;
		2656: Delta = 46'sb0000000000000010000000001000000000000000000000;
		3723: Delta = 46'sb1111111111111110000000001000000000000000000000;
		14890: Delta = 46'sb0000000000000001111111111000000000000000000000;
		15957: Delta = 46'sb1111111111111101111111111000000000000000000000;
		11429: Delta = 46'sb0000000000000100000000001000000000000000000000;
		13563: Delta = 46'sb1111111111111100000000001000000000000000000000;
		5050: Delta = 46'sb0000000000000011111111111000000000000000000000;
		7184: Delta = 46'sb1111111111111011111111111000000000000000000000;
		10362: Delta = 46'sb0000000000001000000000001000000000000000000000;
		14630: Delta = 46'sb1111111111111000000000001000000000000000000000;
		3983: Delta = 46'sb0000000000000111111111111000000000000000000000;
		8251: Delta = 46'sb1111111111110111111111111000000000000000000000;
		8228: Delta = 46'sb0000000000010000000000001000000000000000000000;
		16764: Delta = 46'sb1111111111110000000000001000000000000000000000;
		1849: Delta = 46'sb0000000000001111111111111000000000000000000000;
		10385: Delta = 46'sb1111111111101111111111111000000000000000000000;
		3960: Delta = 46'sb0000000000100000000000001000000000000000000000;
		2419: Delta = 46'sb1111111111100000000000001000000000000000000000;
		16194: Delta = 46'sb0000000000011111111111111000000000000000000000;
		14653: Delta = 46'sb1111111111011111111111111000000000000000000000;
		14037: Delta = 46'sb0000000001000000000000001000000000000000000000;
		10955: Delta = 46'sb1111111111000000000000001000000000000000000000;
		7658: Delta = 46'sb0000000000111111111111111000000000000000000000;
		4576: Delta = 46'sb1111111110111111111111111000000000000000000000;
		15578: Delta = 46'sb0000000010000000000000001000000000000000000000;
		9414: Delta = 46'sb1111111110000000000000001000000000000000000000;
		9199: Delta = 46'sb0000000001111111111111111000000000000000000000;
		3035: Delta = 46'sb1111111101111111111111111000000000000000000000;
		47: Delta = 46'sb0000000100000000000000001000000000000000000000;
		6332: Delta = 46'sb1111111100000000000000001000000000000000000000;
		12281: Delta = 46'sb0000000011111111111111111000000000000000000000;
		18566: Delta = 46'sb1111111011111111111111111000000000000000000000;
		6211: Delta = 46'sb0000001000000000000000001000000000000000000000;
		168: Delta = 46'sb1111111000000000000000001000000000000000000000;
		18445: Delta = 46'sb0000000111111111111111111000000000000000000000;
		12402: Delta = 46'sb1111110111111111111111111000000000000000000000;
		18539: Delta = 46'sb0000010000000000000000001000000000000000000000;
		6453: Delta = 46'sb1111110000000000000000001000000000000000000000;
		12160: Delta = 46'sb0000001111111111111111111000000000000000000000;
		74: Delta = 46'sb1111101111111111111111111000000000000000000000;
		5969: Delta = 46'sb0000100000000000000000001000000000000000000000;
		410: Delta = 46'sb1111100000000000000000001000000000000000000000;
		18203: Delta = 46'sb0000011111111111111111111000000000000000000000;
		12644: Delta = 46'sb1111011111111111111111111000000000000000000000;
		18055: Delta = 46'sb0001000000000000000000001000000000000000000000;
		6937: Delta = 46'sb1111000000000000000000001000000000000000000000;
		11676: Delta = 46'sb0000111111111111111111111000000000000000000000;
		558: Delta = 46'sb1110111111111111111111111000000000000000000000;
		5001: Delta = 46'sb0010000000000000000000001000000000000000000000;
		1378: Delta = 46'sb1110000000000000000000001000000000000000000000;
		17235: Delta = 46'sb0001111111111111111111111000000000000000000000;
		13612: Delta = 46'sb1101111111111111111111111000000000000000000000;
		16119: Delta = 46'sb0100000000000000000000001000000000000000000000;
		8873: Delta = 46'sb1100000000000000000000001000000000000000000000;
		9740: Delta = 46'sb0011111111111111111111111000000000000000000000;
		2494: Delta = 46'sb1011111111111111111111111000000000000000000000;
		524: Delta = 46'sb0000000000000000000000110000000000000000000000;
		18089: Delta = 46'sb1111111111111111111111010000000000000000000000;
		13282: Delta = 46'sb0000000000000000000001010000000000000000000000;
		5331: Delta = 46'sb1111111111111111111110110000000000000000000000;
		1572: Delta = 46'sb0000000000000000000010010000000000000000000000;
		11186: Delta = 46'sb1111111111111111111110010000000000000000000000;
		7427: Delta = 46'sb0000000000000000000001110000000000000000000000;
		17041: Delta = 46'sb1111111111111111111101110000000000000000000000;
		15378: Delta = 46'sb0000000000000000000100010000000000000000000000;
		15993: Delta = 46'sb1111111111111111111100010000000000000000000000;
		2620: Delta = 46'sb0000000000000000000011110000000000000000000000;
		3235: Delta = 46'sb1111111111111111111011110000000000000000000000;
		5764: Delta = 46'sb0000000000000000001000010000000000000000000000;
		6994: Delta = 46'sb1111111111111111111000010000000000000000000000;
		11619: Delta = 46'sb0000000000000000000111110000000000000000000000;
		12849: Delta = 46'sb1111111111111111110111110000000000000000000000;
		5149: Delta = 46'sb0000000000000000010000010000000000000000000000;
		7609: Delta = 46'sb1111111111111111110000010000000000000000000000;
		11004: Delta = 46'sb0000000000000000001111110000000000000000000000;
		13464: Delta = 46'sb1111111111111111101111110000000000000000000000;
		3919: Delta = 46'sb0000000000000000100000010000000000000000000000;
		8839: Delta = 46'sb1111111111111111100000010000000000000000000000;
		9774: Delta = 46'sb0000000000000000011111110000000000000000000000;
		14694: Delta = 46'sb1111111111111111011111110000000000000000000000;
		1459: Delta = 46'sb0000000000000001000000010000000000000000000000;
		11299: Delta = 46'sb1111111111111111000000010000000000000000000000;
		7314: Delta = 46'sb0000000000000000111111110000000000000000000000;
		17154: Delta = 46'sb1111111111111110111111110000000000000000000000;
		15152: Delta = 46'sb0000000000000010000000010000000000000000000000;
		16219: Delta = 46'sb1111111111111110000000010000000000000000000000;
		2394: Delta = 46'sb0000000000000001111111110000000000000000000000;
		3461: Delta = 46'sb1111111111111101111111110000000000000000000000;
		5312: Delta = 46'sb0000000000000100000000010000000000000000000000;
		7446: Delta = 46'sb1111111111111100000000010000000000000000000000;
		11167: Delta = 46'sb0000000000000011111111110000000000000000000000;
		13301: Delta = 46'sb1111111111111011111111110000000000000000000000;
		4245: Delta = 46'sb0000000000001000000000010000000000000000000000;
		8513: Delta = 46'sb1111111111111000000000010000000000000000000000;
		10100: Delta = 46'sb0000000000000111111111110000000000000000000000;
		14368: Delta = 46'sb1111111111110111111111110000000000000000000000;
		2111: Delta = 46'sb0000000000010000000000010000000000000000000000;
		10647: Delta = 46'sb1111111111110000000000010000000000000000000000;
		7966: Delta = 46'sb0000000000001111111111110000000000000000000000;
		16502: Delta = 46'sb1111111111101111111111110000000000000000000000;
		16456: Delta = 46'sb0000000000100000000000010000000000000000000000;
		14915: Delta = 46'sb1111111111100000000000010000000000000000000000;
		3698: Delta = 46'sb0000000000011111111111110000000000000000000000;
		2157: Delta = 46'sb1111111111011111111111110000000000000000000000;
		7920: Delta = 46'sb0000000001000000000000010000000000000000000000;
		4838: Delta = 46'sb1111111111000000000000010000000000000000000000;
		13775: Delta = 46'sb0000000000111111111111110000000000000000000000;
		10693: Delta = 46'sb1111111110111111111111110000000000000000000000;
		9461: Delta = 46'sb0000000010000000000000010000000000000000000000;
		3297: Delta = 46'sb1111111110000000000000010000000000000000000000;
		15316: Delta = 46'sb0000000001111111111111110000000000000000000000;
		9152: Delta = 46'sb1111111101111111111111110000000000000000000000;
		12543: Delta = 46'sb0000000100000000000000010000000000000000000000;
		215: Delta = 46'sb1111111100000000000000010000000000000000000000;
		18398: Delta = 46'sb0000000011111111111111110000000000000000000000;
		6070: Delta = 46'sb1111111011111111111111110000000000000000000000;
		94: Delta = 46'sb0000001000000000000000010000000000000000000000;
		12664: Delta = 46'sb1111111000000000000000010000000000000000000000;
		5949: Delta = 46'sb0000000111111111111111110000000000000000000000;
		18519: Delta = 46'sb1111110111111111111111110000000000000000000000;
		12422: Delta = 46'sb0000010000000000000000010000000000000000000000;
		336: Delta = 46'sb1111110000000000000000010000000000000000000000;
		18277: Delta = 46'sb0000001111111111111111110000000000000000000000;
		6191: Delta = 46'sb1111101111111111111111110000000000000000000000;
		18465: Delta = 46'sb0000100000000000000000010000000000000000000000;
		12906: Delta = 46'sb1111100000000000000000010000000000000000000000;
		5707: Delta = 46'sb0000011111111111111111110000000000000000000000;
		148: Delta = 46'sb1111011111111111111111110000000000000000000000;
		11938: Delta = 46'sb0001000000000000000000010000000000000000000000;
		820: Delta = 46'sb1111000000000000000000010000000000000000000000;
		17793: Delta = 46'sb0000111111111111111111110000000000000000000000;
		6675: Delta = 46'sb1110111111111111111111110000000000000000000000;
		17497: Delta = 46'sb0010000000000000000000010000000000000000000000;
		13874: Delta = 46'sb1110000000000000000000010000000000000000000000;
		4739: Delta = 46'sb0001111111111111111111110000000000000000000000;
		1116: Delta = 46'sb1101111111111111111111110000000000000000000000;
		10002: Delta = 46'sb0100000000000000000000010000000000000000000000;
		2756: Delta = 46'sb1100000000000000000000010000000000000000000000;
		15857: Delta = 46'sb0011111111111111111111110000000000000000000000;
		8611: Delta = 46'sb1011111111111111111111110000000000000000000000;
		1048: Delta = 46'sb0000000000000000000001100000000000000000000000;
		17565: Delta = 46'sb1111111111111111111110100000000000000000000000;
		7951: Delta = 46'sb0000000000000000000010100000000000000000000000;
		10662: Delta = 46'sb1111111111111111111101100000000000000000000000;
		3144: Delta = 46'sb0000000000000000000100100000000000000000000000;
		3759: Delta = 46'sb1111111111111111111100100000000000000000000000;
		14854: Delta = 46'sb0000000000000000000011100000000000000000000000;
		15469: Delta = 46'sb1111111111111111111011100000000000000000000000;
		12143: Delta = 46'sb0000000000000000001000100000000000000000000000;
		13373: Delta = 46'sb1111111111111111111000100000000000000000000000;
		5240: Delta = 46'sb0000000000000000000111100000000000000000000000;
		6470: Delta = 46'sb1111111111111111110111100000000000000000000000;
		11528: Delta = 46'sb0000000000000000010000100000000000000000000000;
		13988: Delta = 46'sb1111111111111111110000100000000000000000000000;
		4625: Delta = 46'sb0000000000000000001111100000000000000000000000;
		7085: Delta = 46'sb1111111111111111101111100000000000000000000000;
		10298: Delta = 46'sb0000000000000000100000100000000000000000000000;
		15218: Delta = 46'sb1111111111111111100000100000000000000000000000;
		3395: Delta = 46'sb0000000000000000011111100000000000000000000000;
		8315: Delta = 46'sb1111111111111111011111100000000000000000000000;
		7838: Delta = 46'sb0000000000000001000000100000000000000000000000;
		17678: Delta = 46'sb1111111111111111000000100000000000000000000000;
		935: Delta = 46'sb0000000000000000111111100000000000000000000000;
		10775: Delta = 46'sb1111111111111110111111100000000000000000000000;
		2918: Delta = 46'sb0000000000000010000000100000000000000000000000;
		3985: Delta = 46'sb1111111111111110000000100000000000000000000000;
		14628: Delta = 46'sb0000000000000001111111100000000000000000000000;
		15695: Delta = 46'sb1111111111111101111111100000000000000000000000;
		11691: Delta = 46'sb0000000000000100000000100000000000000000000000;
		13825: Delta = 46'sb1111111111111100000000100000000000000000000000;
		4788: Delta = 46'sb0000000000000011111111100000000000000000000000;
		6922: Delta = 46'sb1111111111111011111111100000000000000000000000;
		10624: Delta = 46'sb0000000000001000000000100000000000000000000000;
		14892: Delta = 46'sb1111111111111000000000100000000000000000000000;
		3721: Delta = 46'sb0000000000000111111111100000000000000000000000;
		7989: Delta = 46'sb1111111111110111111111100000000000000000000000;
		8490: Delta = 46'sb0000000000010000000000100000000000000000000000;
		17026: Delta = 46'sb1111111111110000000000100000000000000000000000;
		1587: Delta = 46'sb0000000000001111111111100000000000000000000000;
		10123: Delta = 46'sb1111111111101111111111100000000000000000000000;
		4222: Delta = 46'sb0000000000100000000000100000000000000000000000;
		2681: Delta = 46'sb1111111111100000000000100000000000000000000000;
		15932: Delta = 46'sb0000000000011111111111100000000000000000000000;
		14391: Delta = 46'sb1111111111011111111111100000000000000000000000;
		14299: Delta = 46'sb0000000001000000000000100000000000000000000000;
		11217: Delta = 46'sb1111111111000000000000100000000000000000000000;
		7396: Delta = 46'sb0000000000111111111111100000000000000000000000;
		4314: Delta = 46'sb1111111110111111111111100000000000000000000000;
		15840: Delta = 46'sb0000000010000000000000100000000000000000000000;
		9676: Delta = 46'sb1111111110000000000000100000000000000000000000;
		8937: Delta = 46'sb0000000001111111111111100000000000000000000000;
		2773: Delta = 46'sb1111111101111111111111100000000000000000000000;
		309: Delta = 46'sb0000000100000000000000100000000000000000000000;
		6594: Delta = 46'sb1111111100000000000000100000000000000000000000;
		12019: Delta = 46'sb0000000011111111111111100000000000000000000000;
		18304: Delta = 46'sb1111111011111111111111100000000000000000000000;
		6473: Delta = 46'sb0000001000000000000000100000000000000000000000;
		430: Delta = 46'sb1111111000000000000000100000000000000000000000;
		18183: Delta = 46'sb0000000111111111111111100000000000000000000000;
		12140: Delta = 46'sb1111110111111111111111100000000000000000000000;
		188: Delta = 46'sb0000010000000000000000100000000000000000000000;
		6715: Delta = 46'sb1111110000000000000000100000000000000000000000;
		11898: Delta = 46'sb0000001111111111111111100000000000000000000000;
		18425: Delta = 46'sb1111101111111111111111100000000000000000000000;
		6231: Delta = 46'sb0000100000000000000000100000000000000000000000;
		672: Delta = 46'sb1111100000000000000000100000000000000000000000;
		17941: Delta = 46'sb0000011111111111111111100000000000000000000000;
		12382: Delta = 46'sb1111011111111111111111100000000000000000000000;
		18317: Delta = 46'sb0001000000000000000000100000000000000000000000;
		7199: Delta = 46'sb1111000000000000000000100000000000000000000000;
		11414: Delta = 46'sb0000111111111111111111100000000000000000000000;
		296: Delta = 46'sb1110111111111111111111100000000000000000000000;
		5263: Delta = 46'sb0010000000000000000000100000000000000000000000;
		1640: Delta = 46'sb1110000000000000000000100000000000000000000000;
		16973: Delta = 46'sb0001111111111111111111100000000000000000000000;
		13350: Delta = 46'sb1101111111111111111111100000000000000000000000;
		16381: Delta = 46'sb0100000000000000000000100000000000000000000000;
		9135: Delta = 46'sb1100000000000000000000100000000000000000000000;
		9478: Delta = 46'sb0011111111111111111111100000000000000000000000;
		2232: Delta = 46'sb1011111111111111111111100000000000000000000000;
		2096: Delta = 46'sb0000000000000000000011000000000000000000000000;
		16517: Delta = 46'sb1111111111111111111101000000000000000000000000;
		15902: Delta = 46'sb0000000000000000000101000000000000000000000000;
		2711: Delta = 46'sb1111111111111111111011000000000000000000000000;
		6288: Delta = 46'sb0000000000000000001001000000000000000000000000;
		7518: Delta = 46'sb1111111111111111111001000000000000000000000000;
		11095: Delta = 46'sb0000000000000000000111000000000000000000000000;
		12325: Delta = 46'sb1111111111111111110111000000000000000000000000;
		5673: Delta = 46'sb0000000000000000010001000000000000000000000000;
		8133: Delta = 46'sb1111111111111111110001000000000000000000000000;
		10480: Delta = 46'sb0000000000000000001111000000000000000000000000;
		12940: Delta = 46'sb1111111111111111101111000000000000000000000000;
		4443: Delta = 46'sb0000000000000000100001000000000000000000000000;
		9363: Delta = 46'sb1111111111111111100001000000000000000000000000;
		9250: Delta = 46'sb0000000000000000011111000000000000000000000000;
		14170: Delta = 46'sb1111111111111111011111000000000000000000000000;
		1983: Delta = 46'sb0000000000000001000001000000000000000000000000;
		11823: Delta = 46'sb1111111111111111000001000000000000000000000000;
		6790: Delta = 46'sb0000000000000000111111000000000000000000000000;
		16630: Delta = 46'sb1111111111111110111111000000000000000000000000;
		15676: Delta = 46'sb0000000000000010000001000000000000000000000000;
		16743: Delta = 46'sb1111111111111110000001000000000000000000000000;
		1870: Delta = 46'sb0000000000000001111111000000000000000000000000;
		2937: Delta = 46'sb1111111111111101111111000000000000000000000000;
		5836: Delta = 46'sb0000000000000100000001000000000000000000000000;
		7970: Delta = 46'sb1111111111111100000001000000000000000000000000;
		10643: Delta = 46'sb0000000000000011111111000000000000000000000000;
		12777: Delta = 46'sb1111111111111011111111000000000000000000000000;
		4769: Delta = 46'sb0000000000001000000001000000000000000000000000;
		9037: Delta = 46'sb1111111111111000000001000000000000000000000000;
		9576: Delta = 46'sb0000000000000111111111000000000000000000000000;
		13844: Delta = 46'sb1111111111110111111111000000000000000000000000;
		2635: Delta = 46'sb0000000000010000000001000000000000000000000000;
		11171: Delta = 46'sb1111111111110000000001000000000000000000000000;
		7442: Delta = 46'sb0000000000001111111111000000000000000000000000;
		15978: Delta = 46'sb1111111111101111111111000000000000000000000000;
		16980: Delta = 46'sb0000000000100000000001000000000000000000000000;
		15439: Delta = 46'sb1111111111100000000001000000000000000000000000;
		3174: Delta = 46'sb0000000000011111111111000000000000000000000000;
		1633: Delta = 46'sb1111111111011111111111000000000000000000000000;
		8444: Delta = 46'sb0000000001000000000001000000000000000000000000;
		5362: Delta = 46'sb1111111111000000000001000000000000000000000000;
		13251: Delta = 46'sb0000000000111111111111000000000000000000000000;
		10169: Delta = 46'sb1111111110111111111111000000000000000000000000;
		9985: Delta = 46'sb0000000010000000000001000000000000000000000000;
		3821: Delta = 46'sb1111111110000000000001000000000000000000000000;
		14792: Delta = 46'sb0000000001111111111111000000000000000000000000;
		8628: Delta = 46'sb1111111101111111111111000000000000000000000000;
		13067: Delta = 46'sb0000000100000000000001000000000000000000000000;
		739: Delta = 46'sb1111111100000000000001000000000000000000000000;
		17874: Delta = 46'sb0000000011111111111111000000000000000000000000;
		5546: Delta = 46'sb1111111011111111111111000000000000000000000000;
		618: Delta = 46'sb0000001000000000000001000000000000000000000000;
		13188: Delta = 46'sb1111111000000000000001000000000000000000000000;
		5425: Delta = 46'sb0000000111111111111111000000000000000000000000;
		17995: Delta = 46'sb1111110111111111111111000000000000000000000000;
		12946: Delta = 46'sb0000010000000000000001000000000000000000000000;
		860: Delta = 46'sb1111110000000000000001000000000000000000000000;
		17753: Delta = 46'sb0000001111111111111111000000000000000000000000;
		5667: Delta = 46'sb1111101111111111111111000000000000000000000000;
		376: Delta = 46'sb0000100000000000000001000000000000000000000000;
		13430: Delta = 46'sb1111100000000000000001000000000000000000000000;
		5183: Delta = 46'sb0000011111111111111111000000000000000000000000;
		18237: Delta = 46'sb1111011111111111111111000000000000000000000000;
		12462: Delta = 46'sb0001000000000000000001000000000000000000000000;
		1344: Delta = 46'sb1111000000000000000001000000000000000000000000;
		17269: Delta = 46'sb0000111111111111111111000000000000000000000000;
		6151: Delta = 46'sb1110111111111111111111000000000000000000000000;
		18021: Delta = 46'sb0010000000000000000001000000000000000000000000;
		14398: Delta = 46'sb1110000000000000000001000000000000000000000000;
		4215: Delta = 46'sb0001111111111111111111000000000000000000000000;
		592: Delta = 46'sb1101111111111111111111000000000000000000000000;
		10526: Delta = 46'sb0100000000000000000001000000000000000000000000;
		3280: Delta = 46'sb1100000000000000000001000000000000000000000000;
		15333: Delta = 46'sb0011111111111111111111000000000000000000000000;
		8087: Delta = 46'sb1011111111111111111111000000000000000000000000;
		4192: Delta = 46'sb0000000000000000000110000000000000000000000000;
		14421: Delta = 46'sb1111111111111111111010000000000000000000000000;
		13191: Delta = 46'sb0000000000000000001010000000000000000000000000;
		5422: Delta = 46'sb1111111111111111110110000000000000000000000000;
		12576: Delta = 46'sb0000000000000000010010000000000000000000000000;
		15036: Delta = 46'sb1111111111111111110010000000000000000000000000;
		3577: Delta = 46'sb0000000000000000001110000000000000000000000000;
		6037: Delta = 46'sb1111111111111111101110000000000000000000000000;
		11346: Delta = 46'sb0000000000000000100010000000000000000000000000;
		16266: Delta = 46'sb1111111111111111100010000000000000000000000000;
		2347: Delta = 46'sb0000000000000000011110000000000000000000000000;
		7267: Delta = 46'sb1111111111111111011110000000000000000000000000;
		8886: Delta = 46'sb0000000000000001000010000000000000000000000000;
		113: Delta = 46'sb1111111111111111000010000000000000000000000000;
		18500: Delta = 46'sb0000000000000000111110000000000000000000000000;
		9727: Delta = 46'sb1111111111111110111110000000000000000000000000;
		3966: Delta = 46'sb0000000000000010000010000000000000000000000000;
		5033: Delta = 46'sb1111111111111110000010000000000000000000000000;
		13580: Delta = 46'sb0000000000000001111110000000000000000000000000;
		14647: Delta = 46'sb1111111111111101111110000000000000000000000000;
		12739: Delta = 46'sb0000000000000100000010000000000000000000000000;
		14873: Delta = 46'sb1111111111111100000010000000000000000000000000;
		3740: Delta = 46'sb0000000000000011111110000000000000000000000000;
		5874: Delta = 46'sb1111111111111011111110000000000000000000000000;
		11672: Delta = 46'sb0000000000001000000010000000000000000000000000;
		15940: Delta = 46'sb1111111111111000000010000000000000000000000000;
		2673: Delta = 46'sb0000000000000111111110000000000000000000000000;
		6941: Delta = 46'sb1111111111110111111110000000000000000000000000;
		9538: Delta = 46'sb0000000000010000000010000000000000000000000000;
		18074: Delta = 46'sb1111111111110000000010000000000000000000000000;
		539: Delta = 46'sb0000000000001111111110000000000000000000000000;
		9075: Delta = 46'sb1111111111101111111110000000000000000000000000;
		5270: Delta = 46'sb0000000000100000000010000000000000000000000000;
		3729: Delta = 46'sb1111111111100000000010000000000000000000000000;
		14884: Delta = 46'sb0000000000011111111110000000000000000000000000;
		13343: Delta = 46'sb1111111111011111111110000000000000000000000000;
		15347: Delta = 46'sb0000000001000000000010000000000000000000000000;
		12265: Delta = 46'sb1111111111000000000010000000000000000000000000;
		6348: Delta = 46'sb0000000000111111111110000000000000000000000000;
		3266: Delta = 46'sb1111111110111111111110000000000000000000000000;
		16888: Delta = 46'sb0000000010000000000010000000000000000000000000;
		10724: Delta = 46'sb1111111110000000000010000000000000000000000000;
		7889: Delta = 46'sb0000000001111111111110000000000000000000000000;
		1725: Delta = 46'sb1111111101111111111110000000000000000000000000;
		1357: Delta = 46'sb0000000100000000000010000000000000000000000000;
		7642: Delta = 46'sb1111111100000000000010000000000000000000000000;
		10971: Delta = 46'sb0000000011111111111110000000000000000000000000;
		17256: Delta = 46'sb1111111011111111111110000000000000000000000000;
		7521: Delta = 46'sb0000001000000000000010000000000000000000000000;
		1478: Delta = 46'sb1111111000000000000010000000000000000000000000;
		17135: Delta = 46'sb0000000111111111111110000000000000000000000000;
		11092: Delta = 46'sb1111110111111111111110000000000000000000000000;
		1236: Delta = 46'sb0000010000000000000010000000000000000000000000;
		7763: Delta = 46'sb1111110000000000000010000000000000000000000000;
		10850: Delta = 46'sb0000001111111111111110000000000000000000000000;
		17377: Delta = 46'sb1111101111111111111110000000000000000000000000;
		7279: Delta = 46'sb0000100000000000000010000000000000000000000000;
		1720: Delta = 46'sb1111100000000000000010000000000000000000000000;
		16893: Delta = 46'sb0000011111111111111110000000000000000000000000;
		11334: Delta = 46'sb1111011111111111111110000000000000000000000000;
		752: Delta = 46'sb0001000000000000000010000000000000000000000000;
		8247: Delta = 46'sb1111000000000000000010000000000000000000000000;
		10366: Delta = 46'sb0000111111111111111110000000000000000000000000;
		17861: Delta = 46'sb1110111111111111111110000000000000000000000000;
		6311: Delta = 46'sb0010000000000000000010000000000000000000000000;
		2688: Delta = 46'sb1110000000000000000010000000000000000000000000;
		15925: Delta = 46'sb0001111111111111111110000000000000000000000000;
		12302: Delta = 46'sb1101111111111111111110000000000000000000000000;
		17429: Delta = 46'sb0100000000000000000010000000000000000000000000;
		10183: Delta = 46'sb1100000000000000000010000000000000000000000000;
		8430: Delta = 46'sb0011111111111111111110000000000000000000000000;
		1184: Delta = 46'sb1011111111111111111110000000000000000000000000;
		8384: Delta = 46'sb0000000000000000001100000000000000000000000000;
		10229: Delta = 46'sb1111111111111111110100000000000000000000000000;
		7769: Delta = 46'sb0000000000000000010100000000000000000000000000;
		10844: Delta = 46'sb1111111111111111101100000000000000000000000000;
		6539: Delta = 46'sb0000000000000000100100000000000000000000000000;
		11459: Delta = 46'sb1111111111111111100100000000000000000000000000;
		7154: Delta = 46'sb0000000000000000011100000000000000000000000000;
		12074: Delta = 46'sb1111111111111111011100000000000000000000000000;
		4079: Delta = 46'sb0000000000000001000100000000000000000000000000;
		13919: Delta = 46'sb1111111111111111000100000000000000000000000000;
		4694: Delta = 46'sb0000000000000000111100000000000000000000000000;
		14534: Delta = 46'sb1111111111111110111100000000000000000000000000;
		17772: Delta = 46'sb0000000000000010000100000000000000000000000000;
		226: Delta = 46'sb1111111111111110000100000000000000000000000000;
		18387: Delta = 46'sb0000000000000001111100000000000000000000000000;
		841: Delta = 46'sb1111111111111101111100000000000000000000000000;
		7932: Delta = 46'sb0000000000000100000100000000000000000000000000;
		10066: Delta = 46'sb1111111111111100000100000000000000000000000000;
		8547: Delta = 46'sb0000000000000011111100000000000000000000000000;
		10681: Delta = 46'sb1111111111111011111100000000000000000000000000;
		6865: Delta = 46'sb0000000000001000000100000000000000000000000000;
		11133: Delta = 46'sb1111111111111000000100000000000000000000000000;
		7480: Delta = 46'sb0000000000000111111100000000000000000000000000;
		11748: Delta = 46'sb1111111111110111111100000000000000000000000000;
		4731: Delta = 46'sb0000000000010000000100000000000000000000000000;
		13267: Delta = 46'sb1111111111110000000100000000000000000000000000;
		5346: Delta = 46'sb0000000000001111111100000000000000000000000000;
		13882: Delta = 46'sb1111111111101111111100000000000000000000000000;
		463: Delta = 46'sb0000000000100000000100000000000000000000000000;
		17535: Delta = 46'sb1111111111100000000100000000000000000000000000;
		1078: Delta = 46'sb0000000000011111111100000000000000000000000000;
		18150: Delta = 46'sb1111111111011111111100000000000000000000000000;
		10540: Delta = 46'sb0000000001000000000100000000000000000000000000;
		7458: Delta = 46'sb1111111111000000000100000000000000000000000000;
		11155: Delta = 46'sb0000000000111111111100000000000000000000000000;
		8073: Delta = 46'sb1111111110111111111100000000000000000000000000;
		12081: Delta = 46'sb0000000010000000000100000000000000000000000000;
		5917: Delta = 46'sb1111111110000000000100000000000000000000000000;
		12696: Delta = 46'sb0000000001111111111100000000000000000000000000;
		6532: Delta = 46'sb1111111101111111111100000000000000000000000000;
		15163: Delta = 46'sb0000000100000000000100000000000000000000000000;
		2835: Delta = 46'sb1111111100000000000100000000000000000000000000;
		15778: Delta = 46'sb0000000011111111111100000000000000000000000000;
		3450: Delta = 46'sb1111111011111111111100000000000000000000000000;
		2714: Delta = 46'sb0000001000000000000100000000000000000000000000;
		15284: Delta = 46'sb1111111000000000000100000000000000000000000000;
		3329: Delta = 46'sb0000000111111111111100000000000000000000000000;
		15899: Delta = 46'sb1111110111111111111100000000000000000000000000;
		15042: Delta = 46'sb0000010000000000000100000000000000000000000000;
		2956: Delta = 46'sb1111110000000000000100000000000000000000000000;
		15657: Delta = 46'sb0000001111111111111100000000000000000000000000;
		3571: Delta = 46'sb1111101111111111111100000000000000000000000000;
		2472: Delta = 46'sb0000100000000000000100000000000000000000000000;
		15526: Delta = 46'sb1111100000000000000100000000000000000000000000;
		3087: Delta = 46'sb0000011111111111111100000000000000000000000000;
		16141: Delta = 46'sb1111011111111111111100000000000000000000000000;
		14558: Delta = 46'sb0001000000000000000100000000000000000000000000;
		3440: Delta = 46'sb1111000000000000000100000000000000000000000000;
		15173: Delta = 46'sb0000111111111111111100000000000000000000000000;
		4055: Delta = 46'sb1110111111111111111100000000000000000000000000;
		1504: Delta = 46'sb0010000000000000000100000000000000000000000000;
		16494: Delta = 46'sb1110000000000000000100000000000000000000000000;
		2119: Delta = 46'sb0001111111111111111100000000000000000000000000;
		17109: Delta = 46'sb1101111111111111111100000000000000000000000000;
		12622: Delta = 46'sb0100000000000000000100000000000000000000000000;
		5376: Delta = 46'sb1100000000000000000100000000000000000000000000;
		13237: Delta = 46'sb0011111111111111111100000000000000000000000000;
		5991: Delta = 46'sb1011111111111111111100000000000000000000000000;
		16768: Delta = 46'sb0000000000000000011000000000000000000000000000;
		1845: Delta = 46'sb1111111111111111101000000000000000000000000000;
		15538: Delta = 46'sb0000000000000000101000000000000000000000000000;
		3075: Delta = 46'sb1111111111111111011000000000000000000000000000;
		13078: Delta = 46'sb0000000000000001001000000000000000000000000000;
		4305: Delta = 46'sb1111111111111111001000000000000000000000000000;
		14308: Delta = 46'sb0000000000000000111000000000000000000000000000;
		5535: Delta = 46'sb1111111111111110111000000000000000000000000000;
		8158: Delta = 46'sb0000000000000010001000000000000000000000000000;
		9225: Delta = 46'sb1111111111111110001000000000000000000000000000;
		9388: Delta = 46'sb0000000000000001111000000000000000000000000000;
		10455: Delta = 46'sb1111111111111101111000000000000000000000000000;
		16931: Delta = 46'sb0000000000000100001000000000000000000000000000;
		452: Delta = 46'sb1111111111111100001000000000000000000000000000;
		18161: Delta = 46'sb0000000000000011111000000000000000000000000000;
		1682: Delta = 46'sb1111111111111011111000000000000000000000000000;
		15864: Delta = 46'sb0000000000001000001000000000000000000000000000;
		1519: Delta = 46'sb1111111111111000001000000000000000000000000000;
		17094: Delta = 46'sb0000000000000111111000000000000000000000000000;
		2749: Delta = 46'sb1111111111110111111000000000000000000000000000;
		13730: Delta = 46'sb0000000000010000001000000000000000000000000000;
		3653: Delta = 46'sb1111111111110000001000000000000000000000000000;
		14960: Delta = 46'sb0000000000001111111000000000000000000000000000;
		4883: Delta = 46'sb1111111111101111111000000000000000000000000000;
		9462: Delta = 46'sb0000000000100000001000000000000000000000000000;
		7921: Delta = 46'sb1111111111100000001000000000000000000000000000;
		10692: Delta = 46'sb0000000000011111111000000000000000000000000000;
		9151: Delta = 46'sb1111111111011111111000000000000000000000000000;
		926: Delta = 46'sb0000000001000000001000000000000000000000000000;
		16457: Delta = 46'sb1111111111000000001000000000000000000000000000;
		2156: Delta = 46'sb0000000000111111111000000000000000000000000000;
		17687: Delta = 46'sb1111111110111111111000000000000000000000000000;
		2467: Delta = 46'sb0000000010000000001000000000000000000000000000;
		14916: Delta = 46'sb1111111110000000001000000000000000000000000000;
		3697: Delta = 46'sb0000000001111111111000000000000000000000000000;
		16146: Delta = 46'sb1111111101111111111000000000000000000000000000;
		5549: Delta = 46'sb0000000100000000001000000000000000000000000000;
		11834: Delta = 46'sb1111111100000000001000000000000000000000000000;
		6779: Delta = 46'sb0000000011111111111000000000000000000000000000;
		13064: Delta = 46'sb1111111011111111111000000000000000000000000000;
		11713: Delta = 46'sb0000001000000000001000000000000000000000000000;
		5670: Delta = 46'sb1111111000000000001000000000000000000000000000;
		12943: Delta = 46'sb0000000111111111111000000000000000000000000000;
		6900: Delta = 46'sb1111110111111111111000000000000000000000000000;
		5428: Delta = 46'sb0000010000000000001000000000000000000000000000;
		11955: Delta = 46'sb1111110000000000001000000000000000000000000000;
		6658: Delta = 46'sb0000001111111111111000000000000000000000000000;
		13185: Delta = 46'sb1111101111111111111000000000000000000000000000;
		11471: Delta = 46'sb0000100000000000001000000000000000000000000000;
		5912: Delta = 46'sb1111100000000000001000000000000000000000000000;
		12701: Delta = 46'sb0000011111111111111000000000000000000000000000;
		7142: Delta = 46'sb1111011111111111111000000000000000000000000000;
		4944: Delta = 46'sb0001000000000000001000000000000000000000000000;
		12439: Delta = 46'sb1111000000000000001000000000000000000000000000;
		6174: Delta = 46'sb0000111111111111111000000000000000000000000000;
		13669: Delta = 46'sb1110111111111111111000000000000000000000000000;
		10503: Delta = 46'sb0010000000000000001000000000000000000000000000;
		6880: Delta = 46'sb1110000000000000001000000000000000000000000000;
		11733: Delta = 46'sb0001111111111111111000000000000000000000000000;
		8110: Delta = 46'sb1101111111111111111000000000000000000000000000;
		3008: Delta = 46'sb0100000000000000001000000000000000000000000000;
		14375: Delta = 46'sb1100000000000000001000000000000000000000000000;
		4238: Delta = 46'sb0011111111111111111000000000000000000000000000;
		15605: Delta = 46'sb1011111111111111111000000000000000000000000000;
		14923: Delta = 46'sb0000000000000000110000000000000000000000000000;
		3690: Delta = 46'sb1111111111111111010000000000000000000000000000;
		12463: Delta = 46'sb0000000000000001010000000000000000000000000000;
		6150: Delta = 46'sb1111111111111110110000000000000000000000000000;
		7543: Delta = 46'sb0000000000000010010000000000000000000000000000;
		8610: Delta = 46'sb1111111111111110010000000000000000000000000000;
		10003: Delta = 46'sb0000000000000001110000000000000000000000000000;
		11070: Delta = 46'sb1111111111111101110000000000000000000000000000;
		16316: Delta = 46'sb0000000000000100010000000000000000000000000000;
		18450: Delta = 46'sb1111111111111100010000000000000000000000000000;
		163: Delta = 46'sb0000000000000011110000000000000000000000000000;
		2297: Delta = 46'sb1111111111111011110000000000000000000000000000;
		15249: Delta = 46'sb0000000000001000010000000000000000000000000000;
		904: Delta = 46'sb1111111111111000010000000000000000000000000000;
		17709: Delta = 46'sb0000000000000111110000000000000000000000000000;
		3364: Delta = 46'sb1111111111110111110000000000000000000000000000;
		13115: Delta = 46'sb0000000000010000010000000000000000000000000000;
		3038: Delta = 46'sb1111111111110000010000000000000000000000000000;
		15575: Delta = 46'sb0000000000001111110000000000000000000000000000;
		5498: Delta = 46'sb1111111111101111110000000000000000000000000000;
		8847: Delta = 46'sb0000000000100000010000000000000000000000000000;
		7306: Delta = 46'sb1111111111100000010000000000000000000000000000;
		11307: Delta = 46'sb0000000000011111110000000000000000000000000000;
		9766: Delta = 46'sb1111111111011111110000000000000000000000000000;
		311: Delta = 46'sb0000000001000000010000000000000000000000000000;
		15842: Delta = 46'sb1111111111000000010000000000000000000000000000;
		2771: Delta = 46'sb0000000000111111110000000000000000000000000000;
		18302: Delta = 46'sb1111111110111111110000000000000000000000000000;
		1852: Delta = 46'sb0000000010000000010000000000000000000000000000;
		14301: Delta = 46'sb1111111110000000010000000000000000000000000000;
		4312: Delta = 46'sb0000000001111111110000000000000000000000000000;
		16761: Delta = 46'sb1111111101111111110000000000000000000000000000;
		4934: Delta = 46'sb0000000100000000010000000000000000000000000000;
		11219: Delta = 46'sb1111111100000000010000000000000000000000000000;
		7394: Delta = 46'sb0000000011111111110000000000000000000000000000;
		13679: Delta = 46'sb1111111011111111110000000000000000000000000000;
		11098: Delta = 46'sb0000001000000000010000000000000000000000000000;
		5055: Delta = 46'sb1111111000000000010000000000000000000000000000;
		13558: Delta = 46'sb0000000111111111110000000000000000000000000000;
		7515: Delta = 46'sb1111110111111111110000000000000000000000000000;
		4813: Delta = 46'sb0000010000000000010000000000000000000000000000;
		11340: Delta = 46'sb1111110000000000010000000000000000000000000000;
		7273: Delta = 46'sb0000001111111111110000000000000000000000000000;
		13800: Delta = 46'sb1111101111111111110000000000000000000000000000;
		10856: Delta = 46'sb0000100000000000010000000000000000000000000000;
		5297: Delta = 46'sb1111100000000000010000000000000000000000000000;
		13316: Delta = 46'sb0000011111111111110000000000000000000000000000;
		7757: Delta = 46'sb1111011111111111110000000000000000000000000000;
		4329: Delta = 46'sb0001000000000000010000000000000000000000000000;
		11824: Delta = 46'sb1111000000000000010000000000000000000000000000;
		6789: Delta = 46'sb0000111111111111110000000000000000000000000000;
		14284: Delta = 46'sb1110111111111111110000000000000000000000000000;
		9888: Delta = 46'sb0010000000000000010000000000000000000000000000;
		6265: Delta = 46'sb1110000000000000010000000000000000000000000000;
		12348: Delta = 46'sb0001111111111111110000000000000000000000000000;
		8725: Delta = 46'sb1101111111111111110000000000000000000000000000;
		2393: Delta = 46'sb0100000000000000010000000000000000000000000000;
		13760: Delta = 46'sb1100000000000000010000000000000000000000000000;
		4853: Delta = 46'sb0011111111111111110000000000000000000000000000;
		16220: Delta = 46'sb1011111111111111110000000000000000000000000000;
		11233: Delta = 46'sb0000000000000001100000000000000000000000000000;
		7380: Delta = 46'sb1111111111111110100000000000000000000000000000;
		6313: Delta = 46'sb0000000000000010100000000000000000000000000000;
		12300: Delta = 46'sb1111111111111101100000000000000000000000000000;
		15086: Delta = 46'sb0000000000000100100000000000000000000000000000;
		17220: Delta = 46'sb1111111111111100100000000000000000000000000000;
		1393: Delta = 46'sb0000000000000011100000000000000000000000000000;
		3527: Delta = 46'sb1111111111111011100000000000000000000000000000;
		14019: Delta = 46'sb0000000000001000100000000000000000000000000000;
		18287: Delta = 46'sb1111111111111000100000000000000000000000000000;
		326: Delta = 46'sb0000000000000111100000000000000000000000000000;
		4594: Delta = 46'sb1111111111110111100000000000000000000000000000;
		11885: Delta = 46'sb0000000000010000100000000000000000000000000000;
		1808: Delta = 46'sb1111111111110000100000000000000000000000000000;
		16805: Delta = 46'sb0000000000001111100000000000000000000000000000;
		6728: Delta = 46'sb1111111111101111100000000000000000000000000000;
		7617: Delta = 46'sb0000000000100000100000000000000000000000000000;
		6076: Delta = 46'sb1111111111100000100000000000000000000000000000;
		12537: Delta = 46'sb0000000000011111100000000000000000000000000000;
		10996: Delta = 46'sb1111111111011111100000000000000000000000000000;
		17694: Delta = 46'sb0000000001000000100000000000000000000000000000;
		14612: Delta = 46'sb1111111111000000100000000000000000000000000000;
		4001: Delta = 46'sb0000000000111111100000000000000000000000000000;
		919: Delta = 46'sb1111111110111111100000000000000000000000000000;
		622: Delta = 46'sb0000000010000000100000000000000000000000000000;
		13071: Delta = 46'sb1111111110000000100000000000000000000000000000;
		5542: Delta = 46'sb0000000001111111100000000000000000000000000000;
		17991: Delta = 46'sb1111111101111111100000000000000000000000000000;
		3704: Delta = 46'sb0000000100000000100000000000000000000000000000;
		9989: Delta = 46'sb1111111100000000100000000000000000000000000000;
		8624: Delta = 46'sb0000000011111111100000000000000000000000000000;
		14909: Delta = 46'sb1111111011111111100000000000000000000000000000;
		9868: Delta = 46'sb0000001000000000100000000000000000000000000000;
		3825: Delta = 46'sb1111111000000000100000000000000000000000000000;
		14788: Delta = 46'sb0000000111111111100000000000000000000000000000;
		8745: Delta = 46'sb1111110111111111100000000000000000000000000000;
		3583: Delta = 46'sb0000010000000000100000000000000000000000000000;
		10110: Delta = 46'sb1111110000000000100000000000000000000000000000;
		8503: Delta = 46'sb0000001111111111100000000000000000000000000000;
		15030: Delta = 46'sb1111101111111111100000000000000000000000000000;
		9626: Delta = 46'sb0000100000000000100000000000000000000000000000;
		4067: Delta = 46'sb1111100000000000100000000000000000000000000000;
		14546: Delta = 46'sb0000011111111111100000000000000000000000000000;
		8987: Delta = 46'sb1111011111111111100000000000000000000000000000;
		3099: Delta = 46'sb0001000000000000100000000000000000000000000000;
		10594: Delta = 46'sb1111000000000000100000000000000000000000000000;
		8019: Delta = 46'sb0000111111111111100000000000000000000000000000;
		15514: Delta = 46'sb1110111111111111100000000000000000000000000000;
		8658: Delta = 46'sb0010000000000000100000000000000000000000000000;
		5035: Delta = 46'sb1110000000000000100000000000000000000000000000;
		13578: Delta = 46'sb0001111111111111100000000000000000000000000000;
		9955: Delta = 46'sb1101111111111111100000000000000000000000000000;
		1163: Delta = 46'sb0100000000000000100000000000000000000000000000;
		12530: Delta = 46'sb1100000000000000100000000000000000000000000000;
		6083: Delta = 46'sb0011111111111111100000000000000000000000000000;
		17450: Delta = 46'sb1011111111111111100000000000000000000000000000;
		3853: Delta = 46'sb0000000000000011000000000000000000000000000000;
		14760: Delta = 46'sb1111111111111101000000000000000000000000000000;
		12626: Delta = 46'sb0000000000000101000000000000000000000000000000;
		5987: Delta = 46'sb1111111111111011000000000000000000000000000000;
		11559: Delta = 46'sb0000000000001001000000000000000000000000000000;
		15827: Delta = 46'sb1111111111111001000000000000000000000000000000;
		2786: Delta = 46'sb0000000000000111000000000000000000000000000000;
		7054: Delta = 46'sb1111111111110111000000000000000000000000000000;
		9425: Delta = 46'sb0000000000010001000000000000000000000000000000;
		17961: Delta = 46'sb1111111111110001000000000000000000000000000000;
		652: Delta = 46'sb0000000000001111000000000000000000000000000000;
		9188: Delta = 46'sb1111111111101111000000000000000000000000000000;
		5157: Delta = 46'sb0000000000100001000000000000000000000000000000;
		3616: Delta = 46'sb1111111111100001000000000000000000000000000000;
		14997: Delta = 46'sb0000000000011111000000000000000000000000000000;
		13456: Delta = 46'sb1111111111011111000000000000000000000000000000;
		15234: Delta = 46'sb0000000001000001000000000000000000000000000000;
		12152: Delta = 46'sb1111111111000001000000000000000000000000000000;
		6461: Delta = 46'sb0000000000111111000000000000000000000000000000;
		3379: Delta = 46'sb1111111110111111000000000000000000000000000000;
		16775: Delta = 46'sb0000000010000001000000000000000000000000000000;
		10611: Delta = 46'sb1111111110000001000000000000000000000000000000;
		8002: Delta = 46'sb0000000001111111000000000000000000000000000000;
		1838: Delta = 46'sb1111111101111111000000000000000000000000000000;
		1244: Delta = 46'sb0000000100000001000000000000000000000000000000;
		7529: Delta = 46'sb1111111100000001000000000000000000000000000000;
		11084: Delta = 46'sb0000000011111111000000000000000000000000000000;
		17369: Delta = 46'sb1111111011111111000000000000000000000000000000;
		7408: Delta = 46'sb0000001000000001000000000000000000000000000000;
		1365: Delta = 46'sb1111111000000001000000000000000000000000000000;
		17248: Delta = 46'sb0000000111111111000000000000000000000000000000;
		11205: Delta = 46'sb1111110111111111000000000000000000000000000000;
		1123: Delta = 46'sb0000010000000001000000000000000000000000000000;
		7650: Delta = 46'sb1111110000000001000000000000000000000000000000;
		10963: Delta = 46'sb0000001111111111000000000000000000000000000000;
		17490: Delta = 46'sb1111101111111111000000000000000000000000000000;
		7166: Delta = 46'sb0000100000000001000000000000000000000000000000;
		1607: Delta = 46'sb1111100000000001000000000000000000000000000000;
		17006: Delta = 46'sb0000011111111111000000000000000000000000000000;
		11447: Delta = 46'sb1111011111111111000000000000000000000000000000;
		639: Delta = 46'sb0001000000000001000000000000000000000000000000;
		8134: Delta = 46'sb1111000000000001000000000000000000000000000000;
		10479: Delta = 46'sb0000111111111111000000000000000000000000000000;
		17974: Delta = 46'sb1110111111111111000000000000000000000000000000;
		6198: Delta = 46'sb0010000000000001000000000000000000000000000000;
		2575: Delta = 46'sb1110000000000001000000000000000000000000000000;
		16038: Delta = 46'sb0001111111111111000000000000000000000000000000;
		12415: Delta = 46'sb1101111111111111000000000000000000000000000000;
		17316: Delta = 46'sb0100000000000001000000000000000000000000000000;
		10070: Delta = 46'sb1100000000000001000000000000000000000000000000;
		8543: Delta = 46'sb0011111111111111000000000000000000000000000000;
		1297: Delta = 46'sb1011111111111111000000000000000000000000000000;
		7706: Delta = 46'sb0000000000000110000000000000000000000000000000;
		10907: Delta = 46'sb1111111111111010000000000000000000000000000000;
		6639: Delta = 46'sb0000000000001010000000000000000000000000000000;
		11974: Delta = 46'sb1111111111110110000000000000000000000000000000;
		4505: Delta = 46'sb0000000000010010000000000000000000000000000000;
		13041: Delta = 46'sb1111111111110010000000000000000000000000000000;
		5572: Delta = 46'sb0000000000001110000000000000000000000000000000;
		14108: Delta = 46'sb1111111111101110000000000000000000000000000000;
		237: Delta = 46'sb0000000000100010000000000000000000000000000000;
		17309: Delta = 46'sb1111111111100010000000000000000000000000000000;
		1304: Delta = 46'sb0000000000011110000000000000000000000000000000;
		18376: Delta = 46'sb1111111111011110000000000000000000000000000000;
		10314: Delta = 46'sb0000000001000010000000000000000000000000000000;
		7232: Delta = 46'sb1111111111000010000000000000000000000000000000;
		11381: Delta = 46'sb0000000000111110000000000000000000000000000000;
		8299: Delta = 46'sb1111111110111110000000000000000000000000000000;
		11855: Delta = 46'sb0000000010000010000000000000000000000000000000;
		5691: Delta = 46'sb1111111110000010000000000000000000000000000000;
		12922: Delta = 46'sb0000000001111110000000000000000000000000000000;
		6758: Delta = 46'sb1111111101111110000000000000000000000000000000;
		14937: Delta = 46'sb0000000100000010000000000000000000000000000000;
		2609: Delta = 46'sb1111111100000010000000000000000000000000000000;
		16004: Delta = 46'sb0000000011111110000000000000000000000000000000;
		3676: Delta = 46'sb1111111011111110000000000000000000000000000000;
		2488: Delta = 46'sb0000001000000010000000000000000000000000000000;
		15058: Delta = 46'sb1111111000000010000000000000000000000000000000;
		3555: Delta = 46'sb0000000111111110000000000000000000000000000000;
		16125: Delta = 46'sb1111110111111110000000000000000000000000000000;
		14816: Delta = 46'sb0000010000000010000000000000000000000000000000;
		2730: Delta = 46'sb1111110000000010000000000000000000000000000000;
		15883: Delta = 46'sb0000001111111110000000000000000000000000000000;
		3797: Delta = 46'sb1111101111111110000000000000000000000000000000;
		2246: Delta = 46'sb0000100000000010000000000000000000000000000000;
		15300: Delta = 46'sb1111100000000010000000000000000000000000000000;
		3313: Delta = 46'sb0000011111111110000000000000000000000000000000;
		16367: Delta = 46'sb1111011111111110000000000000000000000000000000;
		14332: Delta = 46'sb0001000000000010000000000000000000000000000000;
		3214: Delta = 46'sb1111000000000010000000000000000000000000000000;
		15399: Delta = 46'sb0000111111111110000000000000000000000000000000;
		4281: Delta = 46'sb1110111111111110000000000000000000000000000000;
		1278: Delta = 46'sb0010000000000010000000000000000000000000000000;
		16268: Delta = 46'sb1110000000000010000000000000000000000000000000;
		2345: Delta = 46'sb0001111111111110000000000000000000000000000000;
		17335: Delta = 46'sb1101111111111110000000000000000000000000000000;
		12396: Delta = 46'sb0100000000000010000000000000000000000000000000;
		5150: Delta = 46'sb1100000000000010000000000000000000000000000000;
		13463: Delta = 46'sb0011111111111110000000000000000000000000000000;
		6217: Delta = 46'sb1011111111111110000000000000000000000000000000;
		15412: Delta = 46'sb0000000000001100000000000000000000000000000000;
		3201: Delta = 46'sb1111111111110100000000000000000000000000000000;
		13278: Delta = 46'sb0000000000010100000000000000000000000000000000;
		5335: Delta = 46'sb1111111111101100000000000000000000000000000000;
		9010: Delta = 46'sb0000000000100100000000000000000000000000000000;
		7469: Delta = 46'sb1111111111100100000000000000000000000000000000;
		11144: Delta = 46'sb0000000000011100000000000000000000000000000000;
		9603: Delta = 46'sb1111111111011100000000000000000000000000000000;
		474: Delta = 46'sb0000000001000100000000000000000000000000000000;
		16005: Delta = 46'sb1111111111000100000000000000000000000000000000;
		2608: Delta = 46'sb0000000000111100000000000000000000000000000000;
		18139: Delta = 46'sb1111111110111100000000000000000000000000000000;
		2015: Delta = 46'sb0000000010000100000000000000000000000000000000;
		14464: Delta = 46'sb1111111110000100000000000000000000000000000000;
		4149: Delta = 46'sb0000000001111100000000000000000000000000000000;
		16598: Delta = 46'sb1111111101111100000000000000000000000000000000;
		5097: Delta = 46'sb0000000100000100000000000000000000000000000000;
		11382: Delta = 46'sb1111111100000100000000000000000000000000000000;
		7231: Delta = 46'sb0000000011111100000000000000000000000000000000;
		13516: Delta = 46'sb1111111011111100000000000000000000000000000000;
		11261: Delta = 46'sb0000001000000100000000000000000000000000000000;
		5218: Delta = 46'sb1111111000000100000000000000000000000000000000;
		13395: Delta = 46'sb0000000111111100000000000000000000000000000000;
		7352: Delta = 46'sb1111110111111100000000000000000000000000000000;
		4976: Delta = 46'sb0000010000000100000000000000000000000000000000;
		11503: Delta = 46'sb1111110000000100000000000000000000000000000000;
		7110: Delta = 46'sb0000001111111100000000000000000000000000000000;
		13637: Delta = 46'sb1111101111111100000000000000000000000000000000;
		11019: Delta = 46'sb0000100000000100000000000000000000000000000000;
		5460: Delta = 46'sb1111100000000100000000000000000000000000000000;
		13153: Delta = 46'sb0000011111111100000000000000000000000000000000;
		7594: Delta = 46'sb1111011111111100000000000000000000000000000000;
		4492: Delta = 46'sb0001000000000100000000000000000000000000000000;
		11987: Delta = 46'sb1111000000000100000000000000000000000000000000;
		6626: Delta = 46'sb0000111111111100000000000000000000000000000000;
		14121: Delta = 46'sb1110111111111100000000000000000000000000000000;
		10051: Delta = 46'sb0010000000000100000000000000000000000000000000;
		6428: Delta = 46'sb1110000000000100000000000000000000000000000000;
		12185: Delta = 46'sb0001111111111100000000000000000000000000000000;
		8562: Delta = 46'sb1101111111111100000000000000000000000000000000;
		2556: Delta = 46'sb0100000000000100000000000000000000000000000000;
		13923: Delta = 46'sb1100000000000100000000000000000000000000000000;
		4690: Delta = 46'sb0011111111111100000000000000000000000000000000;
		16057: Delta = 46'sb1011111111111100000000000000000000000000000000;
		12211: Delta = 46'sb0000000000011000000000000000000000000000000000;
		6402: Delta = 46'sb1111111111101000000000000000000000000000000000;
		7943: Delta = 46'sb0000000000101000000000000000000000000000000000;
		10670: Delta = 46'sb1111111111011000000000000000000000000000000000;
		18020: Delta = 46'sb0000000001001000000000000000000000000000000000;
		14938: Delta = 46'sb1111111111001000000000000000000000000000000000;
		3675: Delta = 46'sb0000000000111000000000000000000000000000000000;
		593: Delta = 46'sb1111111110111000000000000000000000000000000000;
		948: Delta = 46'sb0000000010001000000000000000000000000000000000;
		13397: Delta = 46'sb1111111110001000000000000000000000000000000000;
		5216: Delta = 46'sb0000000001111000000000000000000000000000000000;
		17665: Delta = 46'sb1111111101111000000000000000000000000000000000;
		4030: Delta = 46'sb0000000100001000000000000000000000000000000000;
		10315: Delta = 46'sb1111111100001000000000000000000000000000000000;
		8298: Delta = 46'sb0000000011111000000000000000000000000000000000;
		14583: Delta = 46'sb1111111011111000000000000000000000000000000000;
		10194: Delta = 46'sb0000001000001000000000000000000000000000000000;
		4151: Delta = 46'sb1111111000001000000000000000000000000000000000;
		14462: Delta = 46'sb0000000111111000000000000000000000000000000000;
		8419: Delta = 46'sb1111110111111000000000000000000000000000000000;
		3909: Delta = 46'sb0000010000001000000000000000000000000000000000;
		10436: Delta = 46'sb1111110000001000000000000000000000000000000000;
		8177: Delta = 46'sb0000001111111000000000000000000000000000000000;
		14704: Delta = 46'sb1111101111111000000000000000000000000000000000;
		9952: Delta = 46'sb0000100000001000000000000000000000000000000000;
		4393: Delta = 46'sb1111100000001000000000000000000000000000000000;
		14220: Delta = 46'sb0000011111111000000000000000000000000000000000;
		8661: Delta = 46'sb1111011111111000000000000000000000000000000000;
		3425: Delta = 46'sb0001000000001000000000000000000000000000000000;
		10920: Delta = 46'sb1111000000001000000000000000000000000000000000;
		7693: Delta = 46'sb0000111111111000000000000000000000000000000000;
		15188: Delta = 46'sb1110111111111000000000000000000000000000000000;
		8984: Delta = 46'sb0010000000001000000000000000000000000000000000;
		5361: Delta = 46'sb1110000000001000000000000000000000000000000000;
		13252: Delta = 46'sb0001111111111000000000000000000000000000000000;
		9629: Delta = 46'sb1101111111111000000000000000000000000000000000;
		1489: Delta = 46'sb0100000000001000000000000000000000000000000000;
		12856: Delta = 46'sb1100000000001000000000000000000000000000000000;
		5757: Delta = 46'sb0011111111111000000000000000000000000000000000;
		17124: Delta = 46'sb1011111111111000000000000000000000000000000000;
		5809: Delta = 46'sb0000000000110000000000000000000000000000000000;
		12804: Delta = 46'sb1111111111010000000000000000000000000000000000;
		15886: Delta = 46'sb0000000001010000000000000000000000000000000000;
		2727: Delta = 46'sb1111111110110000000000000000000000000000000000;
		17427: Delta = 46'sb0000000010010000000000000000000000000000000000;
		11263: Delta = 46'sb1111111110010000000000000000000000000000000000;
		7350: Delta = 46'sb0000000001110000000000000000000000000000000000;
		1186: Delta = 46'sb1111111101110000000000000000000000000000000000;
		1896: Delta = 46'sb0000000100010000000000000000000000000000000000;
		8181: Delta = 46'sb1111111100010000000000000000000000000000000000;
		10432: Delta = 46'sb0000000011110000000000000000000000000000000000;
		16717: Delta = 46'sb1111111011110000000000000000000000000000000000;
		8060: Delta = 46'sb0000001000010000000000000000000000000000000000;
		2017: Delta = 46'sb1111111000010000000000000000000000000000000000;
		16596: Delta = 46'sb0000000111110000000000000000000000000000000000;
		10553: Delta = 46'sb1111110111110000000000000000000000000000000000;
		1775: Delta = 46'sb0000010000010000000000000000000000000000000000;
		8302: Delta = 46'sb1111110000010000000000000000000000000000000000;
		10311: Delta = 46'sb0000001111110000000000000000000000000000000000;
		16838: Delta = 46'sb1111101111110000000000000000000000000000000000;
		7818: Delta = 46'sb0000100000010000000000000000000000000000000000;
		2259: Delta = 46'sb1111100000010000000000000000000000000000000000;
		16354: Delta = 46'sb0000011111110000000000000000000000000000000000;
		10795: Delta = 46'sb1111011111110000000000000000000000000000000000;
		1291: Delta = 46'sb0001000000010000000000000000000000000000000000;
		8786: Delta = 46'sb1111000000010000000000000000000000000000000000;
		9827: Delta = 46'sb0000111111110000000000000000000000000000000000;
		17322: Delta = 46'sb1110111111110000000000000000000000000000000000;
		6850: Delta = 46'sb0010000000010000000000000000000000000000000000;
		3227: Delta = 46'sb1110000000010000000000000000000000000000000000;
		15386: Delta = 46'sb0001111111110000000000000000000000000000000000;
		11763: Delta = 46'sb1101111111110000000000000000000000000000000000;
		17968: Delta = 46'sb0100000000010000000000000000000000000000000000;
		10722: Delta = 46'sb1100000000010000000000000000000000000000000000;
		7891: Delta = 46'sb0011111111110000000000000000000000000000000000;
		645: Delta = 46'sb1011111111110000000000000000000000000000000000;
		11618: Delta = 46'sb0000000001100000000000000000000000000000000000;
		6995: Delta = 46'sb1111111110100000000000000000000000000000000000;
		13159: Delta = 46'sb0000000010100000000000000000000000000000000000;
		5454: Delta = 46'sb1111111101100000000000000000000000000000000000;
		16241: Delta = 46'sb0000000100100000000000000000000000000000000000;
		3913: Delta = 46'sb1111111100100000000000000000000000000000000000;
		14700: Delta = 46'sb0000000011100000000000000000000000000000000000;
		2372: Delta = 46'sb1111111011100000000000000000000000000000000000;
		3792: Delta = 46'sb0000001000100000000000000000000000000000000000;
		16362: Delta = 46'sb1111111000100000000000000000000000000000000000;
		2251: Delta = 46'sb0000000111100000000000000000000000000000000000;
		14821: Delta = 46'sb1111110111100000000000000000000000000000000000;
		16120: Delta = 46'sb0000010000100000000000000000000000000000000000;
		4034: Delta = 46'sb1111110000100000000000000000000000000000000000;
		14579: Delta = 46'sb0000001111100000000000000000000000000000000000;
		2493: Delta = 46'sb1111101111100000000000000000000000000000000000;
		3550: Delta = 46'sb0000100000100000000000000000000000000000000000;
		16604: Delta = 46'sb1111100000100000000000000000000000000000000000;
		2009: Delta = 46'sb0000011111100000000000000000000000000000000000;
		15063: Delta = 46'sb1111011111100000000000000000000000000000000000;
		15636: Delta = 46'sb0001000000100000000000000000000000000000000000;
		4518: Delta = 46'sb1111000000100000000000000000000000000000000000;
		14095: Delta = 46'sb0000111111100000000000000000000000000000000000;
		2977: Delta = 46'sb1110111111100000000000000000000000000000000000;
		2582: Delta = 46'sb0010000000100000000000000000000000000000000000;
		17572: Delta = 46'sb1110000000100000000000000000000000000000000000;
		1041: Delta = 46'sb0001111111100000000000000000000000000000000000;
		16031: Delta = 46'sb1101111111100000000000000000000000000000000000;
		13700: Delta = 46'sb0100000000100000000000000000000000000000000000;
		6454: Delta = 46'sb1100000000100000000000000000000000000000000000;
		12159: Delta = 46'sb0011111111100000000000000000000000000000000000;
		4913: Delta = 46'sb1011111111100000000000000000000000000000000000;
		4623: Delta = 46'sb0000000011000000000000000000000000000000000000;
		13990: Delta = 46'sb1111111101000000000000000000000000000000000000;
		7705: Delta = 46'sb0000000101000000000000000000000000000000000000;
		10908: Delta = 46'sb1111111011000000000000000000000000000000000000;
		13869: Delta = 46'sb0000001001000000000000000000000000000000000000;
		7826: Delta = 46'sb1111111001000000000000000000000000000000000000;
		10787: Delta = 46'sb0000000111000000000000000000000000000000000000;
		4744: Delta = 46'sb1111110111000000000000000000000000000000000000;
		7584: Delta = 46'sb0000010001000000000000000000000000000000000000;
		14111: Delta = 46'sb1111110001000000000000000000000000000000000000;
		4502: Delta = 46'sb0000001111000000000000000000000000000000000000;
		11029: Delta = 46'sb1111101111000000000000000000000000000000000000;
		13627: Delta = 46'sb0000100001000000000000000000000000000000000000;
		8068: Delta = 46'sb1111100001000000000000000000000000000000000000;
		10545: Delta = 46'sb0000011111000000000000000000000000000000000000;
		4986: Delta = 46'sb1111011111000000000000000000000000000000000000;
		7100: Delta = 46'sb0001000001000000000000000000000000000000000000;
		14595: Delta = 46'sb1111000001000000000000000000000000000000000000;
		4018: Delta = 46'sb0000111111000000000000000000000000000000000000;
		11513: Delta = 46'sb1110111111000000000000000000000000000000000000;
		12659: Delta = 46'sb0010000001000000000000000000000000000000000000;
		9036: Delta = 46'sb1110000001000000000000000000000000000000000000;
		9577: Delta = 46'sb0001111111000000000000000000000000000000000000;
		5954: Delta = 46'sb1101111111000000000000000000000000000000000000;
		5164: Delta = 46'sb0100000001000000000000000000000000000000000000;
		16531: Delta = 46'sb1100000001000000000000000000000000000000000000;
		2082: Delta = 46'sb0011111111000000000000000000000000000000000000;
		13449: Delta = 46'sb1011111111000000000000000000000000000000000000;
		9246: Delta = 46'sb0000000110000000000000000000000000000000000000;
		9367: Delta = 46'sb1111111010000000000000000000000000000000000000;
		15410: Delta = 46'sb0000001010000000000000000000000000000000000000;
		3203: Delta = 46'sb1111110110000000000000000000000000000000000000;
		9125: Delta = 46'sb0000010010000000000000000000000000000000000000;
		15652: Delta = 46'sb1111110010000000000000000000000000000000000000;
		2961: Delta = 46'sb0000001110000000000000000000000000000000000000;
		9488: Delta = 46'sb1111101110000000000000000000000000000000000000;
		15168: Delta = 46'sb0000100010000000000000000000000000000000000000;
		9609: Delta = 46'sb1111100010000000000000000000000000000000000000;
		9004: Delta = 46'sb0000011110000000000000000000000000000000000000;
		3445: Delta = 46'sb1111011110000000000000000000000000000000000000;
		8641: Delta = 46'sb0001000010000000000000000000000000000000000000;
		16136: Delta = 46'sb1111000010000000000000000000000000000000000000;
		2477: Delta = 46'sb0000111110000000000000000000000000000000000000;
		9972: Delta = 46'sb1110111110000000000000000000000000000000000000;
		14200: Delta = 46'sb0010000010000000000000000000000000000000000000;
		10577: Delta = 46'sb1110000010000000000000000000000000000000000000;
		8036: Delta = 46'sb0001111110000000000000000000000000000000000000;
		4413: Delta = 46'sb1101111110000000000000000000000000000000000000;
		6705: Delta = 46'sb0100000010000000000000000000000000000000000000;
		18072: Delta = 46'sb1100000010000000000000000000000000000000000000;
		541: Delta = 46'sb0011111110000000000000000000000000000000000000;
		11908: Delta = 46'sb1011111110000000000000000000000000000000000000;
		18492: Delta = 46'sb0000001100000000000000000000000000000000000000;
		121: Delta = 46'sb1111110100000000000000000000000000000000000000;
		12207: Delta = 46'sb0000010100000000000000000000000000000000000000;
		6406: Delta = 46'sb1111101100000000000000000000000000000000000000;
		18250: Delta = 46'sb0000100100000000000000000000000000000000000000;
		12691: Delta = 46'sb1111100100000000000000000000000000000000000000;
		5922: Delta = 46'sb0000011100000000000000000000000000000000000000;
		363: Delta = 46'sb1111011100000000000000000000000000000000000000;
		11723: Delta = 46'sb0001000100000000000000000000000000000000000000;
		605: Delta = 46'sb1111000100000000000000000000000000000000000000;
		18008: Delta = 46'sb0000111100000000000000000000000000000000000000;
		6890: Delta = 46'sb1110111100000000000000000000000000000000000000;
		17282: Delta = 46'sb0010000100000000000000000000000000000000000000;
		13659: Delta = 46'sb1110000100000000000000000000000000000000000000;
		4954: Delta = 46'sb0001111100000000000000000000000000000000000000;
		1331: Delta = 46'sb1101111100000000000000000000000000000000000000;
		9787: Delta = 46'sb0100000100000000000000000000000000000000000000;
		2541: Delta = 46'sb1100000100000000000000000000000000000000000000;
		16072: Delta = 46'sb0011111100000000000000000000000000000000000000;
		8826: Delta = 46'sb1011111100000000000000000000000000000000000000;
		18371: Delta = 46'sb0000011000000000000000000000000000000000000000;
		242: Delta = 46'sb1111101000000000000000000000000000000000000000;
		5801: Delta = 46'sb0000101000000000000000000000000000000000000000;
		12812: Delta = 46'sb1111011000000000000000000000000000000000000000;
		17887: Delta = 46'sb0001001000000000000000000000000000000000000000;
		6769: Delta = 46'sb1111001000000000000000000000000000000000000000;
		11844: Delta = 46'sb0000111000000000000000000000000000000000000000;
		726: Delta = 46'sb1110111000000000000000000000000000000000000000;
		4833: Delta = 46'sb0010001000000000000000000000000000000000000000;
		1210: Delta = 46'sb1110001000000000000000000000000000000000000000;
		17403: Delta = 46'sb0001111000000000000000000000000000000000000000;
		13780: Delta = 46'sb1101111000000000000000000000000000000000000000;
		15951: Delta = 46'sb0100001000000000000000000000000000000000000000;
		8705: Delta = 46'sb1100001000000000000000000000000000000000000000;
		9908: Delta = 46'sb0011111000000000000000000000000000000000000000;
		2662: Delta = 46'sb1011111000000000000000000000000000000000000000;
		18129: Delta = 46'sb0000110000000000000000000000000000000000000000;
		484: Delta = 46'sb1111010000000000000000000000000000000000000000;
		11602: Delta = 46'sb0001010000000000000000000000000000000000000000;
		7011: Delta = 46'sb1110110000000000000000000000000000000000000000;
		17161: Delta = 46'sb0010010000000000000000000000000000000000000000;
		13538: Delta = 46'sb1110010000000000000000000000000000000000000000;
		5075: Delta = 46'sb0001110000000000000000000000000000000000000000;
		1452: Delta = 46'sb1101110000000000000000000000000000000000000000;
		9666: Delta = 46'sb0100010000000000000000000000000000000000000000;
		2420: Delta = 46'sb1100010000000000000000000000000000000000000000;
		16193: Delta = 46'sb0011110000000000000000000000000000000000000000;
		8947: Delta = 46'sb1011110000000000000000000000000000000000000000;
		17645: Delta = 46'sb0001100000000000000000000000000000000000000000;
		968: Delta = 46'sb1110100000000000000000000000000000000000000000;
		4591: Delta = 46'sb0010100000000000000000000000000000000000000000;
		14022: Delta = 46'sb1101100000000000000000000000000000000000000000;
		15709: Delta = 46'sb0100100000000000000000000000000000000000000000;
		8463: Delta = 46'sb1100100000000000000000000000000000000000000000;
		10150: Delta = 46'sb0011100000000000000000000000000000000000000000;
		2904: Delta = 46'sb1011100000000000000000000000000000000000000000;
		16677: Delta = 46'sb0011000000000000000000000000000000000000000000;
		1936: Delta = 46'sb1101000000000000000000000000000000000000000000;
		9182: Delta = 46'sb0101000000000000000000000000000000000000000000;
		9431: Delta = 46'sb1011000000000000000000000000000000000000000000;
		14741: Delta = 46'sb0110000000000000000000000000000000000000000000;
		3872: Delta = 46'sb1010000000000000000000000000000000000000000000;
		default: Delta =46'sb0;
	endcase
end

wire signed [W_BITS-1:0] W_signed;
assign W_signed = (W - Delta);

always@(posedge clk or negedge rst_n) begin
   if(!rst_n) begin
     	ps <= idle;
    end
   else begin
        case(ps)
            idle: begin
                found <= 0;
                R <= 0;
        	Q <= 0;
                ps <= pre;
                end
	    pre: begin
		 Q <= W / A;
		 ps <= load;
		end
            load: begin
                 R <= W - (A * Q);
		 ps <= LUT;
		end
	    LUT: begin
		  if(Delta != 0)begin
		      N <= W_signed / A ;	
		      found <= 1;
                      ps <= idle;
		  end
		  else begin
		      N <= Q;
		      found <= 1;
                      ps <= idle;
		  end
		end
	endcase
    end
end

endmodule

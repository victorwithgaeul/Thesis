// Product (AN) Code DEC r-LUT
// DEC_rLUT30bits.v
// Used to do DEC, but corrected errors by locations, not AWE
// Received remainder r, output two error locations.
module DEC_rLUT30bits(r, l_1, l_2);
input 	[14:0]	r;
output	reg	signed	[6:0]	l_1;
output	reg	signed	[6:0]	l_2;
always@(*) begin
	case(r)
		1: begin l_1 = -1;
				 l_2 = +2; end
		18612: begin l_1 = +1;
				 l_2 = -2; end
		2: begin l_1 = +1;
				 l_2 = +1; end
		18611: begin l_1 = -1;
				 l_2 = -1; end
		4: begin l_1 = +2;
				 l_2 = +2; end
		18609: begin l_1 = -2;
				 l_2 = -2; end
		8: begin l_1 = +3;
				 l_2 = +3; end
		18605: begin l_1 = -3;
				 l_2 = -3; end
		16: begin l_1 = +4;
				 l_2 = +4; end
		18597: begin l_1 = -4;
				 l_2 = -4; end
		32: begin l_1 = +5;
				 l_2 = +5; end
		18581: begin l_1 = -5;
				 l_2 = -5; end
		64: begin l_1 = +6;
				 l_2 = +6; end
		18549: begin l_1 = -6;
				 l_2 = -6; end
		128: begin l_1 = +7;
				 l_2 = +7; end
		18485: begin l_1 = -7;
				 l_2 = -7; end
		256: begin l_1 = +8;
				 l_2 = +8; end
		18357: begin l_1 = -8;
				 l_2 = -8; end
		512: begin l_1 = +9;
				 l_2 = +9; end
		18101: begin l_1 = -9;
				 l_2 = -9; end
		1024: begin l_1 = +10;
				 l_2 = +10; end
		17589: begin l_1 = -10;
				 l_2 = -10; end
		2048: begin l_1 = +11;
				 l_2 = +11; end
		16565: begin l_1 = -11;
				 l_2 = -11; end
		4096: begin l_1 = +12;
				 l_2 = +12; end
		14517: begin l_1 = -12;
				 l_2 = -12; end
		8192: begin l_1 = +13;
				 l_2 = +13; end
		10421: begin l_1 = -13;
				 l_2 = -13; end
		16384: begin l_1 = +14;
				 l_2 = +14; end
		2229: begin l_1 = -14;
				 l_2 = -14; end
		14155: begin l_1 = +15;
				 l_2 = +15; end
		4458: begin l_1 = -15;
				 l_2 = -15; end
		9697: begin l_1 = +16;
				 l_2 = +16; end
		8916: begin l_1 = -16;
				 l_2 = -16; end
		781: begin l_1 = +17;
				 l_2 = +17; end
		17832: begin l_1 = -17;
				 l_2 = -17; end
		1562: begin l_1 = +18;
				 l_2 = +18; end
		17051: begin l_1 = -18;
				 l_2 = -18; end
		3124: begin l_1 = +19;
				 l_2 = +19; end
		15489: begin l_1 = -19;
				 l_2 = -19; end
		6248: begin l_1 = +20;
				 l_2 = +20; end
		12365: begin l_1 = -20;
				 l_2 = -20; end
		12496: begin l_1 = +21;
				 l_2 = +21; end
		6117: begin l_1 = -21;
				 l_2 = -21; end
		6379: begin l_1 = +22;
				 l_2 = +22; end
		12234: begin l_1 = -22;
				 l_2 = -22; end
		12758: begin l_1 = +23;
				 l_2 = +23; end
		5855: begin l_1 = -23;
				 l_2 = -23; end
		6903: begin l_1 = +24;
				 l_2 = +24; end
		11710: begin l_1 = -24;
				 l_2 = -24; end
		13806: begin l_1 = +25;
				 l_2 = +25; end
		4807: begin l_1 = -25;
				 l_2 = -25; end
		8999: begin l_1 = +26;
				 l_2 = +26; end
		9614: begin l_1 = -26;
				 l_2 = -26; end
		17998: begin l_1 = +27;
				 l_2 = +27; end
		615: begin l_1 = -27;
				 l_2 = -27; end
		17383: begin l_1 = +28;
				 l_2 = +28; end
		1230: begin l_1 = -28;
				 l_2 = -28; end
		16153: begin l_1 = +29;
				 l_2 = +29; end
		2460: begin l_1 = -29;
				 l_2 = -29; end
		13693: begin l_1 = +30;
				 l_2 = +30; end
		4920: begin l_1 = -30;
				 l_2 = -30; end
		8773: begin l_1 = +31;
				 l_2 = +31; end
		9840: begin l_1 = -31;
				 l_2 = -31; end
		17546: begin l_1 = +32;
				 l_2 = +32; end
		1067: begin l_1 = -32;
				 l_2 = -32; end
		16479: begin l_1 = +33;
				 l_2 = +33; end
		2134: begin l_1 = -33;
				 l_2 = -33; end
		14345: begin l_1 = +34;
				 l_2 = +34; end
		4268: begin l_1 = -34;
				 l_2 = -34; end
		10077: begin l_1 = +35;
				 l_2 = +35; end
		8536: begin l_1 = -35;
				 l_2 = -35; end
		1541: begin l_1 = +36;
				 l_2 = +36; end
		17072: begin l_1 = -36;
				 l_2 = -36; end
		3082: begin l_1 = +37;
				 l_2 = +37; end
		15531: begin l_1 = -37;
				 l_2 = -37; end
		6164: begin l_1 = +38;
				 l_2 = +38; end
		12449: begin l_1 = -38;
				 l_2 = -38; end
		12328: begin l_1 = +39;
				 l_2 = +39; end
		6285: begin l_1 = -39;
				 l_2 = -39; end
		6043: begin l_1 = +40;
				 l_2 = +40; end
		12570: begin l_1 = -40;
				 l_2 = -40; end
		12086: begin l_1 = +41;
				 l_2 = +41; end
		6527: begin l_1 = -41;
				 l_2 = -41; end
		5559: begin l_1 = +42;
				 l_2 = +42; end
		13054: begin l_1 = -42;
				 l_2 = -42; end
		11118: begin l_1 = +43;
				 l_2 = +43; end
		7495: begin l_1 = -43;
				 l_2 = -43; end
		3623: begin l_1 = +44;
				 l_2 = +44; end
		14990: begin l_1 = -44;
				 l_2 = -44; end
		3: begin l_1 = -1;
				 l_2 = +3; end
		18610: begin l_1 = -1;
				 l_2 = -2; end
		5: begin l_1 = +1;
				 l_2 = +3; end
		18608: begin l_1 = -1;
				 l_2 = -3; end
		9: begin l_1 = +1;
				 l_2 = +4; end
		18606: begin l_1 = +1;
				 l_2 = -4; end
		7: begin l_1 = -1;
				 l_2 = +4; end
		18604: begin l_1 = -1;
				 l_2 = -4; end
		17: begin l_1 = +1;
				 l_2 = +5; end
		18598: begin l_1 = +1;
				 l_2 = -5; end
		15: begin l_1 = -1;
				 l_2 = +5; end
		18596: begin l_1 = -1;
				 l_2 = -5; end
		33: begin l_1 = +1;
				 l_2 = +6; end
		18582: begin l_1 = +1;
				 l_2 = -6; end
		31: begin l_1 = -1;
				 l_2 = +6; end
		18580: begin l_1 = -1;
				 l_2 = -6; end
		65: begin l_1 = +1;
				 l_2 = +7; end
		18550: begin l_1 = +1;
				 l_2 = -7; end
		63: begin l_1 = -1;
				 l_2 = +7; end
		18548: begin l_1 = -1;
				 l_2 = -7; end
		129: begin l_1 = +1;
				 l_2 = +8; end
		18486: begin l_1 = +1;
				 l_2 = -8; end
		127: begin l_1 = -1;
				 l_2 = +8; end
		18484: begin l_1 = -1;
				 l_2 = -8; end
		257: begin l_1 = +1;
				 l_2 = +9; end
		18358: begin l_1 = +1;
				 l_2 = -9; end
		255: begin l_1 = -1;
				 l_2 = +9; end
		18356: begin l_1 = -1;
				 l_2 = -9; end
		513: begin l_1 = +1;
				 l_2 = +10; end
		18102: begin l_1 = +1;
				 l_2 = -10; end
		511: begin l_1 = -1;
				 l_2 = +10; end
		18100: begin l_1 = -1;
				 l_2 = -10; end
		1025: begin l_1 = +1;
				 l_2 = +11; end
		17590: begin l_1 = +1;
				 l_2 = -11; end
		1023: begin l_1 = -1;
				 l_2 = +11; end
		17588: begin l_1 = -1;
				 l_2 = -11; end
		2049: begin l_1 = +1;
				 l_2 = +12; end
		16566: begin l_1 = +1;
				 l_2 = -12; end
		2047: begin l_1 = -1;
				 l_2 = +12; end
		16564: begin l_1 = -1;
				 l_2 = -12; end
		4097: begin l_1 = +1;
				 l_2 = +13; end
		14518: begin l_1 = +1;
				 l_2 = -13; end
		4095: begin l_1 = -1;
				 l_2 = +13; end
		14516: begin l_1 = -1;
				 l_2 = -13; end
		8193: begin l_1 = +1;
				 l_2 = +14; end
		10422: begin l_1 = +1;
				 l_2 = -14; end
		8191: begin l_1 = -1;
				 l_2 = +14; end
		10420: begin l_1 = -1;
				 l_2 = -14; end
		16385: begin l_1 = +1;
				 l_2 = +15; end
		2230: begin l_1 = +1;
				 l_2 = -15; end
		16383: begin l_1 = -1;
				 l_2 = +15; end
		2228: begin l_1 = -1;
				 l_2 = -15; end
		14156: begin l_1 = +1;
				 l_2 = +16; end
		4459: begin l_1 = +1;
				 l_2 = -16; end
		14154: begin l_1 = -1;
				 l_2 = +16; end
		4457: begin l_1 = -1;
				 l_2 = -16; end
		9698: begin l_1 = +1;
				 l_2 = +17; end
		8917: begin l_1 = +1;
				 l_2 = -17; end
		9696: begin l_1 = -1;
				 l_2 = +17; end
		8915: begin l_1 = -1;
				 l_2 = -17; end
		782: begin l_1 = +1;
				 l_2 = +18; end
		17833: begin l_1 = +1;
				 l_2 = -18; end
		780: begin l_1 = -1;
				 l_2 = +18; end
		17831: begin l_1 = -1;
				 l_2 = -18; end
		1563: begin l_1 = +1;
				 l_2 = +19; end
		17052: begin l_1 = +1;
				 l_2 = -19; end
		1561: begin l_1 = -1;
				 l_2 = +19; end
		17050: begin l_1 = -1;
				 l_2 = -19; end
		3125: begin l_1 = +1;
				 l_2 = +20; end
		15490: begin l_1 = +1;
				 l_2 = -20; end
		3123: begin l_1 = -1;
				 l_2 = +20; end
		15488: begin l_1 = -1;
				 l_2 = -20; end
		6249: begin l_1 = +1;
				 l_2 = +21; end
		12366: begin l_1 = +1;
				 l_2 = -21; end
		6247: begin l_1 = -1;
				 l_2 = +21; end
		12364: begin l_1 = -1;
				 l_2 = -21; end
		12497: begin l_1 = +1;
				 l_2 = +22; end
		6118: begin l_1 = +1;
				 l_2 = -22; end
		12495: begin l_1 = -1;
				 l_2 = +22; end
		6116: begin l_1 = -1;
				 l_2 = -22; end
		6380: begin l_1 = +1;
				 l_2 = +23; end
		12235: begin l_1 = +1;
				 l_2 = -23; end
		6378: begin l_1 = -1;
				 l_2 = +23; end
		12233: begin l_1 = -1;
				 l_2 = -23; end
		12759: begin l_1 = +1;
				 l_2 = +24; end
		5856: begin l_1 = +1;
				 l_2 = -24; end
		12757: begin l_1 = -1;
				 l_2 = +24; end
		5854: begin l_1 = -1;
				 l_2 = -24; end
		6904: begin l_1 = +1;
				 l_2 = +25; end
		11711: begin l_1 = +1;
				 l_2 = -25; end
		6902: begin l_1 = -1;
				 l_2 = +25; end
		11709: begin l_1 = -1;
				 l_2 = -25; end
		13807: begin l_1 = +1;
				 l_2 = +26; end
		4808: begin l_1 = +1;
				 l_2 = -26; end
		13805: begin l_1 = -1;
				 l_2 = +26; end
		4806: begin l_1 = -1;
				 l_2 = -26; end
		9000: begin l_1 = +1;
				 l_2 = +27; end
		9615: begin l_1 = +1;
				 l_2 = -27; end
		8998: begin l_1 = -1;
				 l_2 = +27; end
		9613: begin l_1 = -1;
				 l_2 = -27; end
		17999: begin l_1 = +1;
				 l_2 = +28; end
		616: begin l_1 = +1;
				 l_2 = -28; end
		17997: begin l_1 = -1;
				 l_2 = +28; end
		614: begin l_1 = -1;
				 l_2 = -28; end
		17384: begin l_1 = +1;
				 l_2 = +29; end
		1231: begin l_1 = +1;
				 l_2 = -29; end
		17382: begin l_1 = -1;
				 l_2 = +29; end
		1229: begin l_1 = -1;
				 l_2 = -29; end
		16154: begin l_1 = +1;
				 l_2 = +30; end
		2461: begin l_1 = +1;
				 l_2 = -30; end
		16152: begin l_1 = -1;
				 l_2 = +30; end
		2459: begin l_1 = -1;
				 l_2 = -30; end
		13694: begin l_1 = +1;
				 l_2 = +31; end
		4921: begin l_1 = +1;
				 l_2 = -31; end
		13692: begin l_1 = -1;
				 l_2 = +31; end
		4919: begin l_1 = -1;
				 l_2 = -31; end
		8774: begin l_1 = +1;
				 l_2 = +32; end
		9841: begin l_1 = +1;
				 l_2 = -32; end
		8772: begin l_1 = -1;
				 l_2 = +32; end
		9839: begin l_1 = -1;
				 l_2 = -32; end
		17547: begin l_1 = +1;
				 l_2 = +33; end
		1068: begin l_1 = +1;
				 l_2 = -33; end
		17545: begin l_1 = -1;
				 l_2 = +33; end
		1066: begin l_1 = -1;
				 l_2 = -33; end
		16480: begin l_1 = +1;
				 l_2 = +34; end
		2135: begin l_1 = +1;
				 l_2 = -34; end
		16478: begin l_1 = -1;
				 l_2 = +34; end
		2133: begin l_1 = -1;
				 l_2 = -34; end
		14346: begin l_1 = +1;
				 l_2 = +35; end
		4269: begin l_1 = +1;
				 l_2 = -35; end
		14344: begin l_1 = -1;
				 l_2 = +35; end
		4267: begin l_1 = -1;
				 l_2 = -35; end
		10078: begin l_1 = +1;
				 l_2 = +36; end
		8537: begin l_1 = +1;
				 l_2 = -36; end
		10076: begin l_1 = -1;
				 l_2 = +36; end
		8535: begin l_1 = -1;
				 l_2 = -36; end
		1542: begin l_1 = +1;
				 l_2 = +37; end
		17073: begin l_1 = +1;
				 l_2 = -37; end
		1540: begin l_1 = -1;
				 l_2 = +37; end
		17071: begin l_1 = -1;
				 l_2 = -37; end
		3083: begin l_1 = +1;
				 l_2 = +38; end
		15532: begin l_1 = +1;
				 l_2 = -38; end
		3081: begin l_1 = -1;
				 l_2 = +38; end
		15530: begin l_1 = -1;
				 l_2 = -38; end
		6165: begin l_1 = +1;
				 l_2 = +39; end
		12450: begin l_1 = +1;
				 l_2 = -39; end
		6163: begin l_1 = -1;
				 l_2 = +39; end
		12448: begin l_1 = -1;
				 l_2 = -39; end
		12329: begin l_1 = +1;
				 l_2 = +40; end
		6286: begin l_1 = +1;
				 l_2 = -40; end
		12327: begin l_1 = -1;
				 l_2 = +40; end
		6284: begin l_1 = -1;
				 l_2 = -40; end
		6044: begin l_1 = +1;
				 l_2 = +41; end
		12571: begin l_1 = +1;
				 l_2 = -41; end
		6042: begin l_1 = -1;
				 l_2 = +41; end
		12569: begin l_1 = -1;
				 l_2 = -41; end
		12087: begin l_1 = +1;
				 l_2 = +42; end
		6528: begin l_1 = +1;
				 l_2 = -42; end
		12085: begin l_1 = -1;
				 l_2 = +42; end
		6526: begin l_1 = -1;
				 l_2 = -42; end
		5560: begin l_1 = +1;
				 l_2 = +43; end
		13055: begin l_1 = +1;
				 l_2 = -43; end
		5558: begin l_1 = -1;
				 l_2 = +43; end
		13053: begin l_1 = -1;
				 l_2 = -43; end
		11119: begin l_1 = +1;
				 l_2 = +44; end
		7496: begin l_1 = +1;
				 l_2 = -44; end
		11117: begin l_1 = -1;
				 l_2 = +44; end
		7494: begin l_1 = -1;
				 l_2 = -44; end
		3624: begin l_1 = +1;
				 l_2 = +45; end
		14991: begin l_1 = +1;
				 l_2 = -45; end
		3622: begin l_1 = -1;
				 l_2 = +45; end
		14989: begin l_1 = -1;
				 l_2 = -45; end
		6: begin l_1 = -2;
				 l_2 = +4; end
		18607: begin l_1 = -2;
				 l_2 = -3; end
		10: begin l_1 = +2;
				 l_2 = +4; end
		18603: begin l_1 = -2;
				 l_2 = -4; end
		18: begin l_1 = +2;
				 l_2 = +5; end
		18599: begin l_1 = +2;
				 l_2 = -5; end
		14: begin l_1 = -2;
				 l_2 = +5; end
		18595: begin l_1 = -2;
				 l_2 = -5; end
		34: begin l_1 = +2;
				 l_2 = +6; end
		18583: begin l_1 = +2;
				 l_2 = -6; end
		30: begin l_1 = -2;
				 l_2 = +6; end
		18579: begin l_1 = -2;
				 l_2 = -6; end
		66: begin l_1 = +2;
				 l_2 = +7; end
		18551: begin l_1 = +2;
				 l_2 = -7; end
		62: begin l_1 = -2;
				 l_2 = +7; end
		18547: begin l_1 = -2;
				 l_2 = -7; end
		130: begin l_1 = +2;
				 l_2 = +8; end
		18487: begin l_1 = +2;
				 l_2 = -8; end
		126: begin l_1 = -2;
				 l_2 = +8; end
		18483: begin l_1 = -2;
				 l_2 = -8; end
		258: begin l_1 = +2;
				 l_2 = +9; end
		18359: begin l_1 = +2;
				 l_2 = -9; end
		254: begin l_1 = -2;
				 l_2 = +9; end
		18355: begin l_1 = -2;
				 l_2 = -9; end
		514: begin l_1 = +2;
				 l_2 = +10; end
		18103: begin l_1 = +2;
				 l_2 = -10; end
		510: begin l_1 = -2;
				 l_2 = +10; end
		18099: begin l_1 = -2;
				 l_2 = -10; end
		1026: begin l_1 = +2;
				 l_2 = +11; end
		17591: begin l_1 = +2;
				 l_2 = -11; end
		1022: begin l_1 = -2;
				 l_2 = +11; end
		17587: begin l_1 = -2;
				 l_2 = -11; end
		2050: begin l_1 = +2;
				 l_2 = +12; end
		16567: begin l_1 = +2;
				 l_2 = -12; end
		2046: begin l_1 = -2;
				 l_2 = +12; end
		16563: begin l_1 = -2;
				 l_2 = -12; end
		4098: begin l_1 = +2;
				 l_2 = +13; end
		14519: begin l_1 = +2;
				 l_2 = -13; end
		4094: begin l_1 = -2;
				 l_2 = +13; end
		14515: begin l_1 = -2;
				 l_2 = -13; end
		8194: begin l_1 = +2;
				 l_2 = +14; end
		10423: begin l_1 = +2;
				 l_2 = -14; end
		8190: begin l_1 = -2;
				 l_2 = +14; end
		10419: begin l_1 = -2;
				 l_2 = -14; end
		16386: begin l_1 = +2;
				 l_2 = +15; end
		2231: begin l_1 = +2;
				 l_2 = -15; end
		16382: begin l_1 = -2;
				 l_2 = +15; end
		2227: begin l_1 = -2;
				 l_2 = -15; end
		14157: begin l_1 = +2;
				 l_2 = +16; end
		4460: begin l_1 = +2;
				 l_2 = -16; end
		14153: begin l_1 = -2;
				 l_2 = +16; end
		4456: begin l_1 = -2;
				 l_2 = -16; end
		9699: begin l_1 = +2;
				 l_2 = +17; end
		8918: begin l_1 = +2;
				 l_2 = -17; end
		9695: begin l_1 = -2;
				 l_2 = +17; end
		8914: begin l_1 = -2;
				 l_2 = -17; end
		783: begin l_1 = +2;
				 l_2 = +18; end
		17834: begin l_1 = +2;
				 l_2 = -18; end
		779: begin l_1 = -2;
				 l_2 = +18; end
		17830: begin l_1 = -2;
				 l_2 = -18; end
		1564: begin l_1 = +2;
				 l_2 = +19; end
		17053: begin l_1 = +2;
				 l_2 = -19; end
		1560: begin l_1 = -2;
				 l_2 = +19; end
		17049: begin l_1 = -2;
				 l_2 = -19; end
		3126: begin l_1 = +2;
				 l_2 = +20; end
		15491: begin l_1 = +2;
				 l_2 = -20; end
		3122: begin l_1 = -2;
				 l_2 = +20; end
		15487: begin l_1 = -2;
				 l_2 = -20; end
		6250: begin l_1 = +2;
				 l_2 = +21; end
		12367: begin l_1 = +2;
				 l_2 = -21; end
		6246: begin l_1 = -2;
				 l_2 = +21; end
		12363: begin l_1 = -2;
				 l_2 = -21; end
		12498: begin l_1 = +2;
				 l_2 = +22; end
		6119: begin l_1 = +2;
				 l_2 = -22; end
		12494: begin l_1 = -2;
				 l_2 = +22; end
		6115: begin l_1 = -2;
				 l_2 = -22; end
		6381: begin l_1 = +2;
				 l_2 = +23; end
		12236: begin l_1 = +2;
				 l_2 = -23; end
		6377: begin l_1 = -2;
				 l_2 = +23; end
		12232: begin l_1 = -2;
				 l_2 = -23; end
		12760: begin l_1 = +2;
				 l_2 = +24; end
		5857: begin l_1 = +2;
				 l_2 = -24; end
		12756: begin l_1 = -2;
				 l_2 = +24; end
		5853: begin l_1 = -2;
				 l_2 = -24; end
		6905: begin l_1 = +2;
				 l_2 = +25; end
		11712: begin l_1 = +2;
				 l_2 = -25; end
		6901: begin l_1 = -2;
				 l_2 = +25; end
		11708: begin l_1 = -2;
				 l_2 = -25; end
		13808: begin l_1 = +2;
				 l_2 = +26; end
		4809: begin l_1 = +2;
				 l_2 = -26; end
		13804: begin l_1 = -2;
				 l_2 = +26; end
		4805: begin l_1 = -2;
				 l_2 = -26; end
		9001: begin l_1 = +2;
				 l_2 = +27; end
		9616: begin l_1 = +2;
				 l_2 = -27; end
		8997: begin l_1 = -2;
				 l_2 = +27; end
		9612: begin l_1 = -2;
				 l_2 = -27; end
		18000: begin l_1 = +2;
				 l_2 = +28; end
		617: begin l_1 = +2;
				 l_2 = -28; end
		17996: begin l_1 = -2;
				 l_2 = +28; end
		613: begin l_1 = -2;
				 l_2 = -28; end
		17385: begin l_1 = +2;
				 l_2 = +29; end
		1232: begin l_1 = +2;
				 l_2 = -29; end
		17381: begin l_1 = -2;
				 l_2 = +29; end
		1228: begin l_1 = -2;
				 l_2 = -29; end
		16155: begin l_1 = +2;
				 l_2 = +30; end
		2462: begin l_1 = +2;
				 l_2 = -30; end
		16151: begin l_1 = -2;
				 l_2 = +30; end
		2458: begin l_1 = -2;
				 l_2 = -30; end
		13695: begin l_1 = +2;
				 l_2 = +31; end
		4922: begin l_1 = +2;
				 l_2 = -31; end
		13691: begin l_1 = -2;
				 l_2 = +31; end
		4918: begin l_1 = -2;
				 l_2 = -31; end
		8775: begin l_1 = +2;
				 l_2 = +32; end
		9842: begin l_1 = +2;
				 l_2 = -32; end
		8771: begin l_1 = -2;
				 l_2 = +32; end
		9838: begin l_1 = -2;
				 l_2 = -32; end
		17548: begin l_1 = +2;
				 l_2 = +33; end
		1069: begin l_1 = +2;
				 l_2 = -33; end
		17544: begin l_1 = -2;
				 l_2 = +33; end
		1065: begin l_1 = -2;
				 l_2 = -33; end
		16481: begin l_1 = +2;
				 l_2 = +34; end
		2136: begin l_1 = +2;
				 l_2 = -34; end
		16477: begin l_1 = -2;
				 l_2 = +34; end
		2132: begin l_1 = -2;
				 l_2 = -34; end
		14347: begin l_1 = +2;
				 l_2 = +35; end
		4270: begin l_1 = +2;
				 l_2 = -35; end
		14343: begin l_1 = -2;
				 l_2 = +35; end
		4266: begin l_1 = -2;
				 l_2 = -35; end
		10079: begin l_1 = +2;
				 l_2 = +36; end
		8538: begin l_1 = +2;
				 l_2 = -36; end
		10075: begin l_1 = -2;
				 l_2 = +36; end
		8534: begin l_1 = -2;
				 l_2 = -36; end
		1543: begin l_1 = +2;
				 l_2 = +37; end
		17074: begin l_1 = +2;
				 l_2 = -37; end
		1539: begin l_1 = -2;
				 l_2 = +37; end
		17070: begin l_1 = -2;
				 l_2 = -37; end
		3084: begin l_1 = +2;
				 l_2 = +38; end
		15533: begin l_1 = +2;
				 l_2 = -38; end
		3080: begin l_1 = -2;
				 l_2 = +38; end
		15529: begin l_1 = -2;
				 l_2 = -38; end
		6166: begin l_1 = +2;
				 l_2 = +39; end
		12451: begin l_1 = +2;
				 l_2 = -39; end
		6162: begin l_1 = -2;
				 l_2 = +39; end
		12447: begin l_1 = -2;
				 l_2 = -39; end
		12330: begin l_1 = +2;
				 l_2 = +40; end
		6287: begin l_1 = +2;
				 l_2 = -40; end
		12326: begin l_1 = -2;
				 l_2 = +40; end
		6283: begin l_1 = -2;
				 l_2 = -40; end
		6045: begin l_1 = +2;
				 l_2 = +41; end
		12572: begin l_1 = +2;
				 l_2 = -41; end
		6041: begin l_1 = -2;
				 l_2 = +41; end
		12568: begin l_1 = -2;
				 l_2 = -41; end
		12088: begin l_1 = +2;
				 l_2 = +42; end
		6529: begin l_1 = +2;
				 l_2 = -42; end
		12084: begin l_1 = -2;
				 l_2 = +42; end
		6525: begin l_1 = -2;
				 l_2 = -42; end
		5561: begin l_1 = +2;
				 l_2 = +43; end
		13056: begin l_1 = +2;
				 l_2 = -43; end
		5557: begin l_1 = -2;
				 l_2 = +43; end
		13052: begin l_1 = -2;
				 l_2 = -43; end
		11120: begin l_1 = +2;
				 l_2 = +44; end
		7497: begin l_1 = +2;
				 l_2 = -44; end
		11116: begin l_1 = -2;
				 l_2 = +44; end
		7493: begin l_1 = -2;
				 l_2 = -44; end
		3625: begin l_1 = +2;
				 l_2 = +45; end
		14992: begin l_1 = +2;
				 l_2 = -45; end
		3621: begin l_1 = -2;
				 l_2 = +45; end
		14988: begin l_1 = -2;
				 l_2 = -45; end
		12: begin l_1 = -3;
				 l_2 = +5; end
		18601: begin l_1 = -3;
				 l_2 = -4; end
		20: begin l_1 = +3;
				 l_2 = +5; end
		18593: begin l_1 = -3;
				 l_2 = -5; end
		36: begin l_1 = +3;
				 l_2 = +6; end
		18585: begin l_1 = +3;
				 l_2 = -6; end
		28: begin l_1 = -3;
				 l_2 = +6; end
		18577: begin l_1 = -3;
				 l_2 = -6; end
		68: begin l_1 = +3;
				 l_2 = +7; end
		18553: begin l_1 = +3;
				 l_2 = -7; end
		60: begin l_1 = -3;
				 l_2 = +7; end
		18545: begin l_1 = -3;
				 l_2 = -7; end
		132: begin l_1 = +3;
				 l_2 = +8; end
		18489: begin l_1 = +3;
				 l_2 = -8; end
		124: begin l_1 = -3;
				 l_2 = +8; end
		18481: begin l_1 = -3;
				 l_2 = -8; end
		260: begin l_1 = +3;
				 l_2 = +9; end
		18361: begin l_1 = +3;
				 l_2 = -9; end
		252: begin l_1 = -3;
				 l_2 = +9; end
		18353: begin l_1 = -3;
				 l_2 = -9; end
		516: begin l_1 = +3;
				 l_2 = +10; end
		18105: begin l_1 = +3;
				 l_2 = -10; end
		508: begin l_1 = -3;
				 l_2 = +10; end
		18097: begin l_1 = -3;
				 l_2 = -10; end
		1028: begin l_1 = +3;
				 l_2 = +11; end
		17593: begin l_1 = +3;
				 l_2 = -11; end
		1020: begin l_1 = -3;
				 l_2 = +11; end
		17585: begin l_1 = -3;
				 l_2 = -11; end
		2052: begin l_1 = +3;
				 l_2 = +12; end
		16569: begin l_1 = +3;
				 l_2 = -12; end
		2044: begin l_1 = -3;
				 l_2 = +12; end
		16561: begin l_1 = -3;
				 l_2 = -12; end
		4100: begin l_1 = +3;
				 l_2 = +13; end
		14521: begin l_1 = +3;
				 l_2 = -13; end
		4092: begin l_1 = -3;
				 l_2 = +13; end
		14513: begin l_1 = -3;
				 l_2 = -13; end
		8196: begin l_1 = +3;
				 l_2 = +14; end
		10425: begin l_1 = +3;
				 l_2 = -14; end
		8188: begin l_1 = -3;
				 l_2 = +14; end
		10417: begin l_1 = -3;
				 l_2 = -14; end
		16388: begin l_1 = +3;
				 l_2 = +15; end
		2233: begin l_1 = +3;
				 l_2 = -15; end
		16380: begin l_1 = -3;
				 l_2 = +15; end
		2225: begin l_1 = -3;
				 l_2 = -15; end
		14159: begin l_1 = +3;
				 l_2 = +16; end
		4462: begin l_1 = +3;
				 l_2 = -16; end
		14151: begin l_1 = -3;
				 l_2 = +16; end
		4454: begin l_1 = -3;
				 l_2 = -16; end
		9701: begin l_1 = +3;
				 l_2 = +17; end
		8920: begin l_1 = +3;
				 l_2 = -17; end
		9693: begin l_1 = -3;
				 l_2 = +17; end
		8912: begin l_1 = -3;
				 l_2 = -17; end
		785: begin l_1 = +3;
				 l_2 = +18; end
		17836: begin l_1 = +3;
				 l_2 = -18; end
		777: begin l_1 = -3;
				 l_2 = +18; end
		17828: begin l_1 = -3;
				 l_2 = -18; end
		1566: begin l_1 = +3;
				 l_2 = +19; end
		17055: begin l_1 = +3;
				 l_2 = -19; end
		1558: begin l_1 = -3;
				 l_2 = +19; end
		17047: begin l_1 = -3;
				 l_2 = -19; end
		3128: begin l_1 = +3;
				 l_2 = +20; end
		15493: begin l_1 = +3;
				 l_2 = -20; end
		3120: begin l_1 = -3;
				 l_2 = +20; end
		15485: begin l_1 = -3;
				 l_2 = -20; end
		6252: begin l_1 = +3;
				 l_2 = +21; end
		12369: begin l_1 = +3;
				 l_2 = -21; end
		6244: begin l_1 = -3;
				 l_2 = +21; end
		12361: begin l_1 = -3;
				 l_2 = -21; end
		12500: begin l_1 = +3;
				 l_2 = +22; end
		6121: begin l_1 = +3;
				 l_2 = -22; end
		12492: begin l_1 = -3;
				 l_2 = +22; end
		6113: begin l_1 = -3;
				 l_2 = -22; end
		6383: begin l_1 = +3;
				 l_2 = +23; end
		12238: begin l_1 = +3;
				 l_2 = -23; end
		6375: begin l_1 = -3;
				 l_2 = +23; end
		12230: begin l_1 = -3;
				 l_2 = -23; end
		12762: begin l_1 = +3;
				 l_2 = +24; end
		5859: begin l_1 = +3;
				 l_2 = -24; end
		12754: begin l_1 = -3;
				 l_2 = +24; end
		5851: begin l_1 = -3;
				 l_2 = -24; end
		6907: begin l_1 = +3;
				 l_2 = +25; end
		11714: begin l_1 = +3;
				 l_2 = -25; end
		6899: begin l_1 = -3;
				 l_2 = +25; end
		11706: begin l_1 = -3;
				 l_2 = -25; end
		13810: begin l_1 = +3;
				 l_2 = +26; end
		4811: begin l_1 = +3;
				 l_2 = -26; end
		13802: begin l_1 = -3;
				 l_2 = +26; end
		4803: begin l_1 = -3;
				 l_2 = -26; end
		9003: begin l_1 = +3;
				 l_2 = +27; end
		9618: begin l_1 = +3;
				 l_2 = -27; end
		8995: begin l_1 = -3;
				 l_2 = +27; end
		9610: begin l_1 = -3;
				 l_2 = -27; end
		18002: begin l_1 = +3;
				 l_2 = +28; end
		619: begin l_1 = +3;
				 l_2 = -28; end
		17994: begin l_1 = -3;
				 l_2 = +28; end
		611: begin l_1 = -3;
				 l_2 = -28; end
		17387: begin l_1 = +3;
				 l_2 = +29; end
		1234: begin l_1 = +3;
				 l_2 = -29; end
		17379: begin l_1 = -3;
				 l_2 = +29; end
		1226: begin l_1 = -3;
				 l_2 = -29; end
		16157: begin l_1 = +3;
				 l_2 = +30; end
		2464: begin l_1 = +3;
				 l_2 = -30; end
		16149: begin l_1 = -3;
				 l_2 = +30; end
		2456: begin l_1 = -3;
				 l_2 = -30; end
		13697: begin l_1 = +3;
				 l_2 = +31; end
		4924: begin l_1 = +3;
				 l_2 = -31; end
		13689: begin l_1 = -3;
				 l_2 = +31; end
		4916: begin l_1 = -3;
				 l_2 = -31; end
		8777: begin l_1 = +3;
				 l_2 = +32; end
		9844: begin l_1 = +3;
				 l_2 = -32; end
		8769: begin l_1 = -3;
				 l_2 = +32; end
		9836: begin l_1 = -3;
				 l_2 = -32; end
		17550: begin l_1 = +3;
				 l_2 = +33; end
		1071: begin l_1 = +3;
				 l_2 = -33; end
		17542: begin l_1 = -3;
				 l_2 = +33; end
		1063: begin l_1 = -3;
				 l_2 = -33; end
		16483: begin l_1 = +3;
				 l_2 = +34; end
		2138: begin l_1 = +3;
				 l_2 = -34; end
		16475: begin l_1 = -3;
				 l_2 = +34; end
		2130: begin l_1 = -3;
				 l_2 = -34; end
		14349: begin l_1 = +3;
				 l_2 = +35; end
		4272: begin l_1 = +3;
				 l_2 = -35; end
		14341: begin l_1 = -3;
				 l_2 = +35; end
		4264: begin l_1 = -3;
				 l_2 = -35; end
		10081: begin l_1 = +3;
				 l_2 = +36; end
		8540: begin l_1 = +3;
				 l_2 = -36; end
		10073: begin l_1 = -3;
				 l_2 = +36; end
		8532: begin l_1 = -3;
				 l_2 = -36; end
		1545: begin l_1 = +3;
				 l_2 = +37; end
		17076: begin l_1 = +3;
				 l_2 = -37; end
		1537: begin l_1 = -3;
				 l_2 = +37; end
		17068: begin l_1 = -3;
				 l_2 = -37; end
		3086: begin l_1 = +3;
				 l_2 = +38; end
		15535: begin l_1 = +3;
				 l_2 = -38; end
		3078: begin l_1 = -3;
				 l_2 = +38; end
		15527: begin l_1 = -3;
				 l_2 = -38; end
		6168: begin l_1 = +3;
				 l_2 = +39; end
		12453: begin l_1 = +3;
				 l_2 = -39; end
		6160: begin l_1 = -3;
				 l_2 = +39; end
		12445: begin l_1 = -3;
				 l_2 = -39; end
		12332: begin l_1 = +3;
				 l_2 = +40; end
		6289: begin l_1 = +3;
				 l_2 = -40; end
		12324: begin l_1 = -3;
				 l_2 = +40; end
		6281: begin l_1 = -3;
				 l_2 = -40; end
		6047: begin l_1 = +3;
				 l_2 = +41; end
		12574: begin l_1 = +3;
				 l_2 = -41; end
		6039: begin l_1 = -3;
				 l_2 = +41; end
		12566: begin l_1 = -3;
				 l_2 = -41; end
		12090: begin l_1 = +3;
				 l_2 = +42; end
		6531: begin l_1 = +3;
				 l_2 = -42; end
		12082: begin l_1 = -3;
				 l_2 = +42; end
		6523: begin l_1 = -3;
				 l_2 = -42; end
		5563: begin l_1 = +3;
				 l_2 = +43; end
		13058: begin l_1 = +3;
				 l_2 = -43; end
		5555: begin l_1 = -3;
				 l_2 = +43; end
		13050: begin l_1 = -3;
				 l_2 = -43; end
		11122: begin l_1 = +3;
				 l_2 = +44; end
		7499: begin l_1 = +3;
				 l_2 = -44; end
		11114: begin l_1 = -3;
				 l_2 = +44; end
		7491: begin l_1 = -3;
				 l_2 = -44; end
		3627: begin l_1 = +3;
				 l_2 = +45; end
		14994: begin l_1 = +3;
				 l_2 = -45; end
		3619: begin l_1 = -3;
				 l_2 = +45; end
		14986: begin l_1 = -3;
				 l_2 = -45; end
		24: begin l_1 = -4;
				 l_2 = +6; end
		18589: begin l_1 = -4;
				 l_2 = -5; end
		40: begin l_1 = +4;
				 l_2 = +6; end
		18573: begin l_1 = -4;
				 l_2 = -6; end
		72: begin l_1 = +4;
				 l_2 = +7; end
		18557: begin l_1 = +4;
				 l_2 = -7; end
		56: begin l_1 = -4;
				 l_2 = +7; end
		18541: begin l_1 = -4;
				 l_2 = -7; end
		136: begin l_1 = +4;
				 l_2 = +8; end
		18493: begin l_1 = +4;
				 l_2 = -8; end
		120: begin l_1 = -4;
				 l_2 = +8; end
		18477: begin l_1 = -4;
				 l_2 = -8; end
		264: begin l_1 = +4;
				 l_2 = +9; end
		18365: begin l_1 = +4;
				 l_2 = -9; end
		248: begin l_1 = -4;
				 l_2 = +9; end
		18349: begin l_1 = -4;
				 l_2 = -9; end
		520: begin l_1 = +4;
				 l_2 = +10; end
		18109: begin l_1 = +4;
				 l_2 = -10; end
		504: begin l_1 = -4;
				 l_2 = +10; end
		18093: begin l_1 = -4;
				 l_2 = -10; end
		1032: begin l_1 = +4;
				 l_2 = +11; end
		17597: begin l_1 = +4;
				 l_2 = -11; end
		1016: begin l_1 = -4;
				 l_2 = +11; end
		17581: begin l_1 = -4;
				 l_2 = -11; end
		2056: begin l_1 = +4;
				 l_2 = +12; end
		16573: begin l_1 = +4;
				 l_2 = -12; end
		2040: begin l_1 = -4;
				 l_2 = +12; end
		16557: begin l_1 = -4;
				 l_2 = -12; end
		4104: begin l_1 = +4;
				 l_2 = +13; end
		14525: begin l_1 = +4;
				 l_2 = -13; end
		4088: begin l_1 = -4;
				 l_2 = +13; end
		14509: begin l_1 = -4;
				 l_2 = -13; end
		8200: begin l_1 = +4;
				 l_2 = +14; end
		10429: begin l_1 = +4;
				 l_2 = -14; end
		8184: begin l_1 = -4;
				 l_2 = +14; end
		10413: begin l_1 = -4;
				 l_2 = -14; end
		16392: begin l_1 = +4;
				 l_2 = +15; end
		2237: begin l_1 = +4;
				 l_2 = -15; end
		16376: begin l_1 = -4;
				 l_2 = +15; end
		2221: begin l_1 = -4;
				 l_2 = -15; end
		14163: begin l_1 = +4;
				 l_2 = +16; end
		4466: begin l_1 = +4;
				 l_2 = -16; end
		14147: begin l_1 = -4;
				 l_2 = +16; end
		4450: begin l_1 = -4;
				 l_2 = -16; end
		9705: begin l_1 = +4;
				 l_2 = +17; end
		8924: begin l_1 = +4;
				 l_2 = -17; end
		9689: begin l_1 = -4;
				 l_2 = +17; end
		8908: begin l_1 = -4;
				 l_2 = -17; end
		789: begin l_1 = +4;
				 l_2 = +18; end
		17840: begin l_1 = +4;
				 l_2 = -18; end
		773: begin l_1 = -4;
				 l_2 = +18; end
		17824: begin l_1 = -4;
				 l_2 = -18; end
		1570: begin l_1 = +4;
				 l_2 = +19; end
		17059: begin l_1 = +4;
				 l_2 = -19; end
		1554: begin l_1 = -4;
				 l_2 = +19; end
		17043: begin l_1 = -4;
				 l_2 = -19; end
		3132: begin l_1 = +4;
				 l_2 = +20; end
		15497: begin l_1 = +4;
				 l_2 = -20; end
		3116: begin l_1 = -4;
				 l_2 = +20; end
		15481: begin l_1 = -4;
				 l_2 = -20; end
		6256: begin l_1 = +4;
				 l_2 = +21; end
		12373: begin l_1 = +4;
				 l_2 = -21; end
		6240: begin l_1 = -4;
				 l_2 = +21; end
		12357: begin l_1 = -4;
				 l_2 = -21; end
		12504: begin l_1 = +4;
				 l_2 = +22; end
		6125: begin l_1 = +4;
				 l_2 = -22; end
		12488: begin l_1 = -4;
				 l_2 = +22; end
		6109: begin l_1 = -4;
				 l_2 = -22; end
		6387: begin l_1 = +4;
				 l_2 = +23; end
		12242: begin l_1 = +4;
				 l_2 = -23; end
		6371: begin l_1 = -4;
				 l_2 = +23; end
		12226: begin l_1 = -4;
				 l_2 = -23; end
		12766: begin l_1 = +4;
				 l_2 = +24; end
		5863: begin l_1 = +4;
				 l_2 = -24; end
		12750: begin l_1 = -4;
				 l_2 = +24; end
		5847: begin l_1 = -4;
				 l_2 = -24; end
		6911: begin l_1 = +4;
				 l_2 = +25; end
		11718: begin l_1 = +4;
				 l_2 = -25; end
		6895: begin l_1 = -4;
				 l_2 = +25; end
		11702: begin l_1 = -4;
				 l_2 = -25; end
		13814: begin l_1 = +4;
				 l_2 = +26; end
		4815: begin l_1 = +4;
				 l_2 = -26; end
		13798: begin l_1 = -4;
				 l_2 = +26; end
		4799: begin l_1 = -4;
				 l_2 = -26; end
		9007: begin l_1 = +4;
				 l_2 = +27; end
		9622: begin l_1 = +4;
				 l_2 = -27; end
		8991: begin l_1 = -4;
				 l_2 = +27; end
		9606: begin l_1 = -4;
				 l_2 = -27; end
		18006: begin l_1 = +4;
				 l_2 = +28; end
		623: begin l_1 = +4;
				 l_2 = -28; end
		17990: begin l_1 = -4;
				 l_2 = +28; end
		607: begin l_1 = -4;
				 l_2 = -28; end
		17391: begin l_1 = +4;
				 l_2 = +29; end
		1238: begin l_1 = +4;
				 l_2 = -29; end
		17375: begin l_1 = -4;
				 l_2 = +29; end
		1222: begin l_1 = -4;
				 l_2 = -29; end
		16161: begin l_1 = +4;
				 l_2 = +30; end
		2468: begin l_1 = +4;
				 l_2 = -30; end
		16145: begin l_1 = -4;
				 l_2 = +30; end
		2452: begin l_1 = -4;
				 l_2 = -30; end
		13701: begin l_1 = +4;
				 l_2 = +31; end
		4928: begin l_1 = +4;
				 l_2 = -31; end
		13685: begin l_1 = -4;
				 l_2 = +31; end
		4912: begin l_1 = -4;
				 l_2 = -31; end
		8781: begin l_1 = +4;
				 l_2 = +32; end
		9848: begin l_1 = +4;
				 l_2 = -32; end
		8765: begin l_1 = -4;
				 l_2 = +32; end
		9832: begin l_1 = -4;
				 l_2 = -32; end
		17554: begin l_1 = +4;
				 l_2 = +33; end
		1075: begin l_1 = +4;
				 l_2 = -33; end
		17538: begin l_1 = -4;
				 l_2 = +33; end
		1059: begin l_1 = -4;
				 l_2 = -33; end
		16487: begin l_1 = +4;
				 l_2 = +34; end
		2142: begin l_1 = +4;
				 l_2 = -34; end
		16471: begin l_1 = -4;
				 l_2 = +34; end
		2126: begin l_1 = -4;
				 l_2 = -34; end
		14353: begin l_1 = +4;
				 l_2 = +35; end
		4276: begin l_1 = +4;
				 l_2 = -35; end
		14337: begin l_1 = -4;
				 l_2 = +35; end
		4260: begin l_1 = -4;
				 l_2 = -35; end
		10085: begin l_1 = +4;
				 l_2 = +36; end
		8544: begin l_1 = +4;
				 l_2 = -36; end
		10069: begin l_1 = -4;
				 l_2 = +36; end
		8528: begin l_1 = -4;
				 l_2 = -36; end
		1549: begin l_1 = +4;
				 l_2 = +37; end
		17080: begin l_1 = +4;
				 l_2 = -37; end
		1533: begin l_1 = -4;
				 l_2 = +37; end
		17064: begin l_1 = -4;
				 l_2 = -37; end
		3090: begin l_1 = +4;
				 l_2 = +38; end
		15539: begin l_1 = +4;
				 l_2 = -38; end
		3074: begin l_1 = -4;
				 l_2 = +38; end
		15523: begin l_1 = -4;
				 l_2 = -38; end
		6172: begin l_1 = +4;
				 l_2 = +39; end
		12457: begin l_1 = +4;
				 l_2 = -39; end
		6156: begin l_1 = -4;
				 l_2 = +39; end
		12441: begin l_1 = -4;
				 l_2 = -39; end
		12336: begin l_1 = +4;
				 l_2 = +40; end
		6293: begin l_1 = +4;
				 l_2 = -40; end
		12320: begin l_1 = -4;
				 l_2 = +40; end
		6277: begin l_1 = -4;
				 l_2 = -40; end
		6051: begin l_1 = +4;
				 l_2 = +41; end
		12578: begin l_1 = +4;
				 l_2 = -41; end
		6035: begin l_1 = -4;
				 l_2 = +41; end
		12562: begin l_1 = -4;
				 l_2 = -41; end
		12094: begin l_1 = +4;
				 l_2 = +42; end
		6535: begin l_1 = +4;
				 l_2 = -42; end
		12078: begin l_1 = -4;
				 l_2 = +42; end
		6519: begin l_1 = -4;
				 l_2 = -42; end
		5567: begin l_1 = +4;
				 l_2 = +43; end
		13062: begin l_1 = +4;
				 l_2 = -43; end
		5551: begin l_1 = -4;
				 l_2 = +43; end
		13046: begin l_1 = -4;
				 l_2 = -43; end
		11126: begin l_1 = +4;
				 l_2 = +44; end
		7503: begin l_1 = +4;
				 l_2 = -44; end
		11110: begin l_1 = -4;
				 l_2 = +44; end
		7487: begin l_1 = -4;
				 l_2 = -44; end
		3631: begin l_1 = +4;
				 l_2 = +45; end
		14998: begin l_1 = +4;
				 l_2 = -45; end
		3615: begin l_1 = -4;
				 l_2 = +45; end
		14982: begin l_1 = -4;
				 l_2 = -45; end
		48: begin l_1 = -5;
				 l_2 = +7; end
		18565: begin l_1 = -5;
				 l_2 = -6; end
		80: begin l_1 = +5;
				 l_2 = +7; end
		18533: begin l_1 = -5;
				 l_2 = -7; end
		144: begin l_1 = +5;
				 l_2 = +8; end
		18501: begin l_1 = +5;
				 l_2 = -8; end
		112: begin l_1 = -5;
				 l_2 = +8; end
		18469: begin l_1 = -5;
				 l_2 = -8; end
		272: begin l_1 = +5;
				 l_2 = +9; end
		18373: begin l_1 = +5;
				 l_2 = -9; end
		240: begin l_1 = -5;
				 l_2 = +9; end
		18341: begin l_1 = -5;
				 l_2 = -9; end
		528: begin l_1 = +5;
				 l_2 = +10; end
		18117: begin l_1 = +5;
				 l_2 = -10; end
		496: begin l_1 = -5;
				 l_2 = +10; end
		18085: begin l_1 = -5;
				 l_2 = -10; end
		1040: begin l_1 = +5;
				 l_2 = +11; end
		17605: begin l_1 = +5;
				 l_2 = -11; end
		1008: begin l_1 = -5;
				 l_2 = +11; end
		17573: begin l_1 = -5;
				 l_2 = -11; end
		2064: begin l_1 = +5;
				 l_2 = +12; end
		16581: begin l_1 = +5;
				 l_2 = -12; end
		2032: begin l_1 = -5;
				 l_2 = +12; end
		16549: begin l_1 = -5;
				 l_2 = -12; end
		4112: begin l_1 = +5;
				 l_2 = +13; end
		14533: begin l_1 = +5;
				 l_2 = -13; end
		4080: begin l_1 = -5;
				 l_2 = +13; end
		14501: begin l_1 = -5;
				 l_2 = -13; end
		8208: begin l_1 = +5;
				 l_2 = +14; end
		10437: begin l_1 = +5;
				 l_2 = -14; end
		8176: begin l_1 = -5;
				 l_2 = +14; end
		10405: begin l_1 = -5;
				 l_2 = -14; end
		16400: begin l_1 = +5;
				 l_2 = +15; end
		2245: begin l_1 = +5;
				 l_2 = -15; end
		16368: begin l_1 = -5;
				 l_2 = +15; end
		2213: begin l_1 = -5;
				 l_2 = -15; end
		14171: begin l_1 = +5;
				 l_2 = +16; end
		4474: begin l_1 = +5;
				 l_2 = -16; end
		14139: begin l_1 = -5;
				 l_2 = +16; end
		4442: begin l_1 = -5;
				 l_2 = -16; end
		9713: begin l_1 = +5;
				 l_2 = +17; end
		8932: begin l_1 = +5;
				 l_2 = -17; end
		9681: begin l_1 = -5;
				 l_2 = +17; end
		8900: begin l_1 = -5;
				 l_2 = -17; end
		797: begin l_1 = +5;
				 l_2 = +18; end
		17848: begin l_1 = +5;
				 l_2 = -18; end
		765: begin l_1 = -5;
				 l_2 = +18; end
		17816: begin l_1 = -5;
				 l_2 = -18; end
		1578: begin l_1 = +5;
				 l_2 = +19; end
		17067: begin l_1 = +5;
				 l_2 = -19; end
		1546: begin l_1 = -5;
				 l_2 = +19; end
		17035: begin l_1 = -5;
				 l_2 = -19; end
		3140: begin l_1 = +5;
				 l_2 = +20; end
		15505: begin l_1 = +5;
				 l_2 = -20; end
		3108: begin l_1 = -5;
				 l_2 = +20; end
		15473: begin l_1 = -5;
				 l_2 = -20; end
		6264: begin l_1 = +5;
				 l_2 = +21; end
		12381: begin l_1 = +5;
				 l_2 = -21; end
		6232: begin l_1 = -5;
				 l_2 = +21; end
		12349: begin l_1 = -5;
				 l_2 = -21; end
		12512: begin l_1 = +5;
				 l_2 = +22; end
		6133: begin l_1 = +5;
				 l_2 = -22; end
		12480: begin l_1 = -5;
				 l_2 = +22; end
		6101: begin l_1 = -5;
				 l_2 = -22; end
		6395: begin l_1 = +5;
				 l_2 = +23; end
		12250: begin l_1 = +5;
				 l_2 = -23; end
		6363: begin l_1 = -5;
				 l_2 = +23; end
		12218: begin l_1 = -5;
				 l_2 = -23; end
		12774: begin l_1 = +5;
				 l_2 = +24; end
		5871: begin l_1 = +5;
				 l_2 = -24; end
		12742: begin l_1 = -5;
				 l_2 = +24; end
		5839: begin l_1 = -5;
				 l_2 = -24; end
		6919: begin l_1 = +5;
				 l_2 = +25; end
		11726: begin l_1 = +5;
				 l_2 = -25; end
		6887: begin l_1 = -5;
				 l_2 = +25; end
		11694: begin l_1 = -5;
				 l_2 = -25; end
		13822: begin l_1 = +5;
				 l_2 = +26; end
		4823: begin l_1 = +5;
				 l_2 = -26; end
		13790: begin l_1 = -5;
				 l_2 = +26; end
		4791: begin l_1 = -5;
				 l_2 = -26; end
		9015: begin l_1 = +5;
				 l_2 = +27; end
		9630: begin l_1 = +5;
				 l_2 = -27; end
		8983: begin l_1 = -5;
				 l_2 = +27; end
		9598: begin l_1 = -5;
				 l_2 = -27; end
		18014: begin l_1 = +5;
				 l_2 = +28; end
		631: begin l_1 = +5;
				 l_2 = -28; end
		17982: begin l_1 = -5;
				 l_2 = +28; end
		599: begin l_1 = -5;
				 l_2 = -28; end
		17399: begin l_1 = +5;
				 l_2 = +29; end
		1246: begin l_1 = +5;
				 l_2 = -29; end
		17367: begin l_1 = -5;
				 l_2 = +29; end
		1214: begin l_1 = -5;
				 l_2 = -29; end
		16169: begin l_1 = +5;
				 l_2 = +30; end
		2476: begin l_1 = +5;
				 l_2 = -30; end
		16137: begin l_1 = -5;
				 l_2 = +30; end
		2444: begin l_1 = -5;
				 l_2 = -30; end
		13709: begin l_1 = +5;
				 l_2 = +31; end
		4936: begin l_1 = +5;
				 l_2 = -31; end
		13677: begin l_1 = -5;
				 l_2 = +31; end
		4904: begin l_1 = -5;
				 l_2 = -31; end
		8789: begin l_1 = +5;
				 l_2 = +32; end
		9856: begin l_1 = +5;
				 l_2 = -32; end
		8757: begin l_1 = -5;
				 l_2 = +32; end
		9824: begin l_1 = -5;
				 l_2 = -32; end
		17562: begin l_1 = +5;
				 l_2 = +33; end
		1083: begin l_1 = +5;
				 l_2 = -33; end
		17530: begin l_1 = -5;
				 l_2 = +33; end
		1051: begin l_1 = -5;
				 l_2 = -33; end
		16495: begin l_1 = +5;
				 l_2 = +34; end
		2150: begin l_1 = +5;
				 l_2 = -34; end
		16463: begin l_1 = -5;
				 l_2 = +34; end
		2118: begin l_1 = -5;
				 l_2 = -34; end
		14361: begin l_1 = +5;
				 l_2 = +35; end
		4284: begin l_1 = +5;
				 l_2 = -35; end
		14329: begin l_1 = -5;
				 l_2 = +35; end
		4252: begin l_1 = -5;
				 l_2 = -35; end
		10093: begin l_1 = +5;
				 l_2 = +36; end
		8552: begin l_1 = +5;
				 l_2 = -36; end
		10061: begin l_1 = -5;
				 l_2 = +36; end
		8520: begin l_1 = -5;
				 l_2 = -36; end
		1557: begin l_1 = +5;
				 l_2 = +37; end
		17088: begin l_1 = +5;
				 l_2 = -37; end
		1525: begin l_1 = -5;
				 l_2 = +37; end
		17056: begin l_1 = -5;
				 l_2 = -37; end
		3098: begin l_1 = +5;
				 l_2 = +38; end
		15547: begin l_1 = +5;
				 l_2 = -38; end
		3066: begin l_1 = -5;
				 l_2 = +38; end
		15515: begin l_1 = -5;
				 l_2 = -38; end
		6180: begin l_1 = +5;
				 l_2 = +39; end
		12465: begin l_1 = +5;
				 l_2 = -39; end
		6148: begin l_1 = -5;
				 l_2 = +39; end
		12433: begin l_1 = -5;
				 l_2 = -39; end
		12344: begin l_1 = +5;
				 l_2 = +40; end
		6301: begin l_1 = +5;
				 l_2 = -40; end
		12312: begin l_1 = -5;
				 l_2 = +40; end
		6269: begin l_1 = -5;
				 l_2 = -40; end
		6059: begin l_1 = +5;
				 l_2 = +41; end
		12586: begin l_1 = +5;
				 l_2 = -41; end
		6027: begin l_1 = -5;
				 l_2 = +41; end
		12554: begin l_1 = -5;
				 l_2 = -41; end
		12102: begin l_1 = +5;
				 l_2 = +42; end
		6543: begin l_1 = +5;
				 l_2 = -42; end
		12070: begin l_1 = -5;
				 l_2 = +42; end
		6511: begin l_1 = -5;
				 l_2 = -42; end
		5575: begin l_1 = +5;
				 l_2 = +43; end
		13070: begin l_1 = +5;
				 l_2 = -43; end
		5543: begin l_1 = -5;
				 l_2 = +43; end
		13038: begin l_1 = -5;
				 l_2 = -43; end
		11134: begin l_1 = +5;
				 l_2 = +44; end
		7511: begin l_1 = +5;
				 l_2 = -44; end
		11102: begin l_1 = -5;
				 l_2 = +44; end
		7479: begin l_1 = -5;
				 l_2 = -44; end
		3639: begin l_1 = +5;
				 l_2 = +45; end
		15006: begin l_1 = +5;
				 l_2 = -45; end
		3607: begin l_1 = -5;
				 l_2 = +45; end
		14974: begin l_1 = -5;
				 l_2 = -45; end
		96: begin l_1 = -6;
				 l_2 = +8; end
		18517: begin l_1 = -6;
				 l_2 = -7; end
		160: begin l_1 = +6;
				 l_2 = +8; end
		18453: begin l_1 = -6;
				 l_2 = -8; end
		288: begin l_1 = +6;
				 l_2 = +9; end
		18389: begin l_1 = +6;
				 l_2 = -9; end
		224: begin l_1 = -6;
				 l_2 = +9; end
		18325: begin l_1 = -6;
				 l_2 = -9; end
		544: begin l_1 = +6;
				 l_2 = +10; end
		18133: begin l_1 = +6;
				 l_2 = -10; end
		480: begin l_1 = -6;
				 l_2 = +10; end
		18069: begin l_1 = -6;
				 l_2 = -10; end
		1056: begin l_1 = +6;
				 l_2 = +11; end
		17621: begin l_1 = +6;
				 l_2 = -11; end
		992: begin l_1 = -6;
				 l_2 = +11; end
		17557: begin l_1 = -6;
				 l_2 = -11; end
		2080: begin l_1 = +6;
				 l_2 = +12; end
		16597: begin l_1 = +6;
				 l_2 = -12; end
		2016: begin l_1 = -6;
				 l_2 = +12; end
		16533: begin l_1 = -6;
				 l_2 = -12; end
		4128: begin l_1 = +6;
				 l_2 = +13; end
		14549: begin l_1 = +6;
				 l_2 = -13; end
		4064: begin l_1 = -6;
				 l_2 = +13; end
		14485: begin l_1 = -6;
				 l_2 = -13; end
		8224: begin l_1 = +6;
				 l_2 = +14; end
		10453: begin l_1 = +6;
				 l_2 = -14; end
		8160: begin l_1 = -6;
				 l_2 = +14; end
		10389: begin l_1 = -6;
				 l_2 = -14; end
		16416: begin l_1 = +6;
				 l_2 = +15; end
		2261: begin l_1 = +6;
				 l_2 = -15; end
		16352: begin l_1 = -6;
				 l_2 = +15; end
		2197: begin l_1 = -6;
				 l_2 = -15; end
		14187: begin l_1 = +6;
				 l_2 = +16; end
		4490: begin l_1 = +6;
				 l_2 = -16; end
		14123: begin l_1 = -6;
				 l_2 = +16; end
		4426: begin l_1 = -6;
				 l_2 = -16; end
		9729: begin l_1 = +6;
				 l_2 = +17; end
		8948: begin l_1 = +6;
				 l_2 = -17; end
		9665: begin l_1 = -6;
				 l_2 = +17; end
		8884: begin l_1 = -6;
				 l_2 = -17; end
		813: begin l_1 = +6;
				 l_2 = +18; end
		17864: begin l_1 = +6;
				 l_2 = -18; end
		749: begin l_1 = -6;
				 l_2 = +18; end
		17800: begin l_1 = -6;
				 l_2 = -18; end
		1594: begin l_1 = +6;
				 l_2 = +19; end
		17083: begin l_1 = +6;
				 l_2 = -19; end
		1530: begin l_1 = -6;
				 l_2 = +19; end
		17019: begin l_1 = -6;
				 l_2 = -19; end
		3156: begin l_1 = +6;
				 l_2 = +20; end
		15521: begin l_1 = +6;
				 l_2 = -20; end
		3092: begin l_1 = -6;
				 l_2 = +20; end
		15457: begin l_1 = -6;
				 l_2 = -20; end
		6280: begin l_1 = +6;
				 l_2 = +21; end
		12397: begin l_1 = +6;
				 l_2 = -21; end
		6216: begin l_1 = -6;
				 l_2 = +21; end
		12333: begin l_1 = -6;
				 l_2 = -21; end
		12528: begin l_1 = +6;
				 l_2 = +22; end
		6149: begin l_1 = +6;
				 l_2 = -22; end
		12464: begin l_1 = -6;
				 l_2 = +22; end
		6085: begin l_1 = -6;
				 l_2 = -22; end
		6411: begin l_1 = +6;
				 l_2 = +23; end
		12266: begin l_1 = +6;
				 l_2 = -23; end
		6347: begin l_1 = -6;
				 l_2 = +23; end
		12202: begin l_1 = -6;
				 l_2 = -23; end
		12790: begin l_1 = +6;
				 l_2 = +24; end
		5887: begin l_1 = +6;
				 l_2 = -24; end
		12726: begin l_1 = -6;
				 l_2 = +24; end
		5823: begin l_1 = -6;
				 l_2 = -24; end
		6935: begin l_1 = +6;
				 l_2 = +25; end
		11742: begin l_1 = +6;
				 l_2 = -25; end
		6871: begin l_1 = -6;
				 l_2 = +25; end
		11678: begin l_1 = -6;
				 l_2 = -25; end
		13838: begin l_1 = +6;
				 l_2 = +26; end
		4839: begin l_1 = +6;
				 l_2 = -26; end
		13774: begin l_1 = -6;
				 l_2 = +26; end
		4775: begin l_1 = -6;
				 l_2 = -26; end
		9031: begin l_1 = +6;
				 l_2 = +27; end
		9646: begin l_1 = +6;
				 l_2 = -27; end
		8967: begin l_1 = -6;
				 l_2 = +27; end
		9582: begin l_1 = -6;
				 l_2 = -27; end
		18030: begin l_1 = +6;
				 l_2 = +28; end
		647: begin l_1 = +6;
				 l_2 = -28; end
		17966: begin l_1 = -6;
				 l_2 = +28; end
		583: begin l_1 = -6;
				 l_2 = -28; end
		17415: begin l_1 = +6;
				 l_2 = +29; end
		1262: begin l_1 = +6;
				 l_2 = -29; end
		17351: begin l_1 = -6;
				 l_2 = +29; end
		1198: begin l_1 = -6;
				 l_2 = -29; end
		16185: begin l_1 = +6;
				 l_2 = +30; end
		2492: begin l_1 = +6;
				 l_2 = -30; end
		16121: begin l_1 = -6;
				 l_2 = +30; end
		2428: begin l_1 = -6;
				 l_2 = -30; end
		13725: begin l_1 = +6;
				 l_2 = +31; end
		4952: begin l_1 = +6;
				 l_2 = -31; end
		13661: begin l_1 = -6;
				 l_2 = +31; end
		4888: begin l_1 = -6;
				 l_2 = -31; end
		8805: begin l_1 = +6;
				 l_2 = +32; end
		9872: begin l_1 = +6;
				 l_2 = -32; end
		8741: begin l_1 = -6;
				 l_2 = +32; end
		9808: begin l_1 = -6;
				 l_2 = -32; end
		17578: begin l_1 = +6;
				 l_2 = +33; end
		1099: begin l_1 = +6;
				 l_2 = -33; end
		17514: begin l_1 = -6;
				 l_2 = +33; end
		1035: begin l_1 = -6;
				 l_2 = -33; end
		16511: begin l_1 = +6;
				 l_2 = +34; end
		2166: begin l_1 = +6;
				 l_2 = -34; end
		16447: begin l_1 = -6;
				 l_2 = +34; end
		2102: begin l_1 = -6;
				 l_2 = -34; end
		14377: begin l_1 = +6;
				 l_2 = +35; end
		4300: begin l_1 = +6;
				 l_2 = -35; end
		14313: begin l_1 = -6;
				 l_2 = +35; end
		4236: begin l_1 = -6;
				 l_2 = -35; end
		10109: begin l_1 = +6;
				 l_2 = +36; end
		8568: begin l_1 = +6;
				 l_2 = -36; end
		10045: begin l_1 = -6;
				 l_2 = +36; end
		8504: begin l_1 = -6;
				 l_2 = -36; end
		1573: begin l_1 = +6;
				 l_2 = +37; end
		17104: begin l_1 = +6;
				 l_2 = -37; end
		1509: begin l_1 = -6;
				 l_2 = +37; end
		17040: begin l_1 = -6;
				 l_2 = -37; end
		3114: begin l_1 = +6;
				 l_2 = +38; end
		15563: begin l_1 = +6;
				 l_2 = -38; end
		3050: begin l_1 = -6;
				 l_2 = +38; end
		15499: begin l_1 = -6;
				 l_2 = -38; end
		6196: begin l_1 = +6;
				 l_2 = +39; end
		12481: begin l_1 = +6;
				 l_2 = -39; end
		6132: begin l_1 = -6;
				 l_2 = +39; end
		12417: begin l_1 = -6;
				 l_2 = -39; end
		12360: begin l_1 = +6;
				 l_2 = +40; end
		6317: begin l_1 = +6;
				 l_2 = -40; end
		12296: begin l_1 = -6;
				 l_2 = +40; end
		6253: begin l_1 = -6;
				 l_2 = -40; end
		6075: begin l_1 = +6;
				 l_2 = +41; end
		12602: begin l_1 = +6;
				 l_2 = -41; end
		6011: begin l_1 = -6;
				 l_2 = +41; end
		12538: begin l_1 = -6;
				 l_2 = -41; end
		12118: begin l_1 = +6;
				 l_2 = +42; end
		6559: begin l_1 = +6;
				 l_2 = -42; end
		12054: begin l_1 = -6;
				 l_2 = +42; end
		6495: begin l_1 = -6;
				 l_2 = -42; end
		5591: begin l_1 = +6;
				 l_2 = +43; end
		13086: begin l_1 = +6;
				 l_2 = -43; end
		5527: begin l_1 = -6;
				 l_2 = +43; end
		13022: begin l_1 = -6;
				 l_2 = -43; end
		11150: begin l_1 = +6;
				 l_2 = +44; end
		7527: begin l_1 = +6;
				 l_2 = -44; end
		11086: begin l_1 = -6;
				 l_2 = +44; end
		7463: begin l_1 = -6;
				 l_2 = -44; end
		3655: begin l_1 = +6;
				 l_2 = +45; end
		15022: begin l_1 = +6;
				 l_2 = -45; end
		3591: begin l_1 = -6;
				 l_2 = +45; end
		14958: begin l_1 = -6;
				 l_2 = -45; end
		192: begin l_1 = -7;
				 l_2 = +9; end
		18421: begin l_1 = -7;
				 l_2 = -8; end
		320: begin l_1 = +7;
				 l_2 = +9; end
		18293: begin l_1 = -7;
				 l_2 = -9; end
		576: begin l_1 = +7;
				 l_2 = +10; end
		18165: begin l_1 = +7;
				 l_2 = -10; end
		448: begin l_1 = -7;
				 l_2 = +10; end
		18037: begin l_1 = -7;
				 l_2 = -10; end
		1088: begin l_1 = +7;
				 l_2 = +11; end
		17653: begin l_1 = +7;
				 l_2 = -11; end
		960: begin l_1 = -7;
				 l_2 = +11; end
		17525: begin l_1 = -7;
				 l_2 = -11; end
		2112: begin l_1 = +7;
				 l_2 = +12; end
		16629: begin l_1 = +7;
				 l_2 = -12; end
		1984: begin l_1 = -7;
				 l_2 = +12; end
		16501: begin l_1 = -7;
				 l_2 = -12; end
		4160: begin l_1 = +7;
				 l_2 = +13; end
		14581: begin l_1 = +7;
				 l_2 = -13; end
		4032: begin l_1 = -7;
				 l_2 = +13; end
		14453: begin l_1 = -7;
				 l_2 = -13; end
		8256: begin l_1 = +7;
				 l_2 = +14; end
		10485: begin l_1 = +7;
				 l_2 = -14; end
		8128: begin l_1 = -7;
				 l_2 = +14; end
		10357: begin l_1 = -7;
				 l_2 = -14; end
		16448: begin l_1 = +7;
				 l_2 = +15; end
		2293: begin l_1 = +7;
				 l_2 = -15; end
		16320: begin l_1 = -7;
				 l_2 = +15; end
		2165: begin l_1 = -7;
				 l_2 = -15; end
		14219: begin l_1 = +7;
				 l_2 = +16; end
		4522: begin l_1 = +7;
				 l_2 = -16; end
		14091: begin l_1 = -7;
				 l_2 = +16; end
		4394: begin l_1 = -7;
				 l_2 = -16; end
		9761: begin l_1 = +7;
				 l_2 = +17; end
		8980: begin l_1 = +7;
				 l_2 = -17; end
		9633: begin l_1 = -7;
				 l_2 = +17; end
		8852: begin l_1 = -7;
				 l_2 = -17; end
		845: begin l_1 = +7;
				 l_2 = +18; end
		17896: begin l_1 = +7;
				 l_2 = -18; end
		717: begin l_1 = -7;
				 l_2 = +18; end
		17768: begin l_1 = -7;
				 l_2 = -18; end
		1626: begin l_1 = +7;
				 l_2 = +19; end
		17115: begin l_1 = +7;
				 l_2 = -19; end
		1498: begin l_1 = -7;
				 l_2 = +19; end
		16987: begin l_1 = -7;
				 l_2 = -19; end
		3188: begin l_1 = +7;
				 l_2 = +20; end
		15553: begin l_1 = +7;
				 l_2 = -20; end
		3060: begin l_1 = -7;
				 l_2 = +20; end
		15425: begin l_1 = -7;
				 l_2 = -20; end
		6312: begin l_1 = +7;
				 l_2 = +21; end
		12429: begin l_1 = +7;
				 l_2 = -21; end
		6184: begin l_1 = -7;
				 l_2 = +21; end
		12301: begin l_1 = -7;
				 l_2 = -21; end
		12560: begin l_1 = +7;
				 l_2 = +22; end
		6181: begin l_1 = +7;
				 l_2 = -22; end
		12432: begin l_1 = -7;
				 l_2 = +22; end
		6053: begin l_1 = -7;
				 l_2 = -22; end
		6443: begin l_1 = +7;
				 l_2 = +23; end
		12298: begin l_1 = +7;
				 l_2 = -23; end
		6315: begin l_1 = -7;
				 l_2 = +23; end
		12170: begin l_1 = -7;
				 l_2 = -23; end
		12822: begin l_1 = +7;
				 l_2 = +24; end
		5919: begin l_1 = +7;
				 l_2 = -24; end
		12694: begin l_1 = -7;
				 l_2 = +24; end
		5791: begin l_1 = -7;
				 l_2 = -24; end
		6967: begin l_1 = +7;
				 l_2 = +25; end
		11774: begin l_1 = +7;
				 l_2 = -25; end
		6839: begin l_1 = -7;
				 l_2 = +25; end
		11646: begin l_1 = -7;
				 l_2 = -25; end
		13870: begin l_1 = +7;
				 l_2 = +26; end
		4871: begin l_1 = +7;
				 l_2 = -26; end
		13742: begin l_1 = -7;
				 l_2 = +26; end
		4743: begin l_1 = -7;
				 l_2 = -26; end
		9063: begin l_1 = +7;
				 l_2 = +27; end
		9678: begin l_1 = +7;
				 l_2 = -27; end
		8935: begin l_1 = -7;
				 l_2 = +27; end
		9550: begin l_1 = -7;
				 l_2 = -27; end
		18062: begin l_1 = +7;
				 l_2 = +28; end
		679: begin l_1 = +7;
				 l_2 = -28; end
		17934: begin l_1 = -7;
				 l_2 = +28; end
		551: begin l_1 = -7;
				 l_2 = -28; end
		17447: begin l_1 = +7;
				 l_2 = +29; end
		1294: begin l_1 = +7;
				 l_2 = -29; end
		17319: begin l_1 = -7;
				 l_2 = +29; end
		1166: begin l_1 = -7;
				 l_2 = -29; end
		16217: begin l_1 = +7;
				 l_2 = +30; end
		2524: begin l_1 = +7;
				 l_2 = -30; end
		16089: begin l_1 = -7;
				 l_2 = +30; end
		2396: begin l_1 = -7;
				 l_2 = -30; end
		13757: begin l_1 = +7;
				 l_2 = +31; end
		4984: begin l_1 = +7;
				 l_2 = -31; end
		13629: begin l_1 = -7;
				 l_2 = +31; end
		4856: begin l_1 = -7;
				 l_2 = -31; end
		8837: begin l_1 = +7;
				 l_2 = +32; end
		9904: begin l_1 = +7;
				 l_2 = -32; end
		8709: begin l_1 = -7;
				 l_2 = +32; end
		9776: begin l_1 = -7;
				 l_2 = -32; end
		17610: begin l_1 = +7;
				 l_2 = +33; end
		1131: begin l_1 = +7;
				 l_2 = -33; end
		17482: begin l_1 = -7;
				 l_2 = +33; end
		1003: begin l_1 = -7;
				 l_2 = -33; end
		16543: begin l_1 = +7;
				 l_2 = +34; end
		2198: begin l_1 = +7;
				 l_2 = -34; end
		16415: begin l_1 = -7;
				 l_2 = +34; end
		2070: begin l_1 = -7;
				 l_2 = -34; end
		14409: begin l_1 = +7;
				 l_2 = +35; end
		4332: begin l_1 = +7;
				 l_2 = -35; end
		14281: begin l_1 = -7;
				 l_2 = +35; end
		4204: begin l_1 = -7;
				 l_2 = -35; end
		10141: begin l_1 = +7;
				 l_2 = +36; end
		8600: begin l_1 = +7;
				 l_2 = -36; end
		10013: begin l_1 = -7;
				 l_2 = +36; end
		8472: begin l_1 = -7;
				 l_2 = -36; end
		1605: begin l_1 = +7;
				 l_2 = +37; end
		17136: begin l_1 = +7;
				 l_2 = -37; end
		1477: begin l_1 = -7;
				 l_2 = +37; end
		17008: begin l_1 = -7;
				 l_2 = -37; end
		3146: begin l_1 = +7;
				 l_2 = +38; end
		15595: begin l_1 = +7;
				 l_2 = -38; end
		3018: begin l_1 = -7;
				 l_2 = +38; end
		15467: begin l_1 = -7;
				 l_2 = -38; end
		6228: begin l_1 = +7;
				 l_2 = +39; end
		12513: begin l_1 = +7;
				 l_2 = -39; end
		6100: begin l_1 = -7;
				 l_2 = +39; end
		12385: begin l_1 = -7;
				 l_2 = -39; end
		12392: begin l_1 = +7;
				 l_2 = +40; end
		6349: begin l_1 = +7;
				 l_2 = -40; end
		12264: begin l_1 = -7;
				 l_2 = +40; end
		6221: begin l_1 = -7;
				 l_2 = -40; end
		6107: begin l_1 = +7;
				 l_2 = +41; end
		12634: begin l_1 = +7;
				 l_2 = -41; end
		5979: begin l_1 = -7;
				 l_2 = +41; end
		12506: begin l_1 = -7;
				 l_2 = -41; end
		12150: begin l_1 = +7;
				 l_2 = +42; end
		6591: begin l_1 = +7;
				 l_2 = -42; end
		12022: begin l_1 = -7;
				 l_2 = +42; end
		6463: begin l_1 = -7;
				 l_2 = -42; end
		5623: begin l_1 = +7;
				 l_2 = +43; end
		13118: begin l_1 = +7;
				 l_2 = -43; end
		5495: begin l_1 = -7;
				 l_2 = +43; end
		12990: begin l_1 = -7;
				 l_2 = -43; end
		11182: begin l_1 = +7;
				 l_2 = +44; end
		7559: begin l_1 = +7;
				 l_2 = -44; end
		11054: begin l_1 = -7;
				 l_2 = +44; end
		7431: begin l_1 = -7;
				 l_2 = -44; end
		3687: begin l_1 = +7;
				 l_2 = +45; end
		15054: begin l_1 = +7;
				 l_2 = -45; end
		3559: begin l_1 = -7;
				 l_2 = +45; end
		14926: begin l_1 = -7;
				 l_2 = -45; end
		384: begin l_1 = -8;
				 l_2 = +10; end
		18229: begin l_1 = -8;
				 l_2 = -9; end
		640: begin l_1 = +8;
				 l_2 = +10; end
		17973: begin l_1 = -8;
				 l_2 = -10; end
		1152: begin l_1 = +8;
				 l_2 = +11; end
		17717: begin l_1 = +8;
				 l_2 = -11; end
		896: begin l_1 = -8;
				 l_2 = +11; end
		17461: begin l_1 = -8;
				 l_2 = -11; end
		2176: begin l_1 = +8;
				 l_2 = +12; end
		16693: begin l_1 = +8;
				 l_2 = -12; end
		1920: begin l_1 = -8;
				 l_2 = +12; end
		16437: begin l_1 = -8;
				 l_2 = -12; end
		4224: begin l_1 = +8;
				 l_2 = +13; end
		14645: begin l_1 = +8;
				 l_2 = -13; end
		3968: begin l_1 = -8;
				 l_2 = +13; end
		14389: begin l_1 = -8;
				 l_2 = -13; end
		8320: begin l_1 = +8;
				 l_2 = +14; end
		10549: begin l_1 = +8;
				 l_2 = -14; end
		8064: begin l_1 = -8;
				 l_2 = +14; end
		10293: begin l_1 = -8;
				 l_2 = -14; end
		16512: begin l_1 = +8;
				 l_2 = +15; end
		2357: begin l_1 = +8;
				 l_2 = -15; end
		16256: begin l_1 = -8;
				 l_2 = +15; end
		2101: begin l_1 = -8;
				 l_2 = -15; end
		14283: begin l_1 = +8;
				 l_2 = +16; end
		4586: begin l_1 = +8;
				 l_2 = -16; end
		14027: begin l_1 = -8;
				 l_2 = +16; end
		4330: begin l_1 = -8;
				 l_2 = -16; end
		9825: begin l_1 = +8;
				 l_2 = +17; end
		9044: begin l_1 = +8;
				 l_2 = -17; end
		9569: begin l_1 = -8;
				 l_2 = +17; end
		8788: begin l_1 = -8;
				 l_2 = -17; end
		909: begin l_1 = +8;
				 l_2 = +18; end
		17960: begin l_1 = +8;
				 l_2 = -18; end
		653: begin l_1 = -8;
				 l_2 = +18; end
		17704: begin l_1 = -8;
				 l_2 = -18; end
		1690: begin l_1 = +8;
				 l_2 = +19; end
		17179: begin l_1 = +8;
				 l_2 = -19; end
		1434: begin l_1 = -8;
				 l_2 = +19; end
		16923: begin l_1 = -8;
				 l_2 = -19; end
		3252: begin l_1 = +8;
				 l_2 = +20; end
		15617: begin l_1 = +8;
				 l_2 = -20; end
		2996: begin l_1 = -8;
				 l_2 = +20; end
		15361: begin l_1 = -8;
				 l_2 = -20; end
		6376: begin l_1 = +8;
				 l_2 = +21; end
		12493: begin l_1 = +8;
				 l_2 = -21; end
		6120: begin l_1 = -8;
				 l_2 = +21; end
		12237: begin l_1 = -8;
				 l_2 = -21; end
		12624: begin l_1 = +8;
				 l_2 = +22; end
		6245: begin l_1 = +8;
				 l_2 = -22; end
		12368: begin l_1 = -8;
				 l_2 = +22; end
		5989: begin l_1 = -8;
				 l_2 = -22; end
		6507: begin l_1 = +8;
				 l_2 = +23; end
		12362: begin l_1 = +8;
				 l_2 = -23; end
		6251: begin l_1 = -8;
				 l_2 = +23; end
		12106: begin l_1 = -8;
				 l_2 = -23; end
		12886: begin l_1 = +8;
				 l_2 = +24; end
		5983: begin l_1 = +8;
				 l_2 = -24; end
		12630: begin l_1 = -8;
				 l_2 = +24; end
		5727: begin l_1 = -8;
				 l_2 = -24; end
		7031: begin l_1 = +8;
				 l_2 = +25; end
		11838: begin l_1 = +8;
				 l_2 = -25; end
		6775: begin l_1 = -8;
				 l_2 = +25; end
		11582: begin l_1 = -8;
				 l_2 = -25; end
		13934: begin l_1 = +8;
				 l_2 = +26; end
		4935: begin l_1 = +8;
				 l_2 = -26; end
		13678: begin l_1 = -8;
				 l_2 = +26; end
		4679: begin l_1 = -8;
				 l_2 = -26; end
		9127: begin l_1 = +8;
				 l_2 = +27; end
		9742: begin l_1 = +8;
				 l_2 = -27; end
		8871: begin l_1 = -8;
				 l_2 = +27; end
		9486: begin l_1 = -8;
				 l_2 = -27; end
		18126: begin l_1 = +8;
				 l_2 = +28; end
		743: begin l_1 = +8;
				 l_2 = -28; end
		17870: begin l_1 = -8;
				 l_2 = +28; end
		487: begin l_1 = -8;
				 l_2 = -28; end
		17511: begin l_1 = +8;
				 l_2 = +29; end
		1358: begin l_1 = +8;
				 l_2 = -29; end
		17255: begin l_1 = -8;
				 l_2 = +29; end
		1102: begin l_1 = -8;
				 l_2 = -29; end
		16281: begin l_1 = +8;
				 l_2 = +30; end
		2588: begin l_1 = +8;
				 l_2 = -30; end
		16025: begin l_1 = -8;
				 l_2 = +30; end
		2332: begin l_1 = -8;
				 l_2 = -30; end
		13821: begin l_1 = +8;
				 l_2 = +31; end
		5048: begin l_1 = +8;
				 l_2 = -31; end
		13565: begin l_1 = -8;
				 l_2 = +31; end
		4792: begin l_1 = -8;
				 l_2 = -31; end
		8901: begin l_1 = +8;
				 l_2 = +32; end
		9968: begin l_1 = +8;
				 l_2 = -32; end
		8645: begin l_1 = -8;
				 l_2 = +32; end
		9712: begin l_1 = -8;
				 l_2 = -32; end
		17674: begin l_1 = +8;
				 l_2 = +33; end
		1195: begin l_1 = +8;
				 l_2 = -33; end
		17418: begin l_1 = -8;
				 l_2 = +33; end
		939: begin l_1 = -8;
				 l_2 = -33; end
		16607: begin l_1 = +8;
				 l_2 = +34; end
		2262: begin l_1 = +8;
				 l_2 = -34; end
		16351: begin l_1 = -8;
				 l_2 = +34; end
		2006: begin l_1 = -8;
				 l_2 = -34; end
		14473: begin l_1 = +8;
				 l_2 = +35; end
		4396: begin l_1 = +8;
				 l_2 = -35; end
		14217: begin l_1 = -8;
				 l_2 = +35; end
		4140: begin l_1 = -8;
				 l_2 = -35; end
		10205: begin l_1 = +8;
				 l_2 = +36; end
		8664: begin l_1 = +8;
				 l_2 = -36; end
		9949: begin l_1 = -8;
				 l_2 = +36; end
		8408: begin l_1 = -8;
				 l_2 = -36; end
		1669: begin l_1 = +8;
				 l_2 = +37; end
		17200: begin l_1 = +8;
				 l_2 = -37; end
		1413: begin l_1 = -8;
				 l_2 = +37; end
		16944: begin l_1 = -8;
				 l_2 = -37; end
		3210: begin l_1 = +8;
				 l_2 = +38; end
		15659: begin l_1 = +8;
				 l_2 = -38; end
		2954: begin l_1 = -8;
				 l_2 = +38; end
		15403: begin l_1 = -8;
				 l_2 = -38; end
		6292: begin l_1 = +8;
				 l_2 = +39; end
		12577: begin l_1 = +8;
				 l_2 = -39; end
		6036: begin l_1 = -8;
				 l_2 = +39; end
		12321: begin l_1 = -8;
				 l_2 = -39; end
		12456: begin l_1 = +8;
				 l_2 = +40; end
		6413: begin l_1 = +8;
				 l_2 = -40; end
		12200: begin l_1 = -8;
				 l_2 = +40; end
		6157: begin l_1 = -8;
				 l_2 = -40; end
		6171: begin l_1 = +8;
				 l_2 = +41; end
		12698: begin l_1 = +8;
				 l_2 = -41; end
		5915: begin l_1 = -8;
				 l_2 = +41; end
		12442: begin l_1 = -8;
				 l_2 = -41; end
		12214: begin l_1 = +8;
				 l_2 = +42; end
		6655: begin l_1 = +8;
				 l_2 = -42; end
		11958: begin l_1 = -8;
				 l_2 = +42; end
		6399: begin l_1 = -8;
				 l_2 = -42; end
		5687: begin l_1 = +8;
				 l_2 = +43; end
		13182: begin l_1 = +8;
				 l_2 = -43; end
		5431: begin l_1 = -8;
				 l_2 = +43; end
		12926: begin l_1 = -8;
				 l_2 = -43; end
		11246: begin l_1 = +8;
				 l_2 = +44; end
		7623: begin l_1 = +8;
				 l_2 = -44; end
		10990: begin l_1 = -8;
				 l_2 = +44; end
		7367: begin l_1 = -8;
				 l_2 = -44; end
		3751: begin l_1 = +8;
				 l_2 = +45; end
		15118: begin l_1 = +8;
				 l_2 = -45; end
		3495: begin l_1 = -8;
				 l_2 = +45; end
		14862: begin l_1 = -8;
				 l_2 = -45; end
		768: begin l_1 = -9;
				 l_2 = +11; end
		17845: begin l_1 = -9;
				 l_2 = -10; end
		1280: begin l_1 = +9;
				 l_2 = +11; end
		17333: begin l_1 = -9;
				 l_2 = -11; end
		2304: begin l_1 = +9;
				 l_2 = +12; end
		16821: begin l_1 = +9;
				 l_2 = -12; end
		1792: begin l_1 = -9;
				 l_2 = +12; end
		16309: begin l_1 = -9;
				 l_2 = -12; end
		4352: begin l_1 = +9;
				 l_2 = +13; end
		14773: begin l_1 = +9;
				 l_2 = -13; end
		3840: begin l_1 = -9;
				 l_2 = +13; end
		14261: begin l_1 = -9;
				 l_2 = -13; end
		8448: begin l_1 = +9;
				 l_2 = +14; end
		10677: begin l_1 = +9;
				 l_2 = -14; end
		7936: begin l_1 = -9;
				 l_2 = +14; end
		10165: begin l_1 = -9;
				 l_2 = -14; end
		16640: begin l_1 = +9;
				 l_2 = +15; end
		2485: begin l_1 = +9;
				 l_2 = -15; end
		16128: begin l_1 = -9;
				 l_2 = +15; end
		1973: begin l_1 = -9;
				 l_2 = -15; end
		14411: begin l_1 = +9;
				 l_2 = +16; end
		4714: begin l_1 = +9;
				 l_2 = -16; end
		13899: begin l_1 = -9;
				 l_2 = +16; end
		4202: begin l_1 = -9;
				 l_2 = -16; end
		9953: begin l_1 = +9;
				 l_2 = +17; end
		9172: begin l_1 = +9;
				 l_2 = -17; end
		9441: begin l_1 = -9;
				 l_2 = +17; end
		8660: begin l_1 = -9;
				 l_2 = -17; end
		1037: begin l_1 = +9;
				 l_2 = +18; end
		18088: begin l_1 = +9;
				 l_2 = -18; end
		525: begin l_1 = -9;
				 l_2 = +18; end
		17576: begin l_1 = -9;
				 l_2 = -18; end
		1818: begin l_1 = +9;
				 l_2 = +19; end
		17307: begin l_1 = +9;
				 l_2 = -19; end
		1306: begin l_1 = -9;
				 l_2 = +19; end
		16795: begin l_1 = -9;
				 l_2 = -19; end
		3380: begin l_1 = +9;
				 l_2 = +20; end
		15745: begin l_1 = +9;
				 l_2 = -20; end
		2868: begin l_1 = -9;
				 l_2 = +20; end
		15233: begin l_1 = -9;
				 l_2 = -20; end
		6504: begin l_1 = +9;
				 l_2 = +21; end
		12621: begin l_1 = +9;
				 l_2 = -21; end
		5992: begin l_1 = -9;
				 l_2 = +21; end
		12109: begin l_1 = -9;
				 l_2 = -21; end
		12752: begin l_1 = +9;
				 l_2 = +22; end
		6373: begin l_1 = +9;
				 l_2 = -22; end
		12240: begin l_1 = -9;
				 l_2 = +22; end
		5861: begin l_1 = -9;
				 l_2 = -22; end
		6635: begin l_1 = +9;
				 l_2 = +23; end
		12490: begin l_1 = +9;
				 l_2 = -23; end
		6123: begin l_1 = -9;
				 l_2 = +23; end
		11978: begin l_1 = -9;
				 l_2 = -23; end
		13014: begin l_1 = +9;
				 l_2 = +24; end
		6111: begin l_1 = +9;
				 l_2 = -24; end
		12502: begin l_1 = -9;
				 l_2 = +24; end
		5599: begin l_1 = -9;
				 l_2 = -24; end
		7159: begin l_1 = +9;
				 l_2 = +25; end
		11966: begin l_1 = +9;
				 l_2 = -25; end
		6647: begin l_1 = -9;
				 l_2 = +25; end
		11454: begin l_1 = -9;
				 l_2 = -25; end
		14062: begin l_1 = +9;
				 l_2 = +26; end
		5063: begin l_1 = +9;
				 l_2 = -26; end
		13550: begin l_1 = -9;
				 l_2 = +26; end
		4551: begin l_1 = -9;
				 l_2 = -26; end
		9255: begin l_1 = +9;
				 l_2 = +27; end
		9870: begin l_1 = +9;
				 l_2 = -27; end
		8743: begin l_1 = -9;
				 l_2 = +27; end
		9358: begin l_1 = -9;
				 l_2 = -27; end
		18254: begin l_1 = +9;
				 l_2 = +28; end
		871: begin l_1 = +9;
				 l_2 = -28; end
		17742: begin l_1 = -9;
				 l_2 = +28; end
		359: begin l_1 = -9;
				 l_2 = -28; end
		17639: begin l_1 = +9;
				 l_2 = +29; end
		1486: begin l_1 = +9;
				 l_2 = -29; end
		17127: begin l_1 = -9;
				 l_2 = +29; end
		974: begin l_1 = -9;
				 l_2 = -29; end
		16409: begin l_1 = +9;
				 l_2 = +30; end
		2716: begin l_1 = +9;
				 l_2 = -30; end
		15897: begin l_1 = -9;
				 l_2 = +30; end
		2204: begin l_1 = -9;
				 l_2 = -30; end
		13949: begin l_1 = +9;
				 l_2 = +31; end
		5176: begin l_1 = +9;
				 l_2 = -31; end
		13437: begin l_1 = -9;
				 l_2 = +31; end
		4664: begin l_1 = -9;
				 l_2 = -31; end
		9029: begin l_1 = +9;
				 l_2 = +32; end
		10096: begin l_1 = +9;
				 l_2 = -32; end
		8517: begin l_1 = -9;
				 l_2 = +32; end
		9584: begin l_1 = -9;
				 l_2 = -32; end
		17802: begin l_1 = +9;
				 l_2 = +33; end
		1323: begin l_1 = +9;
				 l_2 = -33; end
		17290: begin l_1 = -9;
				 l_2 = +33; end
		811: begin l_1 = -9;
				 l_2 = -33; end
		16735: begin l_1 = +9;
				 l_2 = +34; end
		2390: begin l_1 = +9;
				 l_2 = -34; end
		16223: begin l_1 = -9;
				 l_2 = +34; end
		1878: begin l_1 = -9;
				 l_2 = -34; end
		14601: begin l_1 = +9;
				 l_2 = +35; end
		4524: begin l_1 = +9;
				 l_2 = -35; end
		14089: begin l_1 = -9;
				 l_2 = +35; end
		4012: begin l_1 = -9;
				 l_2 = -35; end
		10333: begin l_1 = +9;
				 l_2 = +36; end
		8792: begin l_1 = +9;
				 l_2 = -36; end
		9821: begin l_1 = -9;
				 l_2 = +36; end
		8280: begin l_1 = -9;
				 l_2 = -36; end
		1797: begin l_1 = +9;
				 l_2 = +37; end
		17328: begin l_1 = +9;
				 l_2 = -37; end
		1285: begin l_1 = -9;
				 l_2 = +37; end
		16816: begin l_1 = -9;
				 l_2 = -37; end
		3338: begin l_1 = +9;
				 l_2 = +38; end
		15787: begin l_1 = +9;
				 l_2 = -38; end
		2826: begin l_1 = -9;
				 l_2 = +38; end
		15275: begin l_1 = -9;
				 l_2 = -38; end
		6420: begin l_1 = +9;
				 l_2 = +39; end
		12705: begin l_1 = +9;
				 l_2 = -39; end
		5908: begin l_1 = -9;
				 l_2 = +39; end
		12193: begin l_1 = -9;
				 l_2 = -39; end
		12584: begin l_1 = +9;
				 l_2 = +40; end
		6541: begin l_1 = +9;
				 l_2 = -40; end
		12072: begin l_1 = -9;
				 l_2 = +40; end
		6029: begin l_1 = -9;
				 l_2 = -40; end
		6299: begin l_1 = +9;
				 l_2 = +41; end
		12826: begin l_1 = +9;
				 l_2 = -41; end
		5787: begin l_1 = -9;
				 l_2 = +41; end
		12314: begin l_1 = -9;
				 l_2 = -41; end
		12342: begin l_1 = +9;
				 l_2 = +42; end
		6783: begin l_1 = +9;
				 l_2 = -42; end
		11830: begin l_1 = -9;
				 l_2 = +42; end
		6271: begin l_1 = -9;
				 l_2 = -42; end
		5815: begin l_1 = +9;
				 l_2 = +43; end
		13310: begin l_1 = +9;
				 l_2 = -43; end
		5303: begin l_1 = -9;
				 l_2 = +43; end
		12798: begin l_1 = -9;
				 l_2 = -43; end
		11374: begin l_1 = +9;
				 l_2 = +44; end
		7751: begin l_1 = +9;
				 l_2 = -44; end
		10862: begin l_1 = -9;
				 l_2 = +44; end
		7239: begin l_1 = -9;
				 l_2 = -44; end
		3879: begin l_1 = +9;
				 l_2 = +45; end
		15246: begin l_1 = +9;
				 l_2 = -45; end
		3367: begin l_1 = -9;
				 l_2 = +45; end
		14734: begin l_1 = -9;
				 l_2 = -45; end
		1536: begin l_1 = -10;
				 l_2 = +12; end
		17077: begin l_1 = -10;
				 l_2 = -11; end
		2560: begin l_1 = +10;
				 l_2 = +12; end
		16053: begin l_1 = -10;
				 l_2 = -12; end
		4608: begin l_1 = +10;
				 l_2 = +13; end
		15029: begin l_1 = +10;
				 l_2 = -13; end
		3584: begin l_1 = -10;
				 l_2 = +13; end
		14005: begin l_1 = -10;
				 l_2 = -13; end
		8704: begin l_1 = +10;
				 l_2 = +14; end
		10933: begin l_1 = +10;
				 l_2 = -14; end
		7680: begin l_1 = -10;
				 l_2 = +14; end
		9909: begin l_1 = -10;
				 l_2 = -14; end
		16896: begin l_1 = +10;
				 l_2 = +15; end
		2741: begin l_1 = +10;
				 l_2 = -15; end
		15872: begin l_1 = -10;
				 l_2 = +15; end
		1717: begin l_1 = -10;
				 l_2 = -15; end
		14667: begin l_1 = +10;
				 l_2 = +16; end
		4970: begin l_1 = +10;
				 l_2 = -16; end
		13643: begin l_1 = -10;
				 l_2 = +16; end
		3946: begin l_1 = -10;
				 l_2 = -16; end
		10209: begin l_1 = +10;
				 l_2 = +17; end
		9428: begin l_1 = +10;
				 l_2 = -17; end
		9185: begin l_1 = -10;
				 l_2 = +17; end
		8404: begin l_1 = -10;
				 l_2 = -17; end
		1293: begin l_1 = +10;
				 l_2 = +18; end
		18344: begin l_1 = +10;
				 l_2 = -18; end
		269: begin l_1 = -10;
				 l_2 = +18; end
		17320: begin l_1 = -10;
				 l_2 = -18; end
		2074: begin l_1 = +10;
				 l_2 = +19; end
		17563: begin l_1 = +10;
				 l_2 = -19; end
		1050: begin l_1 = -10;
				 l_2 = +19; end
		16539: begin l_1 = -10;
				 l_2 = -19; end
		3636: begin l_1 = +10;
				 l_2 = +20; end
		16001: begin l_1 = +10;
				 l_2 = -20; end
		2612: begin l_1 = -10;
				 l_2 = +20; end
		14977: begin l_1 = -10;
				 l_2 = -20; end
		6760: begin l_1 = +10;
				 l_2 = +21; end
		12877: begin l_1 = +10;
				 l_2 = -21; end
		5736: begin l_1 = -10;
				 l_2 = +21; end
		11853: begin l_1 = -10;
				 l_2 = -21; end
		13008: begin l_1 = +10;
				 l_2 = +22; end
		6629: begin l_1 = +10;
				 l_2 = -22; end
		11984: begin l_1 = -10;
				 l_2 = +22; end
		5605: begin l_1 = -10;
				 l_2 = -22; end
		6891: begin l_1 = +10;
				 l_2 = +23; end
		12746: begin l_1 = +10;
				 l_2 = -23; end
		5867: begin l_1 = -10;
				 l_2 = +23; end
		11722: begin l_1 = -10;
				 l_2 = -23; end
		13270: begin l_1 = +10;
				 l_2 = +24; end
		6367: begin l_1 = +10;
				 l_2 = -24; end
		12246: begin l_1 = -10;
				 l_2 = +24; end
		5343: begin l_1 = -10;
				 l_2 = -24; end
		7415: begin l_1 = +10;
				 l_2 = +25; end
		12222: begin l_1 = +10;
				 l_2 = -25; end
		6391: begin l_1 = -10;
				 l_2 = +25; end
		11198: begin l_1 = -10;
				 l_2 = -25; end
		14318: begin l_1 = +10;
				 l_2 = +26; end
		5319: begin l_1 = +10;
				 l_2 = -26; end
		13294: begin l_1 = -10;
				 l_2 = +26; end
		4295: begin l_1 = -10;
				 l_2 = -26; end
		9511: begin l_1 = +10;
				 l_2 = +27; end
		10126: begin l_1 = +10;
				 l_2 = -27; end
		8487: begin l_1 = -10;
				 l_2 = +27; end
		9102: begin l_1 = -10;
				 l_2 = -27; end
		18510: begin l_1 = +10;
				 l_2 = +28; end
		1127: begin l_1 = +10;
				 l_2 = -28; end
		17486: begin l_1 = -10;
				 l_2 = +28; end
		103: begin l_1 = -10;
				 l_2 = -28; end
		17895: begin l_1 = +10;
				 l_2 = +29; end
		1742: begin l_1 = +10;
				 l_2 = -29; end
		16871: begin l_1 = -10;
				 l_2 = +29; end
		718: begin l_1 = -10;
				 l_2 = -29; end
		16665: begin l_1 = +10;
				 l_2 = +30; end
		2972: begin l_1 = +10;
				 l_2 = -30; end
		15641: begin l_1 = -10;
				 l_2 = +30; end
		1948: begin l_1 = -10;
				 l_2 = -30; end
		14205: begin l_1 = +10;
				 l_2 = +31; end
		5432: begin l_1 = +10;
				 l_2 = -31; end
		13181: begin l_1 = -10;
				 l_2 = +31; end
		4408: begin l_1 = -10;
				 l_2 = -31; end
		9285: begin l_1 = +10;
				 l_2 = +32; end
		10352: begin l_1 = +10;
				 l_2 = -32; end
		8261: begin l_1 = -10;
				 l_2 = +32; end
		9328: begin l_1 = -10;
				 l_2 = -32; end
		18058: begin l_1 = +10;
				 l_2 = +33; end
		1579: begin l_1 = +10;
				 l_2 = -33; end
		17034: begin l_1 = -10;
				 l_2 = +33; end
		555: begin l_1 = -10;
				 l_2 = -33; end
		16991: begin l_1 = +10;
				 l_2 = +34; end
		2646: begin l_1 = +10;
				 l_2 = -34; end
		15967: begin l_1 = -10;
				 l_2 = +34; end
		1622: begin l_1 = -10;
				 l_2 = -34; end
		14857: begin l_1 = +10;
				 l_2 = +35; end
		4780: begin l_1 = +10;
				 l_2 = -35; end
		13833: begin l_1 = -10;
				 l_2 = +35; end
		3756: begin l_1 = -10;
				 l_2 = -35; end
		10589: begin l_1 = +10;
				 l_2 = +36; end
		9048: begin l_1 = +10;
				 l_2 = -36; end
		9565: begin l_1 = -10;
				 l_2 = +36; end
		8024: begin l_1 = -10;
				 l_2 = -36; end
		2053: begin l_1 = +10;
				 l_2 = +37; end
		17584: begin l_1 = +10;
				 l_2 = -37; end
		1029: begin l_1 = -10;
				 l_2 = +37; end
		16560: begin l_1 = -10;
				 l_2 = -37; end
		3594: begin l_1 = +10;
				 l_2 = +38; end
		16043: begin l_1 = +10;
				 l_2 = -38; end
		2570: begin l_1 = -10;
				 l_2 = +38; end
		15019: begin l_1 = -10;
				 l_2 = -38; end
		6676: begin l_1 = +10;
				 l_2 = +39; end
		12961: begin l_1 = +10;
				 l_2 = -39; end
		5652: begin l_1 = -10;
				 l_2 = +39; end
		11937: begin l_1 = -10;
				 l_2 = -39; end
		12840: begin l_1 = +10;
				 l_2 = +40; end
		6797: begin l_1 = +10;
				 l_2 = -40; end
		11816: begin l_1 = -10;
				 l_2 = +40; end
		5773: begin l_1 = -10;
				 l_2 = -40; end
		6555: begin l_1 = +10;
				 l_2 = +41; end
		13082: begin l_1 = +10;
				 l_2 = -41; end
		5531: begin l_1 = -10;
				 l_2 = +41; end
		12058: begin l_1 = -10;
				 l_2 = -41; end
		12598: begin l_1 = +10;
				 l_2 = +42; end
		7039: begin l_1 = +10;
				 l_2 = -42; end
		11574: begin l_1 = -10;
				 l_2 = +42; end
		6015: begin l_1 = -10;
				 l_2 = -42; end
		6071: begin l_1 = +10;
				 l_2 = +43; end
		13566: begin l_1 = +10;
				 l_2 = -43; end
		5047: begin l_1 = -10;
				 l_2 = +43; end
		12542: begin l_1 = -10;
				 l_2 = -43; end
		11630: begin l_1 = +10;
				 l_2 = +44; end
		8007: begin l_1 = +10;
				 l_2 = -44; end
		10606: begin l_1 = -10;
				 l_2 = +44; end
		6983: begin l_1 = -10;
				 l_2 = -44; end
		4135: begin l_1 = +10;
				 l_2 = +45; end
		15502: begin l_1 = +10;
				 l_2 = -45; end
		3111: begin l_1 = -10;
				 l_2 = +45; end
		14478: begin l_1 = -10;
				 l_2 = -45; end
		3072: begin l_1 = -11;
				 l_2 = +13; end
		15541: begin l_1 = -11;
				 l_2 = -12; end
		5120: begin l_1 = +11;
				 l_2 = +13; end
		13493: begin l_1 = -11;
				 l_2 = -13; end
		9216: begin l_1 = +11;
				 l_2 = +14; end
		11445: begin l_1 = +11;
				 l_2 = -14; end
		7168: begin l_1 = -11;
				 l_2 = +14; end
		9397: begin l_1 = -11;
				 l_2 = -14; end
		17408: begin l_1 = +11;
				 l_2 = +15; end
		3253: begin l_1 = +11;
				 l_2 = -15; end
		15360: begin l_1 = -11;
				 l_2 = +15; end
		1205: begin l_1 = -11;
				 l_2 = -15; end
		15179: begin l_1 = +11;
				 l_2 = +16; end
		5482: begin l_1 = +11;
				 l_2 = -16; end
		13131: begin l_1 = -11;
				 l_2 = +16; end
		3434: begin l_1 = -11;
				 l_2 = -16; end
		10721: begin l_1 = +11;
				 l_2 = +17; end
		9940: begin l_1 = +11;
				 l_2 = -17; end
		8673: begin l_1 = -11;
				 l_2 = +17; end
		7892: begin l_1 = -11;
				 l_2 = -17; end
		1805: begin l_1 = +11;
				 l_2 = +18; end
		243: begin l_1 = +11;
				 l_2 = -18; end
		18370: begin l_1 = -11;
				 l_2 = +18; end
		16808: begin l_1 = -11;
				 l_2 = -18; end
		2586: begin l_1 = +11;
				 l_2 = +19; end
		18075: begin l_1 = +11;
				 l_2 = -19; end
		538: begin l_1 = -11;
				 l_2 = +19; end
		16027: begin l_1 = -11;
				 l_2 = -19; end
		4148: begin l_1 = +11;
				 l_2 = +20; end
		16513: begin l_1 = +11;
				 l_2 = -20; end
		2100: begin l_1 = -11;
				 l_2 = +20; end
		14465: begin l_1 = -11;
				 l_2 = -20; end
		7272: begin l_1 = +11;
				 l_2 = +21; end
		13389: begin l_1 = +11;
				 l_2 = -21; end
		5224: begin l_1 = -11;
				 l_2 = +21; end
		11341: begin l_1 = -11;
				 l_2 = -21; end
		13520: begin l_1 = +11;
				 l_2 = +22; end
		7141: begin l_1 = +11;
				 l_2 = -22; end
		11472: begin l_1 = -11;
				 l_2 = +22; end
		5093: begin l_1 = -11;
				 l_2 = -22; end
		7403: begin l_1 = +11;
				 l_2 = +23; end
		13258: begin l_1 = +11;
				 l_2 = -23; end
		5355: begin l_1 = -11;
				 l_2 = +23; end
		11210: begin l_1 = -11;
				 l_2 = -23; end
		13782: begin l_1 = +11;
				 l_2 = +24; end
		6879: begin l_1 = +11;
				 l_2 = -24; end
		11734: begin l_1 = -11;
				 l_2 = +24; end
		4831: begin l_1 = -11;
				 l_2 = -24; end
		7927: begin l_1 = +11;
				 l_2 = +25; end
		12734: begin l_1 = +11;
				 l_2 = -25; end
		5879: begin l_1 = -11;
				 l_2 = +25; end
		10686: begin l_1 = -11;
				 l_2 = -25; end
		14830: begin l_1 = +11;
				 l_2 = +26; end
		5831: begin l_1 = +11;
				 l_2 = -26; end
		12782: begin l_1 = -11;
				 l_2 = +26; end
		3783: begin l_1 = -11;
				 l_2 = -26; end
		10023: begin l_1 = +11;
				 l_2 = +27; end
		10638: begin l_1 = +11;
				 l_2 = -27; end
		7975: begin l_1 = -11;
				 l_2 = +27; end
		8590: begin l_1 = -11;
				 l_2 = -27; end
		409: begin l_1 = +11;
				 l_2 = +28; end
		1639: begin l_1 = +11;
				 l_2 = -28; end
		16974: begin l_1 = -11;
				 l_2 = +28; end
		18204: begin l_1 = -11;
				 l_2 = -28; end
		18407: begin l_1 = +11;
				 l_2 = +29; end
		2254: begin l_1 = +11;
				 l_2 = -29; end
		16359: begin l_1 = -11;
				 l_2 = +29; end
		206: begin l_1 = -11;
				 l_2 = -29; end
		17177: begin l_1 = +11;
				 l_2 = +30; end
		3484: begin l_1 = +11;
				 l_2 = -30; end
		15129: begin l_1 = -11;
				 l_2 = +30; end
		1436: begin l_1 = -11;
				 l_2 = -30; end
		14717: begin l_1 = +11;
				 l_2 = +31; end
		5944: begin l_1 = +11;
				 l_2 = -31; end
		12669: begin l_1 = -11;
				 l_2 = +31; end
		3896: begin l_1 = -11;
				 l_2 = -31; end
		9797: begin l_1 = +11;
				 l_2 = +32; end
		10864: begin l_1 = +11;
				 l_2 = -32; end
		7749: begin l_1 = -11;
				 l_2 = +32; end
		8816: begin l_1 = -11;
				 l_2 = -32; end
		18570: begin l_1 = +11;
				 l_2 = +33; end
		2091: begin l_1 = +11;
				 l_2 = -33; end
		16522: begin l_1 = -11;
				 l_2 = +33; end
		43: begin l_1 = -11;
				 l_2 = -33; end
		17503: begin l_1 = +11;
				 l_2 = +34; end
		3158: begin l_1 = +11;
				 l_2 = -34; end
		15455: begin l_1 = -11;
				 l_2 = +34; end
		1110: begin l_1 = -11;
				 l_2 = -34; end
		15369: begin l_1 = +11;
				 l_2 = +35; end
		5292: begin l_1 = +11;
				 l_2 = -35; end
		13321: begin l_1 = -11;
				 l_2 = +35; end
		3244: begin l_1 = -11;
				 l_2 = -35; end
		11101: begin l_1 = +11;
				 l_2 = +36; end
		9560: begin l_1 = +11;
				 l_2 = -36; end
		9053: begin l_1 = -11;
				 l_2 = +36; end
		7512: begin l_1 = -11;
				 l_2 = -36; end
		2565: begin l_1 = +11;
				 l_2 = +37; end
		18096: begin l_1 = +11;
				 l_2 = -37; end
		517: begin l_1 = -11;
				 l_2 = +37; end
		16048: begin l_1 = -11;
				 l_2 = -37; end
		4106: begin l_1 = +11;
				 l_2 = +38; end
		16555: begin l_1 = +11;
				 l_2 = -38; end
		2058: begin l_1 = -11;
				 l_2 = +38; end
		14507: begin l_1 = -11;
				 l_2 = -38; end
		7188: begin l_1 = +11;
				 l_2 = +39; end
		13473: begin l_1 = +11;
				 l_2 = -39; end
		5140: begin l_1 = -11;
				 l_2 = +39; end
		11425: begin l_1 = -11;
				 l_2 = -39; end
		13352: begin l_1 = +11;
				 l_2 = +40; end
		7309: begin l_1 = +11;
				 l_2 = -40; end
		11304: begin l_1 = -11;
				 l_2 = +40; end
		5261: begin l_1 = -11;
				 l_2 = -40; end
		7067: begin l_1 = +11;
				 l_2 = +41; end
		13594: begin l_1 = +11;
				 l_2 = -41; end
		5019: begin l_1 = -11;
				 l_2 = +41; end
		11546: begin l_1 = -11;
				 l_2 = -41; end
		13110: begin l_1 = +11;
				 l_2 = +42; end
		7551: begin l_1 = +11;
				 l_2 = -42; end
		11062: begin l_1 = -11;
				 l_2 = +42; end
		5503: begin l_1 = -11;
				 l_2 = -42; end
		6583: begin l_1 = +11;
				 l_2 = +43; end
		14078: begin l_1 = +11;
				 l_2 = -43; end
		4535: begin l_1 = -11;
				 l_2 = +43; end
		12030: begin l_1 = -11;
				 l_2 = -43; end
		12142: begin l_1 = +11;
				 l_2 = +44; end
		8519: begin l_1 = +11;
				 l_2 = -44; end
		10094: begin l_1 = -11;
				 l_2 = +44; end
		6471: begin l_1 = -11;
				 l_2 = -44; end
		4647: begin l_1 = +11;
				 l_2 = +45; end
		16014: begin l_1 = +11;
				 l_2 = -45; end
		2599: begin l_1 = -11;
				 l_2 = +45; end
		13966: begin l_1 = -11;
				 l_2 = -45; end
		6144: begin l_1 = -12;
				 l_2 = +14; end
		12469: begin l_1 = -12;
				 l_2 = -13; end
		10240: begin l_1 = +12;
				 l_2 = +14; end
		8373: begin l_1 = -12;
				 l_2 = -14; end
		18432: begin l_1 = +12;
				 l_2 = +15; end
		4277: begin l_1 = +12;
				 l_2 = -15; end
		14336: begin l_1 = -12;
				 l_2 = +15; end
		181: begin l_1 = -12;
				 l_2 = -15; end
		16203: begin l_1 = +12;
				 l_2 = +16; end
		6506: begin l_1 = +12;
				 l_2 = -16; end
		12107: begin l_1 = -12;
				 l_2 = +16; end
		2410: begin l_1 = -12;
				 l_2 = -16; end
		11745: begin l_1 = +12;
				 l_2 = +17; end
		10964: begin l_1 = +12;
				 l_2 = -17; end
		7649: begin l_1 = -12;
				 l_2 = +17; end
		6868: begin l_1 = -12;
				 l_2 = -17; end
		2829: begin l_1 = +12;
				 l_2 = +18; end
		1267: begin l_1 = +12;
				 l_2 = -18; end
		17346: begin l_1 = -12;
				 l_2 = +18; end
		15784: begin l_1 = -12;
				 l_2 = -18; end
		3610: begin l_1 = +12;
				 l_2 = +19; end
		486: begin l_1 = +12;
				 l_2 = -19; end
		18127: begin l_1 = -12;
				 l_2 = +19; end
		15003: begin l_1 = -12;
				 l_2 = -19; end
		5172: begin l_1 = +12;
				 l_2 = +20; end
		17537: begin l_1 = +12;
				 l_2 = -20; end
		1076: begin l_1 = -12;
				 l_2 = +20; end
		13441: begin l_1 = -12;
				 l_2 = -20; end
		8296: begin l_1 = +12;
				 l_2 = +21; end
		14413: begin l_1 = +12;
				 l_2 = -21; end
		4200: begin l_1 = -12;
				 l_2 = +21; end
		10317: begin l_1 = -12;
				 l_2 = -21; end
		14544: begin l_1 = +12;
				 l_2 = +22; end
		8165: begin l_1 = +12;
				 l_2 = -22; end
		10448: begin l_1 = -12;
				 l_2 = +22; end
		4069: begin l_1 = -12;
				 l_2 = -22; end
		8427: begin l_1 = +12;
				 l_2 = +23; end
		14282: begin l_1 = +12;
				 l_2 = -23; end
		4331: begin l_1 = -12;
				 l_2 = +23; end
		10186: begin l_1 = -12;
				 l_2 = -23; end
		14806: begin l_1 = +12;
				 l_2 = +24; end
		7903: begin l_1 = +12;
				 l_2 = -24; end
		10710: begin l_1 = -12;
				 l_2 = +24; end
		3807: begin l_1 = -12;
				 l_2 = -24; end
		8951: begin l_1 = +12;
				 l_2 = +25; end
		13758: begin l_1 = +12;
				 l_2 = -25; end
		4855: begin l_1 = -12;
				 l_2 = +25; end
		9662: begin l_1 = -12;
				 l_2 = -25; end
		15854: begin l_1 = +12;
				 l_2 = +26; end
		6855: begin l_1 = +12;
				 l_2 = -26; end
		11758: begin l_1 = -12;
				 l_2 = +26; end
		2759: begin l_1 = -12;
				 l_2 = -26; end
		11047: begin l_1 = +12;
				 l_2 = +27; end
		11662: begin l_1 = +12;
				 l_2 = -27; end
		6951: begin l_1 = -12;
				 l_2 = +27; end
		7566: begin l_1 = -12;
				 l_2 = -27; end
		1433: begin l_1 = +12;
				 l_2 = +28; end
		2663: begin l_1 = +12;
				 l_2 = -28; end
		15950: begin l_1 = -12;
				 l_2 = +28; end
		17180: begin l_1 = -12;
				 l_2 = -28; end
		818: begin l_1 = +12;
				 l_2 = +29; end
		3278: begin l_1 = +12;
				 l_2 = -29; end
		15335: begin l_1 = -12;
				 l_2 = +29; end
		17795: begin l_1 = -12;
				 l_2 = -29; end
		18201: begin l_1 = +12;
				 l_2 = +30; end
		4508: begin l_1 = +12;
				 l_2 = -30; end
		14105: begin l_1 = -12;
				 l_2 = +30; end
		412: begin l_1 = -12;
				 l_2 = -30; end
		15741: begin l_1 = +12;
				 l_2 = +31; end
		6968: begin l_1 = +12;
				 l_2 = -31; end
		11645: begin l_1 = -12;
				 l_2 = +31; end
		2872: begin l_1 = -12;
				 l_2 = -31; end
		10821: begin l_1 = +12;
				 l_2 = +32; end
		11888: begin l_1 = +12;
				 l_2 = -32; end
		6725: begin l_1 = -12;
				 l_2 = +32; end
		7792: begin l_1 = -12;
				 l_2 = -32; end
		981: begin l_1 = +12;
				 l_2 = +33; end
		3115: begin l_1 = +12;
				 l_2 = -33; end
		15498: begin l_1 = -12;
				 l_2 = +33; end
		17632: begin l_1 = -12;
				 l_2 = -33; end
		18527: begin l_1 = +12;
				 l_2 = +34; end
		4182: begin l_1 = +12;
				 l_2 = -34; end
		14431: begin l_1 = -12;
				 l_2 = +34; end
		86: begin l_1 = -12;
				 l_2 = -34; end
		16393: begin l_1 = +12;
				 l_2 = +35; end
		6316: begin l_1 = +12;
				 l_2 = -35; end
		12297: begin l_1 = -12;
				 l_2 = +35; end
		2220: begin l_1 = -12;
				 l_2 = -35; end
		12125: begin l_1 = +12;
				 l_2 = +36; end
		10584: begin l_1 = +12;
				 l_2 = -36; end
		8029: begin l_1 = -12;
				 l_2 = +36; end
		6488: begin l_1 = -12;
				 l_2 = -36; end
		3589: begin l_1 = +12;
				 l_2 = +37; end
		507: begin l_1 = +12;
				 l_2 = -37; end
		18106: begin l_1 = -12;
				 l_2 = +37; end
		15024: begin l_1 = -12;
				 l_2 = -37; end
		5130: begin l_1 = +12;
				 l_2 = +38; end
		17579: begin l_1 = +12;
				 l_2 = -38; end
		1034: begin l_1 = -12;
				 l_2 = +38; end
		13483: begin l_1 = -12;
				 l_2 = -38; end
		8212: begin l_1 = +12;
				 l_2 = +39; end
		14497: begin l_1 = +12;
				 l_2 = -39; end
		4116: begin l_1 = -12;
				 l_2 = +39; end
		10401: begin l_1 = -12;
				 l_2 = -39; end
		14376: begin l_1 = +12;
				 l_2 = +40; end
		8333: begin l_1 = +12;
				 l_2 = -40; end
		10280: begin l_1 = -12;
				 l_2 = +40; end
		4237: begin l_1 = -12;
				 l_2 = -40; end
		8091: begin l_1 = +12;
				 l_2 = +41; end
		14618: begin l_1 = +12;
				 l_2 = -41; end
		3995: begin l_1 = -12;
				 l_2 = +41; end
		10522: begin l_1 = -12;
				 l_2 = -41; end
		14134: begin l_1 = +12;
				 l_2 = +42; end
		8575: begin l_1 = +12;
				 l_2 = -42; end
		10038: begin l_1 = -12;
				 l_2 = +42; end
		4479: begin l_1 = -12;
				 l_2 = -42; end
		7607: begin l_1 = +12;
				 l_2 = +43; end
		15102: begin l_1 = +12;
				 l_2 = -43; end
		3511: begin l_1 = -12;
				 l_2 = +43; end
		11006: begin l_1 = -12;
				 l_2 = -43; end
		13166: begin l_1 = +12;
				 l_2 = +44; end
		9543: begin l_1 = +12;
				 l_2 = -44; end
		9070: begin l_1 = -12;
				 l_2 = +44; end
		5447: begin l_1 = -12;
				 l_2 = -44; end
		5671: begin l_1 = +12;
				 l_2 = +45; end
		17038: begin l_1 = +12;
				 l_2 = -45; end
		1575: begin l_1 = -12;
				 l_2 = +45; end
		12942: begin l_1 = -12;
				 l_2 = -45; end
		12288: begin l_1 = -13;
				 l_2 = +15; end
		6325: begin l_1 = -13;
				 l_2 = -14; end
		1867: begin l_1 = +13;
				 l_2 = +15; end
		16746: begin l_1 = -13;
				 l_2 = -15; end
		18251: begin l_1 = +13;
				 l_2 = +16; end
		8554: begin l_1 = +13;
				 l_2 = -16; end
		10059: begin l_1 = -13;
				 l_2 = +16; end
		362: begin l_1 = -13;
				 l_2 = -16; end
		13793: begin l_1 = +13;
				 l_2 = +17; end
		13012: begin l_1 = +13;
				 l_2 = -17; end
		5601: begin l_1 = -13;
				 l_2 = +17; end
		4820: begin l_1 = -13;
				 l_2 = -17; end
		4877: begin l_1 = +13;
				 l_2 = +18; end
		3315: begin l_1 = +13;
				 l_2 = -18; end
		15298: begin l_1 = -13;
				 l_2 = +18; end
		13736: begin l_1 = -13;
				 l_2 = -18; end
		5658: begin l_1 = +13;
				 l_2 = +19; end
		2534: begin l_1 = +13;
				 l_2 = -19; end
		16079: begin l_1 = -13;
				 l_2 = +19; end
		12955: begin l_1 = -13;
				 l_2 = -19; end
		7220: begin l_1 = +13;
				 l_2 = +20; end
		972: begin l_1 = +13;
				 l_2 = -20; end
		17641: begin l_1 = -13;
				 l_2 = +20; end
		11393: begin l_1 = -13;
				 l_2 = -20; end
		10344: begin l_1 = +13;
				 l_2 = +21; end
		16461: begin l_1 = +13;
				 l_2 = -21; end
		2152: begin l_1 = -13;
				 l_2 = +21; end
		8269: begin l_1 = -13;
				 l_2 = -21; end
		16592: begin l_1 = +13;
				 l_2 = +22; end
		10213: begin l_1 = +13;
				 l_2 = -22; end
		8400: begin l_1 = -13;
				 l_2 = +22; end
		2021: begin l_1 = -13;
				 l_2 = -22; end
		10475: begin l_1 = +13;
				 l_2 = +23; end
		16330: begin l_1 = +13;
				 l_2 = -23; end
		2283: begin l_1 = -13;
				 l_2 = +23; end
		8138: begin l_1 = -13;
				 l_2 = -23; end
		16854: begin l_1 = +13;
				 l_2 = +24; end
		9951: begin l_1 = +13;
				 l_2 = -24; end
		8662: begin l_1 = -13;
				 l_2 = +24; end
		1759: begin l_1 = -13;
				 l_2 = -24; end
		10999: begin l_1 = +13;
				 l_2 = +25; end
		15806: begin l_1 = +13;
				 l_2 = -25; end
		2807: begin l_1 = -13;
				 l_2 = +25; end
		7614: begin l_1 = -13;
				 l_2 = -25; end
		17902: begin l_1 = +13;
				 l_2 = +26; end
		8903: begin l_1 = +13;
				 l_2 = -26; end
		9710: begin l_1 = -13;
				 l_2 = +26; end
		711: begin l_1 = -13;
				 l_2 = -26; end
		13095: begin l_1 = +13;
				 l_2 = +27; end
		13710: begin l_1 = +13;
				 l_2 = -27; end
		4903: begin l_1 = -13;
				 l_2 = +27; end
		5518: begin l_1 = -13;
				 l_2 = -27; end
		3481: begin l_1 = +13;
				 l_2 = +28; end
		4711: begin l_1 = +13;
				 l_2 = -28; end
		13902: begin l_1 = -13;
				 l_2 = +28; end
		15132: begin l_1 = -13;
				 l_2 = -28; end
		2866: begin l_1 = +13;
				 l_2 = +29; end
		5326: begin l_1 = +13;
				 l_2 = -29; end
		13287: begin l_1 = -13;
				 l_2 = +29; end
		15747: begin l_1 = -13;
				 l_2 = -29; end
		1636: begin l_1 = +13;
				 l_2 = +30; end
		6556: begin l_1 = +13;
				 l_2 = -30; end
		12057: begin l_1 = -13;
				 l_2 = +30; end
		16977: begin l_1 = -13;
				 l_2 = -30; end
		17789: begin l_1 = +13;
				 l_2 = +31; end
		9016: begin l_1 = +13;
				 l_2 = -31; end
		9597: begin l_1 = -13;
				 l_2 = +31; end
		824: begin l_1 = -13;
				 l_2 = -31; end
		12869: begin l_1 = +13;
				 l_2 = +32; end
		13936: begin l_1 = +13;
				 l_2 = -32; end
		4677: begin l_1 = -13;
				 l_2 = +32; end
		5744: begin l_1 = -13;
				 l_2 = -32; end
		3029: begin l_1 = +13;
				 l_2 = +33; end
		5163: begin l_1 = +13;
				 l_2 = -33; end
		13450: begin l_1 = -13;
				 l_2 = +33; end
		15584: begin l_1 = -13;
				 l_2 = -33; end
		1962: begin l_1 = +13;
				 l_2 = +34; end
		6230: begin l_1 = +13;
				 l_2 = -34; end
		12383: begin l_1 = -13;
				 l_2 = +34; end
		16651: begin l_1 = -13;
				 l_2 = -34; end
		18441: begin l_1 = +13;
				 l_2 = +35; end
		8364: begin l_1 = +13;
				 l_2 = -35; end
		10249: begin l_1 = -13;
				 l_2 = +35; end
		172: begin l_1 = -13;
				 l_2 = -35; end
		14173: begin l_1 = +13;
				 l_2 = +36; end
		12632: begin l_1 = +13;
				 l_2 = -36; end
		5981: begin l_1 = -13;
				 l_2 = +36; end
		4440: begin l_1 = -13;
				 l_2 = -36; end
		5637: begin l_1 = +13;
				 l_2 = +37; end
		2555: begin l_1 = +13;
				 l_2 = -37; end
		16058: begin l_1 = -13;
				 l_2 = +37; end
		12976: begin l_1 = -13;
				 l_2 = -37; end
		7178: begin l_1 = +13;
				 l_2 = +38; end
		1014: begin l_1 = +13;
				 l_2 = -38; end
		17599: begin l_1 = -13;
				 l_2 = +38; end
		11435: begin l_1 = -13;
				 l_2 = -38; end
		10260: begin l_1 = +13;
				 l_2 = +39; end
		16545: begin l_1 = +13;
				 l_2 = -39; end
		2068: begin l_1 = -13;
				 l_2 = +39; end
		8353: begin l_1 = -13;
				 l_2 = -39; end
		16424: begin l_1 = +13;
				 l_2 = +40; end
		10381: begin l_1 = +13;
				 l_2 = -40; end
		8232: begin l_1 = -13;
				 l_2 = +40; end
		2189: begin l_1 = -13;
				 l_2 = -40; end
		10139: begin l_1 = +13;
				 l_2 = +41; end
		16666: begin l_1 = +13;
				 l_2 = -41; end
		1947: begin l_1 = -13;
				 l_2 = +41; end
		8474: begin l_1 = -13;
				 l_2 = -41; end
		16182: begin l_1 = +13;
				 l_2 = +42; end
		10623: begin l_1 = +13;
				 l_2 = -42; end
		7990: begin l_1 = -13;
				 l_2 = +42; end
		2431: begin l_1 = -13;
				 l_2 = -42; end
		9655: begin l_1 = +13;
				 l_2 = +43; end
		17150: begin l_1 = +13;
				 l_2 = -43; end
		1463: begin l_1 = -13;
				 l_2 = +43; end
		8958: begin l_1 = -13;
				 l_2 = -43; end
		15214: begin l_1 = +13;
				 l_2 = +44; end
		11591: begin l_1 = +13;
				 l_2 = -44; end
		7022: begin l_1 = -13;
				 l_2 = +44; end
		3399: begin l_1 = -13;
				 l_2 = -44; end
		7719: begin l_1 = +13;
				 l_2 = +45; end
		473: begin l_1 = +13;
				 l_2 = -45; end
		18140: begin l_1 = -13;
				 l_2 = +45; end
		10894: begin l_1 = -13;
				 l_2 = -45; end
		5963: begin l_1 = -14;
				 l_2 = +16; end
		12650: begin l_1 = -14;
				 l_2 = -15; end
		3734: begin l_1 = +14;
				 l_2 = +16; end
		14879: begin l_1 = -14;
				 l_2 = -16; end
		17889: begin l_1 = +14;
				 l_2 = +17; end
		17108: begin l_1 = +14;
				 l_2 = -17; end
		1505: begin l_1 = -14;
				 l_2 = +17; end
		724: begin l_1 = -14;
				 l_2 = -17; end
		8973: begin l_1 = +14;
				 l_2 = +18; end
		7411: begin l_1 = +14;
				 l_2 = -18; end
		11202: begin l_1 = -14;
				 l_2 = +18; end
		9640: begin l_1 = -14;
				 l_2 = -18; end
		9754: begin l_1 = +14;
				 l_2 = +19; end
		6630: begin l_1 = +14;
				 l_2 = -19; end
		11983: begin l_1 = -14;
				 l_2 = +19; end
		8859: begin l_1 = -14;
				 l_2 = -19; end
		11316: begin l_1 = +14;
				 l_2 = +20; end
		5068: begin l_1 = +14;
				 l_2 = -20; end
		13545: begin l_1 = -14;
				 l_2 = +20; end
		7297: begin l_1 = -14;
				 l_2 = -20; end
		14440: begin l_1 = +14;
				 l_2 = +21; end
		1944: begin l_1 = +14;
				 l_2 = -21; end
		16669: begin l_1 = -14;
				 l_2 = +21; end
		4173: begin l_1 = -14;
				 l_2 = -21; end
		2075: begin l_1 = +14;
				 l_2 = +22; end
		14309: begin l_1 = +14;
				 l_2 = -22; end
		4304: begin l_1 = -14;
				 l_2 = +22; end
		16538: begin l_1 = -14;
				 l_2 = -22; end
		14571: begin l_1 = +14;
				 l_2 = +23; end
		1813: begin l_1 = +14;
				 l_2 = -23; end
		16800: begin l_1 = -14;
				 l_2 = +23; end
		4042: begin l_1 = -14;
				 l_2 = -23; end
		2337: begin l_1 = +14;
				 l_2 = +24; end
		14047: begin l_1 = +14;
				 l_2 = -24; end
		4566: begin l_1 = -14;
				 l_2 = +24; end
		16276: begin l_1 = -14;
				 l_2 = -24; end
		15095: begin l_1 = +14;
				 l_2 = +25; end
		1289: begin l_1 = +14;
				 l_2 = -25; end
		17324: begin l_1 = -14;
				 l_2 = +25; end
		3518: begin l_1 = -14;
				 l_2 = -25; end
		3385: begin l_1 = +14;
				 l_2 = +26; end
		12999: begin l_1 = +14;
				 l_2 = -26; end
		5614: begin l_1 = -14;
				 l_2 = +26; end
		15228: begin l_1 = -14;
				 l_2 = -26; end
		17191: begin l_1 = +14;
				 l_2 = +27; end
		17806: begin l_1 = +14;
				 l_2 = -27; end
		807: begin l_1 = -14;
				 l_2 = +27; end
		1422: begin l_1 = -14;
				 l_2 = -27; end
		7577: begin l_1 = +14;
				 l_2 = +28; end
		8807: begin l_1 = +14;
				 l_2 = -28; end
		9806: begin l_1 = -14;
				 l_2 = +28; end
		11036: begin l_1 = -14;
				 l_2 = -28; end
		6962: begin l_1 = +14;
				 l_2 = +29; end
		9422: begin l_1 = +14;
				 l_2 = -29; end
		9191: begin l_1 = -14;
				 l_2 = +29; end
		11651: begin l_1 = -14;
				 l_2 = -29; end
		5732: begin l_1 = +14;
				 l_2 = +30; end
		10652: begin l_1 = +14;
				 l_2 = -30; end
		7961: begin l_1 = -14;
				 l_2 = +30; end
		12881: begin l_1 = -14;
				 l_2 = -30; end
		3272: begin l_1 = +14;
				 l_2 = +31; end
		13112: begin l_1 = +14;
				 l_2 = -31; end
		5501: begin l_1 = -14;
				 l_2 = +31; end
		15341: begin l_1 = -14;
				 l_2 = -31; end
		16965: begin l_1 = +14;
				 l_2 = +32; end
		18032: begin l_1 = +14;
				 l_2 = -32; end
		581: begin l_1 = -14;
				 l_2 = +32; end
		1648: begin l_1 = -14;
				 l_2 = -32; end
		7125: begin l_1 = +14;
				 l_2 = +33; end
		9259: begin l_1 = +14;
				 l_2 = -33; end
		9354: begin l_1 = -14;
				 l_2 = +33; end
		11488: begin l_1 = -14;
				 l_2 = -33; end
		6058: begin l_1 = +14;
				 l_2 = +34; end
		10326: begin l_1 = +14;
				 l_2 = -34; end
		8287: begin l_1 = -14;
				 l_2 = +34; end
		12555: begin l_1 = -14;
				 l_2 = -34; end
		3924: begin l_1 = +14;
				 l_2 = +35; end
		12460: begin l_1 = +14;
				 l_2 = -35; end
		6153: begin l_1 = -14;
				 l_2 = +35; end
		14689: begin l_1 = -14;
				 l_2 = -35; end
		18269: begin l_1 = +14;
				 l_2 = +36; end
		16728: begin l_1 = +14;
				 l_2 = -36; end
		1885: begin l_1 = -14;
				 l_2 = +36; end
		344: begin l_1 = -14;
				 l_2 = -36; end
		9733: begin l_1 = +14;
				 l_2 = +37; end
		6651: begin l_1 = +14;
				 l_2 = -37; end
		11962: begin l_1 = -14;
				 l_2 = +37; end
		8880: begin l_1 = -14;
				 l_2 = -37; end
		11274: begin l_1 = +14;
				 l_2 = +38; end
		5110: begin l_1 = +14;
				 l_2 = -38; end
		13503: begin l_1 = -14;
				 l_2 = +38; end
		7339: begin l_1 = -14;
				 l_2 = -38; end
		14356: begin l_1 = +14;
				 l_2 = +39; end
		2028: begin l_1 = +14;
				 l_2 = -39; end
		16585: begin l_1 = -14;
				 l_2 = +39; end
		4257: begin l_1 = -14;
				 l_2 = -39; end
		1907: begin l_1 = +14;
				 l_2 = +40; end
		14477: begin l_1 = +14;
				 l_2 = -40; end
		4136: begin l_1 = -14;
				 l_2 = +40; end
		16706: begin l_1 = -14;
				 l_2 = -40; end
		14235: begin l_1 = +14;
				 l_2 = +41; end
		2149: begin l_1 = +14;
				 l_2 = -41; end
		16464: begin l_1 = -14;
				 l_2 = +41; end
		4378: begin l_1 = -14;
				 l_2 = -41; end
		1665: begin l_1 = +14;
				 l_2 = +42; end
		14719: begin l_1 = +14;
				 l_2 = -42; end
		3894: begin l_1 = -14;
				 l_2 = +42; end
		16948: begin l_1 = -14;
				 l_2 = -42; end
		13751: begin l_1 = +14;
				 l_2 = +43; end
		2633: begin l_1 = +14;
				 l_2 = -43; end
		15980: begin l_1 = -14;
				 l_2 = +43; end
		4862: begin l_1 = -14;
				 l_2 = -43; end
		697: begin l_1 = +14;
				 l_2 = +44; end
		15687: begin l_1 = +14;
				 l_2 = -44; end
		2926: begin l_1 = -14;
				 l_2 = +44; end
		17916: begin l_1 = -14;
				 l_2 = -44; end
		11815: begin l_1 = +14;
				 l_2 = +45; end
		4569: begin l_1 = +14;
				 l_2 = -45; end
		14044: begin l_1 = -14;
				 l_2 = +45; end
		6798: begin l_1 = -14;
				 l_2 = -45; end
		11926: begin l_1 = -15;
				 l_2 = +17; end
		6687: begin l_1 = -15;
				 l_2 = -16; end
		7468: begin l_1 = +15;
				 l_2 = +17; end
		11145: begin l_1 = -15;
				 l_2 = -17; end
		17165: begin l_1 = +15;
				 l_2 = +18; end
		15603: begin l_1 = +15;
				 l_2 = -18; end
		3010: begin l_1 = -15;
				 l_2 = +18; end
		1448: begin l_1 = -15;
				 l_2 = -18; end
		17946: begin l_1 = +15;
				 l_2 = +19; end
		14822: begin l_1 = +15;
				 l_2 = -19; end
		3791: begin l_1 = -15;
				 l_2 = +19; end
		667: begin l_1 = -15;
				 l_2 = -19; end
		895: begin l_1 = +15;
				 l_2 = +20; end
		13260: begin l_1 = +15;
				 l_2 = -20; end
		5353: begin l_1 = -15;
				 l_2 = +20; end
		17718: begin l_1 = -15;
				 l_2 = -20; end
		4019: begin l_1 = +15;
				 l_2 = +21; end
		10136: begin l_1 = +15;
				 l_2 = -21; end
		8477: begin l_1 = -15;
				 l_2 = +21; end
		14594: begin l_1 = -15;
				 l_2 = -21; end
		10267: begin l_1 = +15;
				 l_2 = +22; end
		3888: begin l_1 = +15;
				 l_2 = -22; end
		14725: begin l_1 = -15;
				 l_2 = +22; end
		8346: begin l_1 = -15;
				 l_2 = -22; end
		4150: begin l_1 = +15;
				 l_2 = +23; end
		10005: begin l_1 = +15;
				 l_2 = -23; end
		8608: begin l_1 = -15;
				 l_2 = +23; end
		14463: begin l_1 = -15;
				 l_2 = -23; end
		10529: begin l_1 = +15;
				 l_2 = +24; end
		3626: begin l_1 = +15;
				 l_2 = -24; end
		14987: begin l_1 = -15;
				 l_2 = +24; end
		8084: begin l_1 = -15;
				 l_2 = -24; end
		4674: begin l_1 = +15;
				 l_2 = +25; end
		9481: begin l_1 = +15;
				 l_2 = -25; end
		9132: begin l_1 = -15;
				 l_2 = +25; end
		13939: begin l_1 = -15;
				 l_2 = -25; end
		11577: begin l_1 = +15;
				 l_2 = +26; end
		2578: begin l_1 = +15;
				 l_2 = -26; end
		16035: begin l_1 = -15;
				 l_2 = +26; end
		7036: begin l_1 = -15;
				 l_2 = -26; end
		6770: begin l_1 = +15;
				 l_2 = +27; end
		7385: begin l_1 = +15;
				 l_2 = -27; end
		11228: begin l_1 = -15;
				 l_2 = +27; end
		11843: begin l_1 = -15;
				 l_2 = -27; end
		15769: begin l_1 = +15;
				 l_2 = +28; end
		16999: begin l_1 = +15;
				 l_2 = -28; end
		1614: begin l_1 = -15;
				 l_2 = +28; end
		2844: begin l_1 = -15;
				 l_2 = -28; end
		15154: begin l_1 = +15;
				 l_2 = +29; end
		17614: begin l_1 = +15;
				 l_2 = -29; end
		999: begin l_1 = -15;
				 l_2 = +29; end
		3459: begin l_1 = -15;
				 l_2 = -29; end
		13924: begin l_1 = +15;
				 l_2 = +30; end
		231: begin l_1 = +15;
				 l_2 = -30; end
		18382: begin l_1 = -15;
				 l_2 = +30; end
		4689: begin l_1 = -15;
				 l_2 = -30; end
		11464: begin l_1 = +15;
				 l_2 = +31; end
		2691: begin l_1 = +15;
				 l_2 = -31; end
		15922: begin l_1 = -15;
				 l_2 = +31; end
		7149: begin l_1 = -15;
				 l_2 = -31; end
		6544: begin l_1 = +15;
				 l_2 = +32; end
		7611: begin l_1 = +15;
				 l_2 = -32; end
		11002: begin l_1 = -15;
				 l_2 = +32; end
		12069: begin l_1 = -15;
				 l_2 = -32; end
		15317: begin l_1 = +15;
				 l_2 = +33; end
		17451: begin l_1 = +15;
				 l_2 = -33; end
		1162: begin l_1 = -15;
				 l_2 = +33; end
		3296: begin l_1 = -15;
				 l_2 = -33; end
		14250: begin l_1 = +15;
				 l_2 = +34; end
		18518: begin l_1 = +15;
				 l_2 = -34; end
		95: begin l_1 = -15;
				 l_2 = +34; end
		4363: begin l_1 = -15;
				 l_2 = -34; end
		12116: begin l_1 = +15;
				 l_2 = +35; end
		2039: begin l_1 = +15;
				 l_2 = -35; end
		16574: begin l_1 = -15;
				 l_2 = +35; end
		6497: begin l_1 = -15;
				 l_2 = -35; end
		7848: begin l_1 = +15;
				 l_2 = +36; end
		6307: begin l_1 = +15;
				 l_2 = -36; end
		12306: begin l_1 = -15;
				 l_2 = +36; end
		10765: begin l_1 = -15;
				 l_2 = -36; end
		17925: begin l_1 = +15;
				 l_2 = +37; end
		14843: begin l_1 = +15;
				 l_2 = -37; end
		3770: begin l_1 = -15;
				 l_2 = +37; end
		688: begin l_1 = -15;
				 l_2 = -37; end
		853: begin l_1 = +15;
				 l_2 = +38; end
		13302: begin l_1 = +15;
				 l_2 = -38; end
		5311: begin l_1 = -15;
				 l_2 = +38; end
		17760: begin l_1 = -15;
				 l_2 = -38; end
		3935: begin l_1 = +15;
				 l_2 = +39; end
		10220: begin l_1 = +15;
				 l_2 = -39; end
		8393: begin l_1 = -15;
				 l_2 = +39; end
		14678: begin l_1 = -15;
				 l_2 = -39; end
		10099: begin l_1 = +15;
				 l_2 = +40; end
		4056: begin l_1 = +15;
				 l_2 = -40; end
		14557: begin l_1 = -15;
				 l_2 = +40; end
		8514: begin l_1 = -15;
				 l_2 = -40; end
		3814: begin l_1 = +15;
				 l_2 = +41; end
		10341: begin l_1 = +15;
				 l_2 = -41; end
		8272: begin l_1 = -15;
				 l_2 = +41; end
		14799: begin l_1 = -15;
				 l_2 = -41; end
		9857: begin l_1 = +15;
				 l_2 = +42; end
		4298: begin l_1 = +15;
				 l_2 = -42; end
		14315: begin l_1 = -15;
				 l_2 = +42; end
		8756: begin l_1 = -15;
				 l_2 = -42; end
		3330: begin l_1 = +15;
				 l_2 = +43; end
		10825: begin l_1 = +15;
				 l_2 = -43; end
		7788: begin l_1 = -15;
				 l_2 = +43; end
		15283: begin l_1 = -15;
				 l_2 = -43; end
		8889: begin l_1 = +15;
				 l_2 = +44; end
		5266: begin l_1 = +15;
				 l_2 = -44; end
		13347: begin l_1 = -15;
				 l_2 = +44; end
		9724: begin l_1 = -15;
				 l_2 = -44; end
		1394: begin l_1 = +15;
				 l_2 = +45; end
		12761: begin l_1 = +15;
				 l_2 = -45; end
		5852: begin l_1 = -15;
				 l_2 = +45; end
		17219: begin l_1 = -15;
				 l_2 = -45; end
		5239: begin l_1 = -16;
				 l_2 = +18; end
		13374: begin l_1 = -16;
				 l_2 = -17; end
		14936: begin l_1 = +16;
				 l_2 = +18; end
		3677: begin l_1 = -16;
				 l_2 = -18; end
		15717: begin l_1 = +16;
				 l_2 = +19; end
		12593: begin l_1 = +16;
				 l_2 = -19; end
		6020: begin l_1 = -16;
				 l_2 = +19; end
		2896: begin l_1 = -16;
				 l_2 = -19; end
		17279: begin l_1 = +16;
				 l_2 = +20; end
		11031: begin l_1 = +16;
				 l_2 = -20; end
		7582: begin l_1 = -16;
				 l_2 = +20; end
		1334: begin l_1 = -16;
				 l_2 = -20; end
		1790: begin l_1 = +16;
				 l_2 = +21; end
		7907: begin l_1 = +16;
				 l_2 = -21; end
		10706: begin l_1 = -16;
				 l_2 = +21; end
		16823: begin l_1 = -16;
				 l_2 = -21; end
		8038: begin l_1 = +16;
				 l_2 = +22; end
		1659: begin l_1 = +16;
				 l_2 = -22; end
		16954: begin l_1 = -16;
				 l_2 = +22; end
		10575: begin l_1 = -16;
				 l_2 = -22; end
		1921: begin l_1 = +16;
				 l_2 = +23; end
		7776: begin l_1 = +16;
				 l_2 = -23; end
		10837: begin l_1 = -16;
				 l_2 = +23; end
		16692: begin l_1 = -16;
				 l_2 = -23; end
		8300: begin l_1 = +16;
				 l_2 = +24; end
		1397: begin l_1 = +16;
				 l_2 = -24; end
		17216: begin l_1 = -16;
				 l_2 = +24; end
		10313: begin l_1 = -16;
				 l_2 = -24; end
		2445: begin l_1 = +16;
				 l_2 = +25; end
		7252: begin l_1 = +16;
				 l_2 = -25; end
		11361: begin l_1 = -16;
				 l_2 = +25; end
		16168: begin l_1 = -16;
				 l_2 = -25; end
		9348: begin l_1 = +16;
				 l_2 = +26; end
		349: begin l_1 = +16;
				 l_2 = -26; end
		18264: begin l_1 = -16;
				 l_2 = +26; end
		9265: begin l_1 = -16;
				 l_2 = -26; end
		4541: begin l_1 = +16;
				 l_2 = +27; end
		5156: begin l_1 = +16;
				 l_2 = -27; end
		13457: begin l_1 = -16;
				 l_2 = +27; end
		14072: begin l_1 = -16;
				 l_2 = -27; end
		13540: begin l_1 = +16;
				 l_2 = +28; end
		14770: begin l_1 = +16;
				 l_2 = -28; end
		3843: begin l_1 = -16;
				 l_2 = +28; end
		5073: begin l_1 = -16;
				 l_2 = -28; end
		12925: begin l_1 = +16;
				 l_2 = +29; end
		15385: begin l_1 = +16;
				 l_2 = -29; end
		3228: begin l_1 = -16;
				 l_2 = +29; end
		5688: begin l_1 = -16;
				 l_2 = -29; end
		11695: begin l_1 = +16;
				 l_2 = +30; end
		16615: begin l_1 = +16;
				 l_2 = -30; end
		1998: begin l_1 = -16;
				 l_2 = +30; end
		6918: begin l_1 = -16;
				 l_2 = -30; end
		9235: begin l_1 = +16;
				 l_2 = +31; end
		462: begin l_1 = +16;
				 l_2 = -31; end
		18151: begin l_1 = -16;
				 l_2 = +31; end
		9378: begin l_1 = -16;
				 l_2 = -31; end
		4315: begin l_1 = +16;
				 l_2 = +32; end
		5382: begin l_1 = +16;
				 l_2 = -32; end
		13231: begin l_1 = -16;
				 l_2 = +32; end
		14298: begin l_1 = -16;
				 l_2 = -32; end
		13088: begin l_1 = +16;
				 l_2 = +33; end
		15222: begin l_1 = +16;
				 l_2 = -33; end
		3391: begin l_1 = -16;
				 l_2 = +33; end
		5525: begin l_1 = -16;
				 l_2 = -33; end
		12021: begin l_1 = +16;
				 l_2 = +34; end
		16289: begin l_1 = +16;
				 l_2 = -34; end
		2324: begin l_1 = -16;
				 l_2 = +34; end
		6592: begin l_1 = -16;
				 l_2 = -34; end
		9887: begin l_1 = +16;
				 l_2 = +35; end
		18423: begin l_1 = +16;
				 l_2 = -35; end
		190: begin l_1 = -16;
				 l_2 = +35; end
		8726: begin l_1 = -16;
				 l_2 = -35; end
		5619: begin l_1 = +16;
				 l_2 = +36; end
		4078: begin l_1 = +16;
				 l_2 = -36; end
		14535: begin l_1 = -16;
				 l_2 = +36; end
		12994: begin l_1 = -16;
				 l_2 = -36; end
		15696: begin l_1 = +16;
				 l_2 = +37; end
		12614: begin l_1 = +16;
				 l_2 = -37; end
		5999: begin l_1 = -16;
				 l_2 = +37; end
		2917: begin l_1 = -16;
				 l_2 = -37; end
		17237: begin l_1 = +16;
				 l_2 = +38; end
		11073: begin l_1 = +16;
				 l_2 = -38; end
		7540: begin l_1 = -16;
				 l_2 = +38; end
		1376: begin l_1 = -16;
				 l_2 = -38; end
		1706: begin l_1 = +16;
				 l_2 = +39; end
		7991: begin l_1 = +16;
				 l_2 = -39; end
		10622: begin l_1 = -16;
				 l_2 = +39; end
		16907: begin l_1 = -16;
				 l_2 = -39; end
		7870: begin l_1 = +16;
				 l_2 = +40; end
		1827: begin l_1 = +16;
				 l_2 = -40; end
		16786: begin l_1 = -16;
				 l_2 = +40; end
		10743: begin l_1 = -16;
				 l_2 = -40; end
		1585: begin l_1 = +16;
				 l_2 = +41; end
		8112: begin l_1 = +16;
				 l_2 = -41; end
		10501: begin l_1 = -16;
				 l_2 = +41; end
		17028: begin l_1 = -16;
				 l_2 = -41; end
		7628: begin l_1 = +16;
				 l_2 = +42; end
		2069: begin l_1 = +16;
				 l_2 = -42; end
		16544: begin l_1 = -16;
				 l_2 = +42; end
		10985: begin l_1 = -16;
				 l_2 = -42; end
		1101: begin l_1 = +16;
				 l_2 = +43; end
		8596: begin l_1 = +16;
				 l_2 = -43; end
		10017: begin l_1 = -16;
				 l_2 = +43; end
		17512: begin l_1 = -16;
				 l_2 = -43; end
		6660: begin l_1 = +16;
				 l_2 = +44; end
		3037: begin l_1 = +16;
				 l_2 = -44; end
		15576: begin l_1 = -16;
				 l_2 = +44; end
		11953: begin l_1 = -16;
				 l_2 = -44; end
		17778: begin l_1 = +16;
				 l_2 = +45; end
		10532: begin l_1 = +16;
				 l_2 = -45; end
		8081: begin l_1 = -16;
				 l_2 = +45; end
		835: begin l_1 = -16;
				 l_2 = -45; end
		10478: begin l_1 = -17;
				 l_2 = +19; end
		8135: begin l_1 = -17;
				 l_2 = -18; end
		11259: begin l_1 = +17;
				 l_2 = +19; end
		7354: begin l_1 = -17;
				 l_2 = -19; end
		12821: begin l_1 = +17;
				 l_2 = +20; end
		6573: begin l_1 = +17;
				 l_2 = -20; end
		12040: begin l_1 = -17;
				 l_2 = +20; end
		5792: begin l_1 = -17;
				 l_2 = -20; end
		15945: begin l_1 = +17;
				 l_2 = +21; end
		3449: begin l_1 = +17;
				 l_2 = -21; end
		15164: begin l_1 = -17;
				 l_2 = +21; end
		2668: begin l_1 = -17;
				 l_2 = -21; end
		3580: begin l_1 = +17;
				 l_2 = +22; end
		15814: begin l_1 = +17;
				 l_2 = -22; end
		2799: begin l_1 = -17;
				 l_2 = +22; end
		15033: begin l_1 = -17;
				 l_2 = -22; end
		16076: begin l_1 = +17;
				 l_2 = +23; end
		3318: begin l_1 = +17;
				 l_2 = -23; end
		15295: begin l_1 = -17;
				 l_2 = +23; end
		2537: begin l_1 = -17;
				 l_2 = -23; end
		3842: begin l_1 = +17;
				 l_2 = +24; end
		15552: begin l_1 = +17;
				 l_2 = -24; end
		3061: begin l_1 = -17;
				 l_2 = +24; end
		14771: begin l_1 = -17;
				 l_2 = -24; end
		16600: begin l_1 = +17;
				 l_2 = +25; end
		2794: begin l_1 = +17;
				 l_2 = -25; end
		15819: begin l_1 = -17;
				 l_2 = +25; end
		2013: begin l_1 = -17;
				 l_2 = -25; end
		4890: begin l_1 = +17;
				 l_2 = +26; end
		14504: begin l_1 = +17;
				 l_2 = -26; end
		4109: begin l_1 = -17;
				 l_2 = +26; end
		13723: begin l_1 = -17;
				 l_2 = -26; end
		83: begin l_1 = +17;
				 l_2 = +27; end
		698: begin l_1 = +17;
				 l_2 = -27; end
		17915: begin l_1 = -17;
				 l_2 = +27; end
		18530: begin l_1 = -17;
				 l_2 = -27; end
		9082: begin l_1 = +17;
				 l_2 = +28; end
		10312: begin l_1 = +17;
				 l_2 = -28; end
		8301: begin l_1 = -17;
				 l_2 = +28; end
		9531: begin l_1 = -17;
				 l_2 = -28; end
		8467: begin l_1 = +17;
				 l_2 = +29; end
		10927: begin l_1 = +17;
				 l_2 = -29; end
		7686: begin l_1 = -17;
				 l_2 = +29; end
		10146: begin l_1 = -17;
				 l_2 = -29; end
		7237: begin l_1 = +17;
				 l_2 = +30; end
		12157: begin l_1 = +17;
				 l_2 = -30; end
		6456: begin l_1 = -17;
				 l_2 = +30; end
		11376: begin l_1 = -17;
				 l_2 = -30; end
		4777: begin l_1 = +17;
				 l_2 = +31; end
		14617: begin l_1 = +17;
				 l_2 = -31; end
		3996: begin l_1 = -17;
				 l_2 = +31; end
		13836: begin l_1 = -17;
				 l_2 = -31; end
		18470: begin l_1 = +17;
				 l_2 = +32; end
		924: begin l_1 = +17;
				 l_2 = -32; end
		17689: begin l_1 = -17;
				 l_2 = +32; end
		143: begin l_1 = -17;
				 l_2 = -32; end
		8630: begin l_1 = +17;
				 l_2 = +33; end
		10764: begin l_1 = +17;
				 l_2 = -33; end
		7849: begin l_1 = -17;
				 l_2 = +33; end
		9983: begin l_1 = -17;
				 l_2 = -33; end
		7563: begin l_1 = +17;
				 l_2 = +34; end
		11831: begin l_1 = +17;
				 l_2 = -34; end
		6782: begin l_1 = -17;
				 l_2 = +34; end
		11050: begin l_1 = -17;
				 l_2 = -34; end
		5429: begin l_1 = +17;
				 l_2 = +35; end
		13965: begin l_1 = +17;
				 l_2 = -35; end
		4648: begin l_1 = -17;
				 l_2 = +35; end
		13184: begin l_1 = -17;
				 l_2 = -35; end
		1161: begin l_1 = +17;
				 l_2 = +36; end
		18233: begin l_1 = +17;
				 l_2 = -36; end
		380: begin l_1 = -17;
				 l_2 = +36; end
		17452: begin l_1 = -17;
				 l_2 = -36; end
		11238: begin l_1 = +17;
				 l_2 = +37; end
		8156: begin l_1 = +17;
				 l_2 = -37; end
		10457: begin l_1 = -17;
				 l_2 = +37; end
		7375: begin l_1 = -17;
				 l_2 = -37; end
		12779: begin l_1 = +17;
				 l_2 = +38; end
		6615: begin l_1 = +17;
				 l_2 = -38; end
		11998: begin l_1 = -17;
				 l_2 = +38; end
		5834: begin l_1 = -17;
				 l_2 = -38; end
		15861: begin l_1 = +17;
				 l_2 = +39; end
		3533: begin l_1 = +17;
				 l_2 = -39; end
		15080: begin l_1 = -17;
				 l_2 = +39; end
		2752: begin l_1 = -17;
				 l_2 = -39; end
		3412: begin l_1 = +17;
				 l_2 = +40; end
		15982: begin l_1 = +17;
				 l_2 = -40; end
		2631: begin l_1 = -17;
				 l_2 = +40; end
		15201: begin l_1 = -17;
				 l_2 = -40; end
		15740: begin l_1 = +17;
				 l_2 = +41; end
		3654: begin l_1 = +17;
				 l_2 = -41; end
		14959: begin l_1 = -17;
				 l_2 = +41; end
		2873: begin l_1 = -17;
				 l_2 = -41; end
		3170: begin l_1 = +17;
				 l_2 = +42; end
		16224: begin l_1 = +17;
				 l_2 = -42; end
		2389: begin l_1 = -17;
				 l_2 = +42; end
		15443: begin l_1 = -17;
				 l_2 = -42; end
		15256: begin l_1 = +17;
				 l_2 = +43; end
		4138: begin l_1 = +17;
				 l_2 = -43; end
		14475: begin l_1 = -17;
				 l_2 = +43; end
		3357: begin l_1 = -17;
				 l_2 = -43; end
		2202: begin l_1 = +17;
				 l_2 = +44; end
		17192: begin l_1 = +17;
				 l_2 = -44; end
		1421: begin l_1 = -17;
				 l_2 = +44; end
		16411: begin l_1 = -17;
				 l_2 = -44; end
		13320: begin l_1 = +17;
				 l_2 = +45; end
		6074: begin l_1 = +17;
				 l_2 = -45; end
		12539: begin l_1 = -17;
				 l_2 = +45; end
		5293: begin l_1 = -17;
				 l_2 = -45; end
		2343: begin l_1 = -18;
				 l_2 = +20; end
		16270: begin l_1 = -18;
				 l_2 = -19; end
		3905: begin l_1 = +18;
				 l_2 = +20; end
		14708: begin l_1 = -18;
				 l_2 = -20; end
		7029: begin l_1 = +18;
				 l_2 = +21; end
		13146: begin l_1 = +18;
				 l_2 = -21; end
		5467: begin l_1 = -18;
				 l_2 = +21; end
		11584: begin l_1 = -18;
				 l_2 = -21; end
		13277: begin l_1 = +18;
				 l_2 = +22; end
		6898: begin l_1 = +18;
				 l_2 = -22; end
		11715: begin l_1 = -18;
				 l_2 = +22; end
		5336: begin l_1 = -18;
				 l_2 = -22; end
		7160: begin l_1 = +18;
				 l_2 = +23; end
		13015: begin l_1 = +18;
				 l_2 = -23; end
		5598: begin l_1 = -18;
				 l_2 = +23; end
		11453: begin l_1 = -18;
				 l_2 = -23; end
		13539: begin l_1 = +18;
				 l_2 = +24; end
		6636: begin l_1 = +18;
				 l_2 = -24; end
		11977: begin l_1 = -18;
				 l_2 = +24; end
		5074: begin l_1 = -18;
				 l_2 = -24; end
		7684: begin l_1 = +18;
				 l_2 = +25; end
		12491: begin l_1 = +18;
				 l_2 = -25; end
		6122: begin l_1 = -18;
				 l_2 = +25; end
		10929: begin l_1 = -18;
				 l_2 = -25; end
		14587: begin l_1 = +18;
				 l_2 = +26; end
		5588: begin l_1 = +18;
				 l_2 = -26; end
		13025: begin l_1 = -18;
				 l_2 = +26; end
		4026: begin l_1 = -18;
				 l_2 = -26; end
		9780: begin l_1 = +18;
				 l_2 = +27; end
		10395: begin l_1 = +18;
				 l_2 = -27; end
		8218: begin l_1 = -18;
				 l_2 = +27; end
		8833: begin l_1 = -18;
				 l_2 = -27; end
		166: begin l_1 = +18;
				 l_2 = +28; end
		1396: begin l_1 = +18;
				 l_2 = -28; end
		17217: begin l_1 = -18;
				 l_2 = +28; end
		18447: begin l_1 = -18;
				 l_2 = -28; end
		18164: begin l_1 = +18;
				 l_2 = +29; end
		2011: begin l_1 = +18;
				 l_2 = -29; end
		16602: begin l_1 = -18;
				 l_2 = +29; end
		449: begin l_1 = -18;
				 l_2 = -29; end
		16934: begin l_1 = +18;
				 l_2 = +30; end
		3241: begin l_1 = +18;
				 l_2 = -30; end
		15372: begin l_1 = -18;
				 l_2 = +30; end
		1679: begin l_1 = -18;
				 l_2 = -30; end
		14474: begin l_1 = +18;
				 l_2 = +31; end
		5701: begin l_1 = +18;
				 l_2 = -31; end
		12912: begin l_1 = -18;
				 l_2 = +31; end
		4139: begin l_1 = -18;
				 l_2 = -31; end
		9554: begin l_1 = +18;
				 l_2 = +32; end
		10621: begin l_1 = +18;
				 l_2 = -32; end
		7992: begin l_1 = -18;
				 l_2 = +32; end
		9059: begin l_1 = -18;
				 l_2 = -32; end
		18327: begin l_1 = +18;
				 l_2 = +33; end
		1848: begin l_1 = +18;
				 l_2 = -33; end
		16765: begin l_1 = -18;
				 l_2 = +33; end
		286: begin l_1 = -18;
				 l_2 = -33; end
		17260: begin l_1 = +18;
				 l_2 = +34; end
		2915: begin l_1 = +18;
				 l_2 = -34; end
		15698: begin l_1 = -18;
				 l_2 = +34; end
		1353: begin l_1 = -18;
				 l_2 = -34; end
		15126: begin l_1 = +18;
				 l_2 = +35; end
		5049: begin l_1 = +18;
				 l_2 = -35; end
		13564: begin l_1 = -18;
				 l_2 = +35; end
		3487: begin l_1 = -18;
				 l_2 = -35; end
		10858: begin l_1 = +18;
				 l_2 = +36; end
		9317: begin l_1 = +18;
				 l_2 = -36; end
		9296: begin l_1 = -18;
				 l_2 = +36; end
		7755: begin l_1 = -18;
				 l_2 = -36; end
		2322: begin l_1 = +18;
				 l_2 = +37; end
		17853: begin l_1 = +18;
				 l_2 = -37; end
		760: begin l_1 = -18;
				 l_2 = +37; end
		16291: begin l_1 = -18;
				 l_2 = -37; end
		3863: begin l_1 = +18;
				 l_2 = +38; end
		16312: begin l_1 = +18;
				 l_2 = -38; end
		2301: begin l_1 = -18;
				 l_2 = +38; end
		14750: begin l_1 = -18;
				 l_2 = -38; end
		6945: begin l_1 = +18;
				 l_2 = +39; end
		13230: begin l_1 = +18;
				 l_2 = -39; end
		5383: begin l_1 = -18;
				 l_2 = +39; end
		11668: begin l_1 = -18;
				 l_2 = -39; end
		13109: begin l_1 = +18;
				 l_2 = +40; end
		7066: begin l_1 = +18;
				 l_2 = -40; end
		11547: begin l_1 = -18;
				 l_2 = +40; end
		5504: begin l_1 = -18;
				 l_2 = -40; end
		6824: begin l_1 = +18;
				 l_2 = +41; end
		13351: begin l_1 = +18;
				 l_2 = -41; end
		5262: begin l_1 = -18;
				 l_2 = +41; end
		11789: begin l_1 = -18;
				 l_2 = -41; end
		12867: begin l_1 = +18;
				 l_2 = +42; end
		7308: begin l_1 = +18;
				 l_2 = -42; end
		11305: begin l_1 = -18;
				 l_2 = +42; end
		5746: begin l_1 = -18;
				 l_2 = -42; end
		6340: begin l_1 = +18;
				 l_2 = +43; end
		13835: begin l_1 = +18;
				 l_2 = -43; end
		4778: begin l_1 = -18;
				 l_2 = +43; end
		12273: begin l_1 = -18;
				 l_2 = -43; end
		11899: begin l_1 = +18;
				 l_2 = +44; end
		8276: begin l_1 = +18;
				 l_2 = -44; end
		10337: begin l_1 = -18;
				 l_2 = +44; end
		6714: begin l_1 = -18;
				 l_2 = -44; end
		4404: begin l_1 = +18;
				 l_2 = +45; end
		15771: begin l_1 = +18;
				 l_2 = -45; end
		2842: begin l_1 = -18;
				 l_2 = +45; end
		14209: begin l_1 = -18;
				 l_2 = -45; end
		4686: begin l_1 = -19;
				 l_2 = +21; end
		13927: begin l_1 = -19;
				 l_2 = -20; end
		7810: begin l_1 = +19;
				 l_2 = +21; end
		10803: begin l_1 = -19;
				 l_2 = -21; end
		14058: begin l_1 = +19;
				 l_2 = +22; end
		7679: begin l_1 = +19;
				 l_2 = -22; end
		10934: begin l_1 = -19;
				 l_2 = +22; end
		4555: begin l_1 = -19;
				 l_2 = -22; end
		7941: begin l_1 = +19;
				 l_2 = +23; end
		13796: begin l_1 = +19;
				 l_2 = -23; end
		4817: begin l_1 = -19;
				 l_2 = +23; end
		10672: begin l_1 = -19;
				 l_2 = -23; end
		14320: begin l_1 = +19;
				 l_2 = +24; end
		7417: begin l_1 = +19;
				 l_2 = -24; end
		11196: begin l_1 = -19;
				 l_2 = +24; end
		4293: begin l_1 = -19;
				 l_2 = -24; end
		8465: begin l_1 = +19;
				 l_2 = +25; end
		13272: begin l_1 = +19;
				 l_2 = -25; end
		5341: begin l_1 = -19;
				 l_2 = +25; end
		10148: begin l_1 = -19;
				 l_2 = -25; end
		15368: begin l_1 = +19;
				 l_2 = +26; end
		6369: begin l_1 = +19;
				 l_2 = -26; end
		12244: begin l_1 = -19;
				 l_2 = +26; end
		3245: begin l_1 = -19;
				 l_2 = -26; end
		10561: begin l_1 = +19;
				 l_2 = +27; end
		11176: begin l_1 = +19;
				 l_2 = -27; end
		7437: begin l_1 = -19;
				 l_2 = +27; end
		8052: begin l_1 = -19;
				 l_2 = -27; end
		947: begin l_1 = +19;
				 l_2 = +28; end
		2177: begin l_1 = +19;
				 l_2 = -28; end
		16436: begin l_1 = -19;
				 l_2 = +28; end
		17666: begin l_1 = -19;
				 l_2 = -28; end
		332: begin l_1 = +19;
				 l_2 = +29; end
		2792: begin l_1 = +19;
				 l_2 = -29; end
		15821: begin l_1 = -19;
				 l_2 = +29; end
		18281: begin l_1 = -19;
				 l_2 = -29; end
		17715: begin l_1 = +19;
				 l_2 = +30; end
		4022: begin l_1 = +19;
				 l_2 = -30; end
		14591: begin l_1 = -19;
				 l_2 = +30; end
		898: begin l_1 = -19;
				 l_2 = -30; end
		15255: begin l_1 = +19;
				 l_2 = +31; end
		6482: begin l_1 = +19;
				 l_2 = -31; end
		12131: begin l_1 = -19;
				 l_2 = +31; end
		3358: begin l_1 = -19;
				 l_2 = -31; end
		10335: begin l_1 = +19;
				 l_2 = +32; end
		11402: begin l_1 = +19;
				 l_2 = -32; end
		7211: begin l_1 = -19;
				 l_2 = +32; end
		8278: begin l_1 = -19;
				 l_2 = -32; end
		495: begin l_1 = +19;
				 l_2 = +33; end
		2629: begin l_1 = +19;
				 l_2 = -33; end
		15984: begin l_1 = -19;
				 l_2 = +33; end
		18118: begin l_1 = -19;
				 l_2 = -33; end
		18041: begin l_1 = +19;
				 l_2 = +34; end
		3696: begin l_1 = +19;
				 l_2 = -34; end
		14917: begin l_1 = -19;
				 l_2 = +34; end
		572: begin l_1 = -19;
				 l_2 = -34; end
		15907: begin l_1 = +19;
				 l_2 = +35; end
		5830: begin l_1 = +19;
				 l_2 = -35; end
		12783: begin l_1 = -19;
				 l_2 = +35; end
		2706: begin l_1 = -19;
				 l_2 = -35; end
		11639: begin l_1 = +19;
				 l_2 = +36; end
		10098: begin l_1 = +19;
				 l_2 = -36; end
		8515: begin l_1 = -19;
				 l_2 = +36; end
		6974: begin l_1 = -19;
				 l_2 = -36; end
		3103: begin l_1 = +19;
				 l_2 = +37; end
		21: begin l_1 = +19;
				 l_2 = -37; end
		18592: begin l_1 = -19;
				 l_2 = +37; end
		15510: begin l_1 = -19;
				 l_2 = -37; end
		4644: begin l_1 = +19;
				 l_2 = +38; end
		17093: begin l_1 = +19;
				 l_2 = -38; end
		1520: begin l_1 = -19;
				 l_2 = +38; end
		13969: begin l_1 = -19;
				 l_2 = -38; end
		7726: begin l_1 = +19;
				 l_2 = +39; end
		14011: begin l_1 = +19;
				 l_2 = -39; end
		4602: begin l_1 = -19;
				 l_2 = +39; end
		10887: begin l_1 = -19;
				 l_2 = -39; end
		13890: begin l_1 = +19;
				 l_2 = +40; end
		7847: begin l_1 = +19;
				 l_2 = -40; end
		10766: begin l_1 = -19;
				 l_2 = +40; end
		4723: begin l_1 = -19;
				 l_2 = -40; end
		7605: begin l_1 = +19;
				 l_2 = +41; end
		14132: begin l_1 = +19;
				 l_2 = -41; end
		4481: begin l_1 = -19;
				 l_2 = +41; end
		11008: begin l_1 = -19;
				 l_2 = -41; end
		13648: begin l_1 = +19;
				 l_2 = +42; end
		8089: begin l_1 = +19;
				 l_2 = -42; end
		10524: begin l_1 = -19;
				 l_2 = +42; end
		4965: begin l_1 = -19;
				 l_2 = -42; end
		7121: begin l_1 = +19;
				 l_2 = +43; end
		14616: begin l_1 = +19;
				 l_2 = -43; end
		3997: begin l_1 = -19;
				 l_2 = +43; end
		11492: begin l_1 = -19;
				 l_2 = -43; end
		12680: begin l_1 = +19;
				 l_2 = +44; end
		9057: begin l_1 = +19;
				 l_2 = -44; end
		9556: begin l_1 = -19;
				 l_2 = +44; end
		5933: begin l_1 = -19;
				 l_2 = -44; end
		5185: begin l_1 = +19;
				 l_2 = +45; end
		16552: begin l_1 = +19;
				 l_2 = -45; end
		2061: begin l_1 = -19;
				 l_2 = +45; end
		13428: begin l_1 = -19;
				 l_2 = -45; end
		9372: begin l_1 = -20;
				 l_2 = +22; end
		9241: begin l_1 = -20;
				 l_2 = -21; end
		15620: begin l_1 = +20;
				 l_2 = +22; end
		2993: begin l_1 = -20;
				 l_2 = -22; end
		9503: begin l_1 = +20;
				 l_2 = +23; end
		15358: begin l_1 = +20;
				 l_2 = -23; end
		3255: begin l_1 = -20;
				 l_2 = +23; end
		9110: begin l_1 = -20;
				 l_2 = -23; end
		15882: begin l_1 = +20;
				 l_2 = +24; end
		8979: begin l_1 = +20;
				 l_2 = -24; end
		9634: begin l_1 = -20;
				 l_2 = +24; end
		2731: begin l_1 = -20;
				 l_2 = -24; end
		10027: begin l_1 = +20;
				 l_2 = +25; end
		14834: begin l_1 = +20;
				 l_2 = -25; end
		3779: begin l_1 = -20;
				 l_2 = +25; end
		8586: begin l_1 = -20;
				 l_2 = -25; end
		16930: begin l_1 = +20;
				 l_2 = +26; end
		7931: begin l_1 = +20;
				 l_2 = -26; end
		10682: begin l_1 = -20;
				 l_2 = +26; end
		1683: begin l_1 = -20;
				 l_2 = -26; end
		12123: begin l_1 = +20;
				 l_2 = +27; end
		12738: begin l_1 = +20;
				 l_2 = -27; end
		5875: begin l_1 = -20;
				 l_2 = +27; end
		6490: begin l_1 = -20;
				 l_2 = -27; end
		2509: begin l_1 = +20;
				 l_2 = +28; end
		3739: begin l_1 = +20;
				 l_2 = -28; end
		14874: begin l_1 = -20;
				 l_2 = +28; end
		16104: begin l_1 = -20;
				 l_2 = -28; end
		1894: begin l_1 = +20;
				 l_2 = +29; end
		4354: begin l_1 = +20;
				 l_2 = -29; end
		14259: begin l_1 = -20;
				 l_2 = +29; end
		16719: begin l_1 = -20;
				 l_2 = -29; end
		664: begin l_1 = +20;
				 l_2 = +30; end
		5584: begin l_1 = +20;
				 l_2 = -30; end
		13029: begin l_1 = -20;
				 l_2 = +30; end
		17949: begin l_1 = -20;
				 l_2 = -30; end
		16817: begin l_1 = +20;
				 l_2 = +31; end
		8044: begin l_1 = +20;
				 l_2 = -31; end
		10569: begin l_1 = -20;
				 l_2 = +31; end
		1796: begin l_1 = -20;
				 l_2 = -31; end
		11897: begin l_1 = +20;
				 l_2 = +32; end
		12964: begin l_1 = +20;
				 l_2 = -32; end
		5649: begin l_1 = -20;
				 l_2 = +32; end
		6716: begin l_1 = -20;
				 l_2 = -32; end
		2057: begin l_1 = +20;
				 l_2 = +33; end
		4191: begin l_1 = +20;
				 l_2 = -33; end
		14422: begin l_1 = -20;
				 l_2 = +33; end
		16556: begin l_1 = -20;
				 l_2 = -33; end
		990: begin l_1 = +20;
				 l_2 = +34; end
		5258: begin l_1 = +20;
				 l_2 = -34; end
		13355: begin l_1 = -20;
				 l_2 = +34; end
		17623: begin l_1 = -20;
				 l_2 = -34; end
		17469: begin l_1 = +20;
				 l_2 = +35; end
		7392: begin l_1 = +20;
				 l_2 = -35; end
		11221: begin l_1 = -20;
				 l_2 = +35; end
		1144: begin l_1 = -20;
				 l_2 = -35; end
		13201: begin l_1 = +20;
				 l_2 = +36; end
		11660: begin l_1 = +20;
				 l_2 = -36; end
		6953: begin l_1 = -20;
				 l_2 = +36; end
		5412: begin l_1 = -20;
				 l_2 = -36; end
		4665: begin l_1 = +20;
				 l_2 = +37; end
		1583: begin l_1 = +20;
				 l_2 = -37; end
		17030: begin l_1 = -20;
				 l_2 = +37; end
		13948: begin l_1 = -20;
				 l_2 = -37; end
		6206: begin l_1 = +20;
				 l_2 = +38; end
		42: begin l_1 = +20;
				 l_2 = -38; end
		18571: begin l_1 = -20;
				 l_2 = +38; end
		12407: begin l_1 = -20;
				 l_2 = -38; end
		9288: begin l_1 = +20;
				 l_2 = +39; end
		15573: begin l_1 = +20;
				 l_2 = -39; end
		3040: begin l_1 = -20;
				 l_2 = +39; end
		9325: begin l_1 = -20;
				 l_2 = -39; end
		15452: begin l_1 = +20;
				 l_2 = +40; end
		9409: begin l_1 = +20;
				 l_2 = -40; end
		9204: begin l_1 = -20;
				 l_2 = +40; end
		3161: begin l_1 = -20;
				 l_2 = -40; end
		9167: begin l_1 = +20;
				 l_2 = +41; end
		15694: begin l_1 = +20;
				 l_2 = -41; end
		2919: begin l_1 = -20;
				 l_2 = +41; end
		9446: begin l_1 = -20;
				 l_2 = -41; end
		15210: begin l_1 = +20;
				 l_2 = +42; end
		9651: begin l_1 = +20;
				 l_2 = -42; end
		8962: begin l_1 = -20;
				 l_2 = +42; end
		3403: begin l_1 = -20;
				 l_2 = -42; end
		8683: begin l_1 = +20;
				 l_2 = +43; end
		16178: begin l_1 = +20;
				 l_2 = -43; end
		2435: begin l_1 = -20;
				 l_2 = +43; end
		9930: begin l_1 = -20;
				 l_2 = -43; end
		14242: begin l_1 = +20;
				 l_2 = +44; end
		10619: begin l_1 = +20;
				 l_2 = -44; end
		7994: begin l_1 = -20;
				 l_2 = +44; end
		4371: begin l_1 = -20;
				 l_2 = -44; end
		6747: begin l_1 = +20;
				 l_2 = +45; end
		18114: begin l_1 = +20;
				 l_2 = -45; end
		499: begin l_1 = -20;
				 l_2 = +45; end
		11866: begin l_1 = -20;
				 l_2 = -45; end
		131: begin l_1 = -21;
				 l_2 = +23; end
		18482: begin l_1 = -21;
				 l_2 = -22; end
		12627: begin l_1 = +21;
				 l_2 = +23; end
		5986: begin l_1 = -21;
				 l_2 = -23; end
		393: begin l_1 = +21;
				 l_2 = +24; end
		12103: begin l_1 = +21;
				 l_2 = -24; end
		6510: begin l_1 = -21;
				 l_2 = +24; end
		18220: begin l_1 = -21;
				 l_2 = -24; end
		13151: begin l_1 = +21;
				 l_2 = +25; end
		17958: begin l_1 = +21;
				 l_2 = -25; end
		655: begin l_1 = -21;
				 l_2 = +25; end
		5462: begin l_1 = -21;
				 l_2 = -25; end
		1441: begin l_1 = +21;
				 l_2 = +26; end
		11055: begin l_1 = +21;
				 l_2 = -26; end
		7558: begin l_1 = -21;
				 l_2 = +26; end
		17172: begin l_1 = -21;
				 l_2 = -26; end
		15247: begin l_1 = +21;
				 l_2 = +27; end
		15862: begin l_1 = +21;
				 l_2 = -27; end
		2751: begin l_1 = -21;
				 l_2 = +27; end
		3366: begin l_1 = -21;
				 l_2 = -27; end
		5633: begin l_1 = +21;
				 l_2 = +28; end
		6863: begin l_1 = +21;
				 l_2 = -28; end
		11750: begin l_1 = -21;
				 l_2 = +28; end
		12980: begin l_1 = -21;
				 l_2 = -28; end
		5018: begin l_1 = +21;
				 l_2 = +29; end
		7478: begin l_1 = +21;
				 l_2 = -29; end
		11135: begin l_1 = -21;
				 l_2 = +29; end
		13595: begin l_1 = -21;
				 l_2 = -29; end
		3788: begin l_1 = +21;
				 l_2 = +30; end
		8708: begin l_1 = +21;
				 l_2 = -30; end
		9905: begin l_1 = -21;
				 l_2 = +30; end
		14825: begin l_1 = -21;
				 l_2 = -30; end
		1328: begin l_1 = +21;
				 l_2 = +31; end
		11168: begin l_1 = +21;
				 l_2 = -31; end
		7445: begin l_1 = -21;
				 l_2 = +31; end
		17285: begin l_1 = -21;
				 l_2 = -31; end
		15021: begin l_1 = +21;
				 l_2 = +32; end
		16088: begin l_1 = +21;
				 l_2 = -32; end
		2525: begin l_1 = -21;
				 l_2 = +32; end
		3592: begin l_1 = -21;
				 l_2 = -32; end
		5181: begin l_1 = +21;
				 l_2 = +33; end
		7315: begin l_1 = +21;
				 l_2 = -33; end
		11298: begin l_1 = -21;
				 l_2 = +33; end
		13432: begin l_1 = -21;
				 l_2 = -33; end
		4114: begin l_1 = +21;
				 l_2 = +34; end
		8382: begin l_1 = +21;
				 l_2 = -34; end
		10231: begin l_1 = -21;
				 l_2 = +34; end
		14499: begin l_1 = -21;
				 l_2 = -34; end
		1980: begin l_1 = +21;
				 l_2 = +35; end
		10516: begin l_1 = +21;
				 l_2 = -35; end
		8097: begin l_1 = -21;
				 l_2 = +35; end
		16633: begin l_1 = -21;
				 l_2 = -35; end
		16325: begin l_1 = +21;
				 l_2 = +36; end
		14784: begin l_1 = +21;
				 l_2 = -36; end
		3829: begin l_1 = -21;
				 l_2 = +36; end
		2288: begin l_1 = -21;
				 l_2 = -36; end
		7789: begin l_1 = +21;
				 l_2 = +37; end
		4707: begin l_1 = +21;
				 l_2 = -37; end
		13906: begin l_1 = -21;
				 l_2 = +37; end
		10824: begin l_1 = -21;
				 l_2 = -37; end
		9330: begin l_1 = +21;
				 l_2 = +38; end
		3166: begin l_1 = +21;
				 l_2 = -38; end
		15447: begin l_1 = -21;
				 l_2 = +38; end
		9283: begin l_1 = -21;
				 l_2 = -38; end
		12412: begin l_1 = +21;
				 l_2 = +39; end
		84: begin l_1 = +21;
				 l_2 = -39; end
		18529: begin l_1 = -21;
				 l_2 = +39; end
		6201: begin l_1 = -21;
				 l_2 = -39; end
		18576: begin l_1 = +21;
				 l_2 = +40; end
		12533: begin l_1 = +21;
				 l_2 = -40; end
		6080: begin l_1 = -21;
				 l_2 = +40; end
		37: begin l_1 = -21;
				 l_2 = -40; end
		12291: begin l_1 = +21;
				 l_2 = +41; end
		205: begin l_1 = +21;
				 l_2 = -41; end
		18408: begin l_1 = -21;
				 l_2 = +41; end
		6322: begin l_1 = -21;
				 l_2 = -41; end
		18334: begin l_1 = +21;
				 l_2 = +42; end
		12775: begin l_1 = +21;
				 l_2 = -42; end
		5838: begin l_1 = -21;
				 l_2 = +42; end
		279: begin l_1 = -21;
				 l_2 = -42; end
		11807: begin l_1 = +21;
				 l_2 = +43; end
		689: begin l_1 = +21;
				 l_2 = -43; end
		17924: begin l_1 = -21;
				 l_2 = +43; end
		6806: begin l_1 = -21;
				 l_2 = -43; end
		17366: begin l_1 = +21;
				 l_2 = +44; end
		13743: begin l_1 = +21;
				 l_2 = -44; end
		4870: begin l_1 = -21;
				 l_2 = +44; end
		1247: begin l_1 = -21;
				 l_2 = -44; end
		9871: begin l_1 = +21;
				 l_2 = +45; end
		2625: begin l_1 = +21;
				 l_2 = -45; end
		15988: begin l_1 = -21;
				 l_2 = +45; end
		8742: begin l_1 = -21;
				 l_2 = -45; end
		262: begin l_1 = -22;
				 l_2 = +24; end
		18351: begin l_1 = -22;
				 l_2 = -23; end
		6641: begin l_1 = +22;
				 l_2 = +24; end
		11972: begin l_1 = -22;
				 l_2 = -24; end
		786: begin l_1 = +22;
				 l_2 = +25; end
		5593: begin l_1 = +22;
				 l_2 = -25; end
		13020: begin l_1 = -22;
				 l_2 = +25; end
		17827: begin l_1 = -22;
				 l_2 = -25; end
		7689: begin l_1 = +22;
				 l_2 = +26; end
		17303: begin l_1 = +22;
				 l_2 = -26; end
		1310: begin l_1 = -22;
				 l_2 = +26; end
		10924: begin l_1 = -22;
				 l_2 = -26; end
		2882: begin l_1 = +22;
				 l_2 = +27; end
		3497: begin l_1 = +22;
				 l_2 = -27; end
		15116: begin l_1 = -22;
				 l_2 = +27; end
		15731: begin l_1 = -22;
				 l_2 = -27; end
		11881: begin l_1 = +22;
				 l_2 = +28; end
		13111: begin l_1 = +22;
				 l_2 = -28; end
		5502: begin l_1 = -22;
				 l_2 = +28; end
		6732: begin l_1 = -22;
				 l_2 = -28; end
		11266: begin l_1 = +22;
				 l_2 = +29; end
		13726: begin l_1 = +22;
				 l_2 = -29; end
		4887: begin l_1 = -22;
				 l_2 = +29; end
		7347: begin l_1 = -22;
				 l_2 = -29; end
		10036: begin l_1 = +22;
				 l_2 = +30; end
		14956: begin l_1 = +22;
				 l_2 = -30; end
		3657: begin l_1 = -22;
				 l_2 = +30; end
		8577: begin l_1 = -22;
				 l_2 = -30; end
		7576: begin l_1 = +22;
				 l_2 = +31; end
		17416: begin l_1 = +22;
				 l_2 = -31; end
		1197: begin l_1 = -22;
				 l_2 = +31; end
		11037: begin l_1 = -22;
				 l_2 = -31; end
		2656: begin l_1 = +22;
				 l_2 = +32; end
		3723: begin l_1 = +22;
				 l_2 = -32; end
		14890: begin l_1 = -22;
				 l_2 = +32; end
		15957: begin l_1 = -22;
				 l_2 = -32; end
		11429: begin l_1 = +22;
				 l_2 = +33; end
		13563: begin l_1 = +22;
				 l_2 = -33; end
		5050: begin l_1 = -22;
				 l_2 = +33; end
		7184: begin l_1 = -22;
				 l_2 = -33; end
		10362: begin l_1 = +22;
				 l_2 = +34; end
		14630: begin l_1 = +22;
				 l_2 = -34; end
		3983: begin l_1 = -22;
				 l_2 = +34; end
		8251: begin l_1 = -22;
				 l_2 = -34; end
		8228: begin l_1 = +22;
				 l_2 = +35; end
		16764: begin l_1 = +22;
				 l_2 = -35; end
		1849: begin l_1 = -22;
				 l_2 = +35; end
		10385: begin l_1 = -22;
				 l_2 = -35; end
		3960: begin l_1 = +22;
				 l_2 = +36; end
		2419: begin l_1 = +22;
				 l_2 = -36; end
		16194: begin l_1 = -22;
				 l_2 = +36; end
		14653: begin l_1 = -22;
				 l_2 = -36; end
		14037: begin l_1 = +22;
				 l_2 = +37; end
		10955: begin l_1 = +22;
				 l_2 = -37; end
		7658: begin l_1 = -22;
				 l_2 = +37; end
		4576: begin l_1 = -22;
				 l_2 = -37; end
		15578: begin l_1 = +22;
				 l_2 = +38; end
		9414: begin l_1 = +22;
				 l_2 = -38; end
		9199: begin l_1 = -22;
				 l_2 = +38; end
		3035: begin l_1 = -22;
				 l_2 = -38; end
		47: begin l_1 = +22;
				 l_2 = +39; end
		6332: begin l_1 = +22;
				 l_2 = -39; end
		12281: begin l_1 = -22;
				 l_2 = +39; end
		18566: begin l_1 = -22;
				 l_2 = -39; end
		6211: begin l_1 = +22;
				 l_2 = +40; end
		168: begin l_1 = +22;
				 l_2 = -40; end
		18445: begin l_1 = -22;
				 l_2 = +40; end
		12402: begin l_1 = -22;
				 l_2 = -40; end
		18539: begin l_1 = +22;
				 l_2 = +41; end
		6453: begin l_1 = +22;
				 l_2 = -41; end
		12160: begin l_1 = -22;
				 l_2 = +41; end
		74: begin l_1 = -22;
				 l_2 = -41; end
		5969: begin l_1 = +22;
				 l_2 = +42; end
		410: begin l_1 = +22;
				 l_2 = -42; end
		18203: begin l_1 = -22;
				 l_2 = +42; end
		12644: begin l_1 = -22;
				 l_2 = -42; end
		18055: begin l_1 = +22;
				 l_2 = +43; end
		6937: begin l_1 = +22;
				 l_2 = -43; end
		11676: begin l_1 = -22;
				 l_2 = +43; end
		558: begin l_1 = -22;
				 l_2 = -43; end
		5001: begin l_1 = +22;
				 l_2 = +44; end
		1378: begin l_1 = +22;
				 l_2 = -44; end
		17235: begin l_1 = -22;
				 l_2 = +44; end
		13612: begin l_1 = -22;
				 l_2 = -44; end
		16119: begin l_1 = +22;
				 l_2 = +45; end
		8873: begin l_1 = +22;
				 l_2 = -45; end
		9740: begin l_1 = -22;
				 l_2 = +45; end
		2494: begin l_1 = -22;
				 l_2 = -45; end
		524: begin l_1 = -23;
				 l_2 = +25; end
		18089: begin l_1 = -23;
				 l_2 = -24; end
		13282: begin l_1 = +23;
				 l_2 = +25; end
		5331: begin l_1 = -23;
				 l_2 = -25; end
		1572: begin l_1 = +23;
				 l_2 = +26; end
		11186: begin l_1 = +23;
				 l_2 = -26; end
		7427: begin l_1 = -23;
				 l_2 = +26; end
		17041: begin l_1 = -23;
				 l_2 = -26; end
		15378: begin l_1 = +23;
				 l_2 = +27; end
		15993: begin l_1 = +23;
				 l_2 = -27; end
		2620: begin l_1 = -23;
				 l_2 = +27; end
		3235: begin l_1 = -23;
				 l_2 = -27; end
		5764: begin l_1 = +23;
				 l_2 = +28; end
		6994: begin l_1 = +23;
				 l_2 = -28; end
		11619: begin l_1 = -23;
				 l_2 = +28; end
		12849: begin l_1 = -23;
				 l_2 = -28; end
		5149: begin l_1 = +23;
				 l_2 = +29; end
		7609: begin l_1 = +23;
				 l_2 = -29; end
		11004: begin l_1 = -23;
				 l_2 = +29; end
		13464: begin l_1 = -23;
				 l_2 = -29; end
		3919: begin l_1 = +23;
				 l_2 = +30; end
		8839: begin l_1 = +23;
				 l_2 = -30; end
		9774: begin l_1 = -23;
				 l_2 = +30; end
		14694: begin l_1 = -23;
				 l_2 = -30; end
		1459: begin l_1 = +23;
				 l_2 = +31; end
		11299: begin l_1 = +23;
				 l_2 = -31; end
		7314: begin l_1 = -23;
				 l_2 = +31; end
		17154: begin l_1 = -23;
				 l_2 = -31; end
		15152: begin l_1 = +23;
				 l_2 = +32; end
		16219: begin l_1 = +23;
				 l_2 = -32; end
		2394: begin l_1 = -23;
				 l_2 = +32; end
		3461: begin l_1 = -23;
				 l_2 = -32; end
		5312: begin l_1 = +23;
				 l_2 = +33; end
		7446: begin l_1 = +23;
				 l_2 = -33; end
		11167: begin l_1 = -23;
				 l_2 = +33; end
		13301: begin l_1 = -23;
				 l_2 = -33; end
		4245: begin l_1 = +23;
				 l_2 = +34; end
		8513: begin l_1 = +23;
				 l_2 = -34; end
		10100: begin l_1 = -23;
				 l_2 = +34; end
		14368: begin l_1 = -23;
				 l_2 = -34; end
		2111: begin l_1 = +23;
				 l_2 = +35; end
		10647: begin l_1 = +23;
				 l_2 = -35; end
		7966: begin l_1 = -23;
				 l_2 = +35; end
		16502: begin l_1 = -23;
				 l_2 = -35; end
		16456: begin l_1 = +23;
				 l_2 = +36; end
		14915: begin l_1 = +23;
				 l_2 = -36; end
		3698: begin l_1 = -23;
				 l_2 = +36; end
		2157: begin l_1 = -23;
				 l_2 = -36; end
		7920: begin l_1 = +23;
				 l_2 = +37; end
		4838: begin l_1 = +23;
				 l_2 = -37; end
		13775: begin l_1 = -23;
				 l_2 = +37; end
		10693: begin l_1 = -23;
				 l_2 = -37; end
		9461: begin l_1 = +23;
				 l_2 = +38; end
		3297: begin l_1 = +23;
				 l_2 = -38; end
		15316: begin l_1 = -23;
				 l_2 = +38; end
		9152: begin l_1 = -23;
				 l_2 = -38; end
		12543: begin l_1 = +23;
				 l_2 = +39; end
		215: begin l_1 = +23;
				 l_2 = -39; end
		18398: begin l_1 = -23;
				 l_2 = +39; end
		6070: begin l_1 = -23;
				 l_2 = -39; end
		94: begin l_1 = +23;
				 l_2 = +40; end
		12664: begin l_1 = +23;
				 l_2 = -40; end
		5949: begin l_1 = -23;
				 l_2 = +40; end
		18519: begin l_1 = -23;
				 l_2 = -40; end
		12422: begin l_1 = +23;
				 l_2 = +41; end
		336: begin l_1 = +23;
				 l_2 = -41; end
		18277: begin l_1 = -23;
				 l_2 = +41; end
		6191: begin l_1 = -23;
				 l_2 = -41; end
		18465: begin l_1 = +23;
				 l_2 = +42; end
		12906: begin l_1 = +23;
				 l_2 = -42; end
		5707: begin l_1 = -23;
				 l_2 = +42; end
		148: begin l_1 = -23;
				 l_2 = -42; end
		11938: begin l_1 = +23;
				 l_2 = +43; end
		820: begin l_1 = +23;
				 l_2 = -43; end
		17793: begin l_1 = -23;
				 l_2 = +43; end
		6675: begin l_1 = -23;
				 l_2 = -43; end
		17497: begin l_1 = +23;
				 l_2 = +44; end
		13874: begin l_1 = +23;
				 l_2 = -44; end
		4739: begin l_1 = -23;
				 l_2 = +44; end
		1116: begin l_1 = -23;
				 l_2 = -44; end
		10002: begin l_1 = +23;
				 l_2 = +45; end
		2756: begin l_1 = +23;
				 l_2 = -45; end
		15857: begin l_1 = -23;
				 l_2 = +45; end
		8611: begin l_1 = -23;
				 l_2 = -45; end
		1048: begin l_1 = -24;
				 l_2 = +26; end
		17565: begin l_1 = -24;
				 l_2 = -25; end
		7951: begin l_1 = +24;
				 l_2 = +26; end
		10662: begin l_1 = -24;
				 l_2 = -26; end
		3144: begin l_1 = +24;
				 l_2 = +27; end
		3759: begin l_1 = +24;
				 l_2 = -27; end
		14854: begin l_1 = -24;
				 l_2 = +27; end
		15469: begin l_1 = -24;
				 l_2 = -27; end
		12143: begin l_1 = +24;
				 l_2 = +28; end
		13373: begin l_1 = +24;
				 l_2 = -28; end
		5240: begin l_1 = -24;
				 l_2 = +28; end
		6470: begin l_1 = -24;
				 l_2 = -28; end
		11528: begin l_1 = +24;
				 l_2 = +29; end
		13988: begin l_1 = +24;
				 l_2 = -29; end
		4625: begin l_1 = -24;
				 l_2 = +29; end
		7085: begin l_1 = -24;
				 l_2 = -29; end
		10298: begin l_1 = +24;
				 l_2 = +30; end
		15218: begin l_1 = +24;
				 l_2 = -30; end
		3395: begin l_1 = -24;
				 l_2 = +30; end
		8315: begin l_1 = -24;
				 l_2 = -30; end
		7838: begin l_1 = +24;
				 l_2 = +31; end
		17678: begin l_1 = +24;
				 l_2 = -31; end
		935: begin l_1 = -24;
				 l_2 = +31; end
		10775: begin l_1 = -24;
				 l_2 = -31; end
		2918: begin l_1 = +24;
				 l_2 = +32; end
		3985: begin l_1 = +24;
				 l_2 = -32; end
		14628: begin l_1 = -24;
				 l_2 = +32; end
		15695: begin l_1 = -24;
				 l_2 = -32; end
		11691: begin l_1 = +24;
				 l_2 = +33; end
		13825: begin l_1 = +24;
				 l_2 = -33; end
		4788: begin l_1 = -24;
				 l_2 = +33; end
		6922: begin l_1 = -24;
				 l_2 = -33; end
		10624: begin l_1 = +24;
				 l_2 = +34; end
		14892: begin l_1 = +24;
				 l_2 = -34; end
		3721: begin l_1 = -24;
				 l_2 = +34; end
		7989: begin l_1 = -24;
				 l_2 = -34; end
		8490: begin l_1 = +24;
				 l_2 = +35; end
		17026: begin l_1 = +24;
				 l_2 = -35; end
		1587: begin l_1 = -24;
				 l_2 = +35; end
		10123: begin l_1 = -24;
				 l_2 = -35; end
		4222: begin l_1 = +24;
				 l_2 = +36; end
		2681: begin l_1 = +24;
				 l_2 = -36; end
		15932: begin l_1 = -24;
				 l_2 = +36; end
		14391: begin l_1 = -24;
				 l_2 = -36; end
		14299: begin l_1 = +24;
				 l_2 = +37; end
		11217: begin l_1 = +24;
				 l_2 = -37; end
		7396: begin l_1 = -24;
				 l_2 = +37; end
		4314: begin l_1 = -24;
				 l_2 = -37; end
		15840: begin l_1 = +24;
				 l_2 = +38; end
		9676: begin l_1 = +24;
				 l_2 = -38; end
		8937: begin l_1 = -24;
				 l_2 = +38; end
		2773: begin l_1 = -24;
				 l_2 = -38; end
		309: begin l_1 = +24;
				 l_2 = +39; end
		6594: begin l_1 = +24;
				 l_2 = -39; end
		12019: begin l_1 = -24;
				 l_2 = +39; end
		18304: begin l_1 = -24;
				 l_2 = -39; end
		6473: begin l_1 = +24;
				 l_2 = +40; end
		430: begin l_1 = +24;
				 l_2 = -40; end
		18183: begin l_1 = -24;
				 l_2 = +40; end
		12140: begin l_1 = -24;
				 l_2 = -40; end
		188: begin l_1 = +24;
				 l_2 = +41; end
		6715: begin l_1 = +24;
				 l_2 = -41; end
		11898: begin l_1 = -24;
				 l_2 = +41; end
		18425: begin l_1 = -24;
				 l_2 = -41; end
		6231: begin l_1 = +24;
				 l_2 = +42; end
		672: begin l_1 = +24;
				 l_2 = -42; end
		17941: begin l_1 = -24;
				 l_2 = +42; end
		12382: begin l_1 = -24;
				 l_2 = -42; end
		18317: begin l_1 = +24;
				 l_2 = +43; end
		7199: begin l_1 = +24;
				 l_2 = -43; end
		11414: begin l_1 = -24;
				 l_2 = +43; end
		296: begin l_1 = -24;
				 l_2 = -43; end
		5263: begin l_1 = +24;
				 l_2 = +44; end
		1640: begin l_1 = +24;
				 l_2 = -44; end
		16973: begin l_1 = -24;
				 l_2 = +44; end
		13350: begin l_1 = -24;
				 l_2 = -44; end
		16381: begin l_1 = +24;
				 l_2 = +45; end
		9135: begin l_1 = +24;
				 l_2 = -45; end
		9478: begin l_1 = -24;
				 l_2 = +45; end
		2232: begin l_1 = -24;
				 l_2 = -45; end
		2096: begin l_1 = -25;
				 l_2 = +27; end
		16517: begin l_1 = -25;
				 l_2 = -26; end
		15902: begin l_1 = +25;
				 l_2 = +27; end
		2711: begin l_1 = -25;
				 l_2 = -27; end
		6288: begin l_1 = +25;
				 l_2 = +28; end
		7518: begin l_1 = +25;
				 l_2 = -28; end
		11095: begin l_1 = -25;
				 l_2 = +28; end
		12325: begin l_1 = -25;
				 l_2 = -28; end
		5673: begin l_1 = +25;
				 l_2 = +29; end
		8133: begin l_1 = +25;
				 l_2 = -29; end
		10480: begin l_1 = -25;
				 l_2 = +29; end
		12940: begin l_1 = -25;
				 l_2 = -29; end
		4443: begin l_1 = +25;
				 l_2 = +30; end
		9363: begin l_1 = +25;
				 l_2 = -30; end
		9250: begin l_1 = -25;
				 l_2 = +30; end
		14170: begin l_1 = -25;
				 l_2 = -30; end
		1983: begin l_1 = +25;
				 l_2 = +31; end
		11823: begin l_1 = +25;
				 l_2 = -31; end
		6790: begin l_1 = -25;
				 l_2 = +31; end
		16630: begin l_1 = -25;
				 l_2 = -31; end
		15676: begin l_1 = +25;
				 l_2 = +32; end
		16743: begin l_1 = +25;
				 l_2 = -32; end
		1870: begin l_1 = -25;
				 l_2 = +32; end
		2937: begin l_1 = -25;
				 l_2 = -32; end
		5836: begin l_1 = +25;
				 l_2 = +33; end
		7970: begin l_1 = +25;
				 l_2 = -33; end
		10643: begin l_1 = -25;
				 l_2 = +33; end
		12777: begin l_1 = -25;
				 l_2 = -33; end
		4769: begin l_1 = +25;
				 l_2 = +34; end
		9037: begin l_1 = +25;
				 l_2 = -34; end
		9576: begin l_1 = -25;
				 l_2 = +34; end
		13844: begin l_1 = -25;
				 l_2 = -34; end
		2635: begin l_1 = +25;
				 l_2 = +35; end
		11171: begin l_1 = +25;
				 l_2 = -35; end
		7442: begin l_1 = -25;
				 l_2 = +35; end
		15978: begin l_1 = -25;
				 l_2 = -35; end
		16980: begin l_1 = +25;
				 l_2 = +36; end
		15439: begin l_1 = +25;
				 l_2 = -36; end
		3174: begin l_1 = -25;
				 l_2 = +36; end
		1633: begin l_1 = -25;
				 l_2 = -36; end
		8444: begin l_1 = +25;
				 l_2 = +37; end
		5362: begin l_1 = +25;
				 l_2 = -37; end
		13251: begin l_1 = -25;
				 l_2 = +37; end
		10169: begin l_1 = -25;
				 l_2 = -37; end
		9985: begin l_1 = +25;
				 l_2 = +38; end
		3821: begin l_1 = +25;
				 l_2 = -38; end
		14792: begin l_1 = -25;
				 l_2 = +38; end
		8628: begin l_1 = -25;
				 l_2 = -38; end
		13067: begin l_1 = +25;
				 l_2 = +39; end
		739: begin l_1 = +25;
				 l_2 = -39; end
		17874: begin l_1 = -25;
				 l_2 = +39; end
		5546: begin l_1 = -25;
				 l_2 = -39; end
		618: begin l_1 = +25;
				 l_2 = +40; end
		13188: begin l_1 = +25;
				 l_2 = -40; end
		5425: begin l_1 = -25;
				 l_2 = +40; end
		17995: begin l_1 = -25;
				 l_2 = -40; end
		12946: begin l_1 = +25;
				 l_2 = +41; end
		860: begin l_1 = +25;
				 l_2 = -41; end
		17753: begin l_1 = -25;
				 l_2 = +41; end
		5667: begin l_1 = -25;
				 l_2 = -41; end
		376: begin l_1 = +25;
				 l_2 = +42; end
		13430: begin l_1 = +25;
				 l_2 = -42; end
		5183: begin l_1 = -25;
				 l_2 = +42; end
		18237: begin l_1 = -25;
				 l_2 = -42; end
		12462: begin l_1 = +25;
				 l_2 = +43; end
		1344: begin l_1 = +25;
				 l_2 = -43; end
		17269: begin l_1 = -25;
				 l_2 = +43; end
		6151: begin l_1 = -25;
				 l_2 = -43; end
		18021: begin l_1 = +25;
				 l_2 = +44; end
		14398: begin l_1 = +25;
				 l_2 = -44; end
		4215: begin l_1 = -25;
				 l_2 = +44; end
		592: begin l_1 = -25;
				 l_2 = -44; end
		10526: begin l_1 = +25;
				 l_2 = +45; end
		3280: begin l_1 = +25;
				 l_2 = -45; end
		15333: begin l_1 = -25;
				 l_2 = +45; end
		8087: begin l_1 = -25;
				 l_2 = -45; end
		4192: begin l_1 = -26;
				 l_2 = +28; end
		14421: begin l_1 = -26;
				 l_2 = -27; end
		13191: begin l_1 = +26;
				 l_2 = +28; end
		5422: begin l_1 = -26;
				 l_2 = -28; end
		12576: begin l_1 = +26;
				 l_2 = +29; end
		15036: begin l_1 = +26;
				 l_2 = -29; end
		3577: begin l_1 = -26;
				 l_2 = +29; end
		6037: begin l_1 = -26;
				 l_2 = -29; end
		11346: begin l_1 = +26;
				 l_2 = +30; end
		16266: begin l_1 = +26;
				 l_2 = -30; end
		2347: begin l_1 = -26;
				 l_2 = +30; end
		7267: begin l_1 = -26;
				 l_2 = -30; end
		8886: begin l_1 = +26;
				 l_2 = +31; end
		113: begin l_1 = +26;
				 l_2 = -31; end
		18500: begin l_1 = -26;
				 l_2 = +31; end
		9727: begin l_1 = -26;
				 l_2 = -31; end
		3966: begin l_1 = +26;
				 l_2 = +32; end
		5033: begin l_1 = +26;
				 l_2 = -32; end
		13580: begin l_1 = -26;
				 l_2 = +32; end
		14647: begin l_1 = -26;
				 l_2 = -32; end
		12739: begin l_1 = +26;
				 l_2 = +33; end
		14873: begin l_1 = +26;
				 l_2 = -33; end
		3740: begin l_1 = -26;
				 l_2 = +33; end
		5874: begin l_1 = -26;
				 l_2 = -33; end
		11672: begin l_1 = +26;
				 l_2 = +34; end
		15940: begin l_1 = +26;
				 l_2 = -34; end
		2673: begin l_1 = -26;
				 l_2 = +34; end
		6941: begin l_1 = -26;
				 l_2 = -34; end
		9538: begin l_1 = +26;
				 l_2 = +35; end
		18074: begin l_1 = +26;
				 l_2 = -35; end
		539: begin l_1 = -26;
				 l_2 = +35; end
		9075: begin l_1 = -26;
				 l_2 = -35; end
		5270: begin l_1 = +26;
				 l_2 = +36; end
		3729: begin l_1 = +26;
				 l_2 = -36; end
		14884: begin l_1 = -26;
				 l_2 = +36; end
		13343: begin l_1 = -26;
				 l_2 = -36; end
		15347: begin l_1 = +26;
				 l_2 = +37; end
		12265: begin l_1 = +26;
				 l_2 = -37; end
		6348: begin l_1 = -26;
				 l_2 = +37; end
		3266: begin l_1 = -26;
				 l_2 = -37; end
		16888: begin l_1 = +26;
				 l_2 = +38; end
		10724: begin l_1 = +26;
				 l_2 = -38; end
		7889: begin l_1 = -26;
				 l_2 = +38; end
		1725: begin l_1 = -26;
				 l_2 = -38; end
		1357: begin l_1 = +26;
				 l_2 = +39; end
		7642: begin l_1 = +26;
				 l_2 = -39; end
		10971: begin l_1 = -26;
				 l_2 = +39; end
		17256: begin l_1 = -26;
				 l_2 = -39; end
		7521: begin l_1 = +26;
				 l_2 = +40; end
		1478: begin l_1 = +26;
				 l_2 = -40; end
		17135: begin l_1 = -26;
				 l_2 = +40; end
		11092: begin l_1 = -26;
				 l_2 = -40; end
		1236: begin l_1 = +26;
				 l_2 = +41; end
		7763: begin l_1 = +26;
				 l_2 = -41; end
		10850: begin l_1 = -26;
				 l_2 = +41; end
		17377: begin l_1 = -26;
				 l_2 = -41; end
		7279: begin l_1 = +26;
				 l_2 = +42; end
		1720: begin l_1 = +26;
				 l_2 = -42; end
		16893: begin l_1 = -26;
				 l_2 = +42; end
		11334: begin l_1 = -26;
				 l_2 = -42; end
		752: begin l_1 = +26;
				 l_2 = +43; end
		8247: begin l_1 = +26;
				 l_2 = -43; end
		10366: begin l_1 = -26;
				 l_2 = +43; end
		17861: begin l_1 = -26;
				 l_2 = -43; end
		6311: begin l_1 = +26;
				 l_2 = +44; end
		2688: begin l_1 = +26;
				 l_2 = -44; end
		15925: begin l_1 = -26;
				 l_2 = +44; end
		12302: begin l_1 = -26;
				 l_2 = -44; end
		17429: begin l_1 = +26;
				 l_2 = +45; end
		10183: begin l_1 = +26;
				 l_2 = -45; end
		8430: begin l_1 = -26;
				 l_2 = +45; end
		1184: begin l_1 = -26;
				 l_2 = -45; end
		8384: begin l_1 = -27;
				 l_2 = +29; end
		10229: begin l_1 = -27;
				 l_2 = -28; end
		7769: begin l_1 = +27;
				 l_2 = +29; end
		10844: begin l_1 = -27;
				 l_2 = -29; end
		6539: begin l_1 = +27;
				 l_2 = +30; end
		11459: begin l_1 = +27;
				 l_2 = -30; end
		7154: begin l_1 = -27;
				 l_2 = +30; end
		12074: begin l_1 = -27;
				 l_2 = -30; end
		4079: begin l_1 = +27;
				 l_2 = +31; end
		13919: begin l_1 = +27;
				 l_2 = -31; end
		4694: begin l_1 = -27;
				 l_2 = +31; end
		14534: begin l_1 = -27;
				 l_2 = -31; end
		17772: begin l_1 = +27;
				 l_2 = +32; end
		226: begin l_1 = +27;
				 l_2 = -32; end
		18387: begin l_1 = -27;
				 l_2 = +32; end
		841: begin l_1 = -27;
				 l_2 = -32; end
		7932: begin l_1 = +27;
				 l_2 = +33; end
		10066: begin l_1 = +27;
				 l_2 = -33; end
		8547: begin l_1 = -27;
				 l_2 = +33; end
		10681: begin l_1 = -27;
				 l_2 = -33; end
		6865: begin l_1 = +27;
				 l_2 = +34; end
		11133: begin l_1 = +27;
				 l_2 = -34; end
		7480: begin l_1 = -27;
				 l_2 = +34; end
		11748: begin l_1 = -27;
				 l_2 = -34; end
		4731: begin l_1 = +27;
				 l_2 = +35; end
		13267: begin l_1 = +27;
				 l_2 = -35; end
		5346: begin l_1 = -27;
				 l_2 = +35; end
		13882: begin l_1 = -27;
				 l_2 = -35; end
		463: begin l_1 = +27;
				 l_2 = +36; end
		17535: begin l_1 = +27;
				 l_2 = -36; end
		1078: begin l_1 = -27;
				 l_2 = +36; end
		18150: begin l_1 = -27;
				 l_2 = -36; end
		10540: begin l_1 = +27;
				 l_2 = +37; end
		7458: begin l_1 = +27;
				 l_2 = -37; end
		11155: begin l_1 = -27;
				 l_2 = +37; end
		8073: begin l_1 = -27;
				 l_2 = -37; end
		12081: begin l_1 = +27;
				 l_2 = +38; end
		5917: begin l_1 = +27;
				 l_2 = -38; end
		12696: begin l_1 = -27;
				 l_2 = +38; end
		6532: begin l_1 = -27;
				 l_2 = -38; end
		15163: begin l_1 = +27;
				 l_2 = +39; end
		2835: begin l_1 = +27;
				 l_2 = -39; end
		15778: begin l_1 = -27;
				 l_2 = +39; end
		3450: begin l_1 = -27;
				 l_2 = -39; end
		2714: begin l_1 = +27;
				 l_2 = +40; end
		15284: begin l_1 = +27;
				 l_2 = -40; end
		3329: begin l_1 = -27;
				 l_2 = +40; end
		15899: begin l_1 = -27;
				 l_2 = -40; end
		15042: begin l_1 = +27;
				 l_2 = +41; end
		2956: begin l_1 = +27;
				 l_2 = -41; end
		15657: begin l_1 = -27;
				 l_2 = +41; end
		3571: begin l_1 = -27;
				 l_2 = -41; end
		2472: begin l_1 = +27;
				 l_2 = +42; end
		15526: begin l_1 = +27;
				 l_2 = -42; end
		3087: begin l_1 = -27;
				 l_2 = +42; end
		16141: begin l_1 = -27;
				 l_2 = -42; end
		14558: begin l_1 = +27;
				 l_2 = +43; end
		3440: begin l_1 = +27;
				 l_2 = -43; end
		15173: begin l_1 = -27;
				 l_2 = +43; end
		4055: begin l_1 = -27;
				 l_2 = -43; end
		1504: begin l_1 = +27;
				 l_2 = +44; end
		16494: begin l_1 = +27;
				 l_2 = -44; end
		2119: begin l_1 = -27;
				 l_2 = +44; end
		17109: begin l_1 = -27;
				 l_2 = -44; end
		12622: begin l_1 = +27;
				 l_2 = +45; end
		5376: begin l_1 = +27;
				 l_2 = -45; end
		13237: begin l_1 = -27;
				 l_2 = +45; end
		5991: begin l_1 = -27;
				 l_2 = -45; end
		16768: begin l_1 = -28;
				 l_2 = +30; end
		1845: begin l_1 = -28;
				 l_2 = -29; end
		15538: begin l_1 = +28;
				 l_2 = +30; end
		3075: begin l_1 = -28;
				 l_2 = -30; end
		13078: begin l_1 = +28;
				 l_2 = +31; end
		4305: begin l_1 = +28;
				 l_2 = -31; end
		14308: begin l_1 = -28;
				 l_2 = +31; end
		5535: begin l_1 = -28;
				 l_2 = -31; end
		8158: begin l_1 = +28;
				 l_2 = +32; end
		9225: begin l_1 = +28;
				 l_2 = -32; end
		9388: begin l_1 = -28;
				 l_2 = +32; end
		10455: begin l_1 = -28;
				 l_2 = -32; end
		16931: begin l_1 = +28;
				 l_2 = +33; end
		452: begin l_1 = +28;
				 l_2 = -33; end
		18161: begin l_1 = -28;
				 l_2 = +33; end
		1682: begin l_1 = -28;
				 l_2 = -33; end
		15864: begin l_1 = +28;
				 l_2 = +34; end
		1519: begin l_1 = +28;
				 l_2 = -34; end
		17094: begin l_1 = -28;
				 l_2 = +34; end
		2749: begin l_1 = -28;
				 l_2 = -34; end
		13730: begin l_1 = +28;
				 l_2 = +35; end
		3653: begin l_1 = +28;
				 l_2 = -35; end
		14960: begin l_1 = -28;
				 l_2 = +35; end
		4883: begin l_1 = -28;
				 l_2 = -35; end
		9462: begin l_1 = +28;
				 l_2 = +36; end
		7921: begin l_1 = +28;
				 l_2 = -36; end
		10692: begin l_1 = -28;
				 l_2 = +36; end
		9151: begin l_1 = -28;
				 l_2 = -36; end
		926: begin l_1 = +28;
				 l_2 = +37; end
		16457: begin l_1 = +28;
				 l_2 = -37; end
		2156: begin l_1 = -28;
				 l_2 = +37; end
		17687: begin l_1 = -28;
				 l_2 = -37; end
		2467: begin l_1 = +28;
				 l_2 = +38; end
		14916: begin l_1 = +28;
				 l_2 = -38; end
		3697: begin l_1 = -28;
				 l_2 = +38; end
		16146: begin l_1 = -28;
				 l_2 = -38; end
		5549: begin l_1 = +28;
				 l_2 = +39; end
		11834: begin l_1 = +28;
				 l_2 = -39; end
		6779: begin l_1 = -28;
				 l_2 = +39; end
		13064: begin l_1 = -28;
				 l_2 = -39; end
		11713: begin l_1 = +28;
				 l_2 = +40; end
		5670: begin l_1 = +28;
				 l_2 = -40; end
		12943: begin l_1 = -28;
				 l_2 = +40; end
		6900: begin l_1 = -28;
				 l_2 = -40; end
		5428: begin l_1 = +28;
				 l_2 = +41; end
		11955: begin l_1 = +28;
				 l_2 = -41; end
		6658: begin l_1 = -28;
				 l_2 = +41; end
		13185: begin l_1 = -28;
				 l_2 = -41; end
		11471: begin l_1 = +28;
				 l_2 = +42; end
		5912: begin l_1 = +28;
				 l_2 = -42; end
		12701: begin l_1 = -28;
				 l_2 = +42; end
		7142: begin l_1 = -28;
				 l_2 = -42; end
		4944: begin l_1 = +28;
				 l_2 = +43; end
		12439: begin l_1 = +28;
				 l_2 = -43; end
		6174: begin l_1 = -28;
				 l_2 = +43; end
		13669: begin l_1 = -28;
				 l_2 = -43; end
		10503: begin l_1 = +28;
				 l_2 = +44; end
		6880: begin l_1 = +28;
				 l_2 = -44; end
		11733: begin l_1 = -28;
				 l_2 = +44; end
		8110: begin l_1 = -28;
				 l_2 = -44; end
		3008: begin l_1 = +28;
				 l_2 = +45; end
		14375: begin l_1 = +28;
				 l_2 = -45; end
		4238: begin l_1 = -28;
				 l_2 = +45; end
		15605: begin l_1 = -28;
				 l_2 = -45; end
		14923: begin l_1 = -29;
				 l_2 = +31; end
		3690: begin l_1 = -29;
				 l_2 = -30; end
		12463: begin l_1 = +29;
				 l_2 = +31; end
		6150: begin l_1 = -29;
				 l_2 = -31; end
		7543: begin l_1 = +29;
				 l_2 = +32; end
		8610: begin l_1 = +29;
				 l_2 = -32; end
		10003: begin l_1 = -29;
				 l_2 = +32; end
		11070: begin l_1 = -29;
				 l_2 = -32; end
		16316: begin l_1 = +29;
				 l_2 = +33; end
		18450: begin l_1 = +29;
				 l_2 = -33; end
		163: begin l_1 = -29;
				 l_2 = +33; end
		2297: begin l_1 = -29;
				 l_2 = -33; end
		15249: begin l_1 = +29;
				 l_2 = +34; end
		904: begin l_1 = +29;
				 l_2 = -34; end
		17709: begin l_1 = -29;
				 l_2 = +34; end
		3364: begin l_1 = -29;
				 l_2 = -34; end
		13115: begin l_1 = +29;
				 l_2 = +35; end
		3038: begin l_1 = +29;
				 l_2 = -35; end
		15575: begin l_1 = -29;
				 l_2 = +35; end
		5498: begin l_1 = -29;
				 l_2 = -35; end
		8847: begin l_1 = +29;
				 l_2 = +36; end
		7306: begin l_1 = +29;
				 l_2 = -36; end
		11307: begin l_1 = -29;
				 l_2 = +36; end
		9766: begin l_1 = -29;
				 l_2 = -36; end
		311: begin l_1 = +29;
				 l_2 = +37; end
		15842: begin l_1 = +29;
				 l_2 = -37; end
		2771: begin l_1 = -29;
				 l_2 = +37; end
		18302: begin l_1 = -29;
				 l_2 = -37; end
		1852: begin l_1 = +29;
				 l_2 = +38; end
		14301: begin l_1 = +29;
				 l_2 = -38; end
		4312: begin l_1 = -29;
				 l_2 = +38; end
		16761: begin l_1 = -29;
				 l_2 = -38; end
		4934: begin l_1 = +29;
				 l_2 = +39; end
		11219: begin l_1 = +29;
				 l_2 = -39; end
		7394: begin l_1 = -29;
				 l_2 = +39; end
		13679: begin l_1 = -29;
				 l_2 = -39; end
		11098: begin l_1 = +29;
				 l_2 = +40; end
		5055: begin l_1 = +29;
				 l_2 = -40; end
		13558: begin l_1 = -29;
				 l_2 = +40; end
		7515: begin l_1 = -29;
				 l_2 = -40; end
		4813: begin l_1 = +29;
				 l_2 = +41; end
		11340: begin l_1 = +29;
				 l_2 = -41; end
		7273: begin l_1 = -29;
				 l_2 = +41; end
		13800: begin l_1 = -29;
				 l_2 = -41; end
		10856: begin l_1 = +29;
				 l_2 = +42; end
		5297: begin l_1 = +29;
				 l_2 = -42; end
		13316: begin l_1 = -29;
				 l_2 = +42; end
		7757: begin l_1 = -29;
				 l_2 = -42; end
		4329: begin l_1 = +29;
				 l_2 = +43; end
		11824: begin l_1 = +29;
				 l_2 = -43; end
		6789: begin l_1 = -29;
				 l_2 = +43; end
		14284: begin l_1 = -29;
				 l_2 = -43; end
		9888: begin l_1 = +29;
				 l_2 = +44; end
		6265: begin l_1 = +29;
				 l_2 = -44; end
		12348: begin l_1 = -29;
				 l_2 = +44; end
		8725: begin l_1 = -29;
				 l_2 = -44; end
		2393: begin l_1 = +29;
				 l_2 = +45; end
		13760: begin l_1 = +29;
				 l_2 = -45; end
		4853: begin l_1 = -29;
				 l_2 = +45; end
		16220: begin l_1 = -29;
				 l_2 = -45; end
		11233: begin l_1 = -30;
				 l_2 = +32; end
		7380: begin l_1 = -30;
				 l_2 = -31; end
		6313: begin l_1 = +30;
				 l_2 = +32; end
		12300: begin l_1 = -30;
				 l_2 = -32; end
		15086: begin l_1 = +30;
				 l_2 = +33; end
		17220: begin l_1 = +30;
				 l_2 = -33; end
		1393: begin l_1 = -30;
				 l_2 = +33; end
		3527: begin l_1 = -30;
				 l_2 = -33; end
		14019: begin l_1 = +30;
				 l_2 = +34; end
		18287: begin l_1 = +30;
				 l_2 = -34; end
		326: begin l_1 = -30;
				 l_2 = +34; end
		4594: begin l_1 = -30;
				 l_2 = -34; end
		11885: begin l_1 = +30;
				 l_2 = +35; end
		1808: begin l_1 = +30;
				 l_2 = -35; end
		16805: begin l_1 = -30;
				 l_2 = +35; end
		6728: begin l_1 = -30;
				 l_2 = -35; end
		7617: begin l_1 = +30;
				 l_2 = +36; end
		6076: begin l_1 = +30;
				 l_2 = -36; end
		12537: begin l_1 = -30;
				 l_2 = +36; end
		10996: begin l_1 = -30;
				 l_2 = -36; end
		17694: begin l_1 = +30;
				 l_2 = +37; end
		14612: begin l_1 = +30;
				 l_2 = -37; end
		4001: begin l_1 = -30;
				 l_2 = +37; end
		919: begin l_1 = -30;
				 l_2 = -37; end
		622: begin l_1 = +30;
				 l_2 = +38; end
		13071: begin l_1 = +30;
				 l_2 = -38; end
		5542: begin l_1 = -30;
				 l_2 = +38; end
		17991: begin l_1 = -30;
				 l_2 = -38; end
		3704: begin l_1 = +30;
				 l_2 = +39; end
		9989: begin l_1 = +30;
				 l_2 = -39; end
		8624: begin l_1 = -30;
				 l_2 = +39; end
		14909: begin l_1 = -30;
				 l_2 = -39; end
		9868: begin l_1 = +30;
				 l_2 = +40; end
		3825: begin l_1 = +30;
				 l_2 = -40; end
		14788: begin l_1 = -30;
				 l_2 = +40; end
		8745: begin l_1 = -30;
				 l_2 = -40; end
		3583: begin l_1 = +30;
				 l_2 = +41; end
		10110: begin l_1 = +30;
				 l_2 = -41; end
		8503: begin l_1 = -30;
				 l_2 = +41; end
		15030: begin l_1 = -30;
				 l_2 = -41; end
		9626: begin l_1 = +30;
				 l_2 = +42; end
		4067: begin l_1 = +30;
				 l_2 = -42; end
		14546: begin l_1 = -30;
				 l_2 = +42; end
		8987: begin l_1 = -30;
				 l_2 = -42; end
		3099: begin l_1 = +30;
				 l_2 = +43; end
		10594: begin l_1 = +30;
				 l_2 = -43; end
		8019: begin l_1 = -30;
				 l_2 = +43; end
		15514: begin l_1 = -30;
				 l_2 = -43; end
		8658: begin l_1 = +30;
				 l_2 = +44; end
		5035: begin l_1 = +30;
				 l_2 = -44; end
		13578: begin l_1 = -30;
				 l_2 = +44; end
		9955: begin l_1 = -30;
				 l_2 = -44; end
		1163: begin l_1 = +30;
				 l_2 = +45; end
		12530: begin l_1 = +30;
				 l_2 = -45; end
		6083: begin l_1 = -30;
				 l_2 = +45; end
		17450: begin l_1 = -30;
				 l_2 = -45; end
		3853: begin l_1 = -31;
				 l_2 = +33; end
		14760: begin l_1 = -31;
				 l_2 = -32; end
		12626: begin l_1 = +31;
				 l_2 = +33; end
		5987: begin l_1 = -31;
				 l_2 = -33; end
		11559: begin l_1 = +31;
				 l_2 = +34; end
		15827: begin l_1 = +31;
				 l_2 = -34; end
		2786: begin l_1 = -31;
				 l_2 = +34; end
		7054: begin l_1 = -31;
				 l_2 = -34; end
		9425: begin l_1 = +31;
				 l_2 = +35; end
		17961: begin l_1 = +31;
				 l_2 = -35; end
		652: begin l_1 = -31;
				 l_2 = +35; end
		9188: begin l_1 = -31;
				 l_2 = -35; end
		5157: begin l_1 = +31;
				 l_2 = +36; end
		3616: begin l_1 = +31;
				 l_2 = -36; end
		14997: begin l_1 = -31;
				 l_2 = +36; end
		13456: begin l_1 = -31;
				 l_2 = -36; end
		15234: begin l_1 = +31;
				 l_2 = +37; end
		12152: begin l_1 = +31;
				 l_2 = -37; end
		6461: begin l_1 = -31;
				 l_2 = +37; end
		3379: begin l_1 = -31;
				 l_2 = -37; end
		16775: begin l_1 = +31;
				 l_2 = +38; end
		10611: begin l_1 = +31;
				 l_2 = -38; end
		8002: begin l_1 = -31;
				 l_2 = +38; end
		1838: begin l_1 = -31;
				 l_2 = -38; end
		1244: begin l_1 = +31;
				 l_2 = +39; end
		7529: begin l_1 = +31;
				 l_2 = -39; end
		11084: begin l_1 = -31;
				 l_2 = +39; end
		17369: begin l_1 = -31;
				 l_2 = -39; end
		7408: begin l_1 = +31;
				 l_2 = +40; end
		1365: begin l_1 = +31;
				 l_2 = -40; end
		17248: begin l_1 = -31;
				 l_2 = +40; end
		11205: begin l_1 = -31;
				 l_2 = -40; end
		1123: begin l_1 = +31;
				 l_2 = +41; end
		7650: begin l_1 = +31;
				 l_2 = -41; end
		10963: begin l_1 = -31;
				 l_2 = +41; end
		17490: begin l_1 = -31;
				 l_2 = -41; end
		7166: begin l_1 = +31;
				 l_2 = +42; end
		1607: begin l_1 = +31;
				 l_2 = -42; end
		17006: begin l_1 = -31;
				 l_2 = +42; end
		11447: begin l_1 = -31;
				 l_2 = -42; end
		639: begin l_1 = +31;
				 l_2 = +43; end
		8134: begin l_1 = +31;
				 l_2 = -43; end
		10479: begin l_1 = -31;
				 l_2 = +43; end
		17974: begin l_1 = -31;
				 l_2 = -43; end
		6198: begin l_1 = +31;
				 l_2 = +44; end
		2575: begin l_1 = +31;
				 l_2 = -44; end
		16038: begin l_1 = -31;
				 l_2 = +44; end
		12415: begin l_1 = -31;
				 l_2 = -44; end
		17316: begin l_1 = +31;
				 l_2 = +45; end
		10070: begin l_1 = +31;
				 l_2 = -45; end
		8543: begin l_1 = -31;
				 l_2 = +45; end
		1297: begin l_1 = -31;
				 l_2 = -45; end
		7706: begin l_1 = -32;
				 l_2 = +34; end
		10907: begin l_1 = -32;
				 l_2 = -33; end
		6639: begin l_1 = +32;
				 l_2 = +34; end
		11974: begin l_1 = -32;
				 l_2 = -34; end
		4505: begin l_1 = +32;
				 l_2 = +35; end
		13041: begin l_1 = +32;
				 l_2 = -35; end
		5572: begin l_1 = -32;
				 l_2 = +35; end
		14108: begin l_1 = -32;
				 l_2 = -35; end
		237: begin l_1 = +32;
				 l_2 = +36; end
		17309: begin l_1 = +32;
				 l_2 = -36; end
		1304: begin l_1 = -32;
				 l_2 = +36; end
		18376: begin l_1 = -32;
				 l_2 = -36; end
		10314: begin l_1 = +32;
				 l_2 = +37; end
		7232: begin l_1 = +32;
				 l_2 = -37; end
		11381: begin l_1 = -32;
				 l_2 = +37; end
		8299: begin l_1 = -32;
				 l_2 = -37; end
		11855: begin l_1 = +32;
				 l_2 = +38; end
		5691: begin l_1 = +32;
				 l_2 = -38; end
		12922: begin l_1 = -32;
				 l_2 = +38; end
		6758: begin l_1 = -32;
				 l_2 = -38; end
		14937: begin l_1 = +32;
				 l_2 = +39; end
		2609: begin l_1 = +32;
				 l_2 = -39; end
		16004: begin l_1 = -32;
				 l_2 = +39; end
		3676: begin l_1 = -32;
				 l_2 = -39; end
		2488: begin l_1 = +32;
				 l_2 = +40; end
		15058: begin l_1 = +32;
				 l_2 = -40; end
		3555: begin l_1 = -32;
				 l_2 = +40; end
		16125: begin l_1 = -32;
				 l_2 = -40; end
		14816: begin l_1 = +32;
				 l_2 = +41; end
		2730: begin l_1 = +32;
				 l_2 = -41; end
		15883: begin l_1 = -32;
				 l_2 = +41; end
		3797: begin l_1 = -32;
				 l_2 = -41; end
		2246: begin l_1 = +32;
				 l_2 = +42; end
		15300: begin l_1 = +32;
				 l_2 = -42; end
		3313: begin l_1 = -32;
				 l_2 = +42; end
		16367: begin l_1 = -32;
				 l_2 = -42; end
		14332: begin l_1 = +32;
				 l_2 = +43; end
		3214: begin l_1 = +32;
				 l_2 = -43; end
		15399: begin l_1 = -32;
				 l_2 = +43; end
		4281: begin l_1 = -32;
				 l_2 = -43; end
		1278: begin l_1 = +32;
				 l_2 = +44; end
		16268: begin l_1 = +32;
				 l_2 = -44; end
		2345: begin l_1 = -32;
				 l_2 = +44; end
		17335: begin l_1 = -32;
				 l_2 = -44; end
		12396: begin l_1 = +32;
				 l_2 = +45; end
		5150: begin l_1 = +32;
				 l_2 = -45; end
		13463: begin l_1 = -32;
				 l_2 = +45; end
		6217: begin l_1 = -32;
				 l_2 = -45; end
		15412: begin l_1 = -33;
				 l_2 = +35; end
		3201: begin l_1 = -33;
				 l_2 = -34; end
		13278: begin l_1 = +33;
				 l_2 = +35; end
		5335: begin l_1 = -33;
				 l_2 = -35; end
		9010: begin l_1 = +33;
				 l_2 = +36; end
		7469: begin l_1 = +33;
				 l_2 = -36; end
		11144: begin l_1 = -33;
				 l_2 = +36; end
		9603: begin l_1 = -33;
				 l_2 = -36; end
		474: begin l_1 = +33;
				 l_2 = +37; end
		16005: begin l_1 = +33;
				 l_2 = -37; end
		2608: begin l_1 = -33;
				 l_2 = +37; end
		18139: begin l_1 = -33;
				 l_2 = -37; end
		2015: begin l_1 = +33;
				 l_2 = +38; end
		14464: begin l_1 = +33;
				 l_2 = -38; end
		4149: begin l_1 = -33;
				 l_2 = +38; end
		16598: begin l_1 = -33;
				 l_2 = -38; end
		5097: begin l_1 = +33;
				 l_2 = +39; end
		11382: begin l_1 = +33;
				 l_2 = -39; end
		7231: begin l_1 = -33;
				 l_2 = +39; end
		13516: begin l_1 = -33;
				 l_2 = -39; end
		11261: begin l_1 = +33;
				 l_2 = +40; end
		5218: begin l_1 = +33;
				 l_2 = -40; end
		13395: begin l_1 = -33;
				 l_2 = +40; end
		7352: begin l_1 = -33;
				 l_2 = -40; end
		4976: begin l_1 = +33;
				 l_2 = +41; end
		11503: begin l_1 = +33;
				 l_2 = -41; end
		7110: begin l_1 = -33;
				 l_2 = +41; end
		13637: begin l_1 = -33;
				 l_2 = -41; end
		11019: begin l_1 = +33;
				 l_2 = +42; end
		5460: begin l_1 = +33;
				 l_2 = -42; end
		13153: begin l_1 = -33;
				 l_2 = +42; end
		7594: begin l_1 = -33;
				 l_2 = -42; end
		4492: begin l_1 = +33;
				 l_2 = +43; end
		11987: begin l_1 = +33;
				 l_2 = -43; end
		6626: begin l_1 = -33;
				 l_2 = +43; end
		14121: begin l_1 = -33;
				 l_2 = -43; end
		10051: begin l_1 = +33;
				 l_2 = +44; end
		6428: begin l_1 = +33;
				 l_2 = -44; end
		12185: begin l_1 = -33;
				 l_2 = +44; end
		8562: begin l_1 = -33;
				 l_2 = -44; end
		2556: begin l_1 = +33;
				 l_2 = +45; end
		13923: begin l_1 = +33;
				 l_2 = -45; end
		4690: begin l_1 = -33;
				 l_2 = +45; end
		16057: begin l_1 = -33;
				 l_2 = -45; end
		12211: begin l_1 = -34;
				 l_2 = +36; end
		6402: begin l_1 = -34;
				 l_2 = -35; end
		7943: begin l_1 = +34;
				 l_2 = +36; end
		10670: begin l_1 = -34;
				 l_2 = -36; end
		18020: begin l_1 = +34;
				 l_2 = +37; end
		14938: begin l_1 = +34;
				 l_2 = -37; end
		3675: begin l_1 = -34;
				 l_2 = +37; end
		593: begin l_1 = -34;
				 l_2 = -37; end
		948: begin l_1 = +34;
				 l_2 = +38; end
		13397: begin l_1 = +34;
				 l_2 = -38; end
		5216: begin l_1 = -34;
				 l_2 = +38; end
		17665: begin l_1 = -34;
				 l_2 = -38; end
		4030: begin l_1 = +34;
				 l_2 = +39; end
		10315: begin l_1 = +34;
				 l_2 = -39; end
		8298: begin l_1 = -34;
				 l_2 = +39; end
		14583: begin l_1 = -34;
				 l_2 = -39; end
		10194: begin l_1 = +34;
				 l_2 = +40; end
		4151: begin l_1 = +34;
				 l_2 = -40; end
		14462: begin l_1 = -34;
				 l_2 = +40; end
		8419: begin l_1 = -34;
				 l_2 = -40; end
		3909: begin l_1 = +34;
				 l_2 = +41; end
		10436: begin l_1 = +34;
				 l_2 = -41; end
		8177: begin l_1 = -34;
				 l_2 = +41; end
		14704: begin l_1 = -34;
				 l_2 = -41; end
		9952: begin l_1 = +34;
				 l_2 = +42; end
		4393: begin l_1 = +34;
				 l_2 = -42; end
		14220: begin l_1 = -34;
				 l_2 = +42; end
		8661: begin l_1 = -34;
				 l_2 = -42; end
		3425: begin l_1 = +34;
				 l_2 = +43; end
		10920: begin l_1 = +34;
				 l_2 = -43; end
		7693: begin l_1 = -34;
				 l_2 = +43; end
		15188: begin l_1 = -34;
				 l_2 = -43; end
		8984: begin l_1 = +34;
				 l_2 = +44; end
		5361: begin l_1 = +34;
				 l_2 = -44; end
		13252: begin l_1 = -34;
				 l_2 = +44; end
		9629: begin l_1 = -34;
				 l_2 = -44; end
		1489: begin l_1 = +34;
				 l_2 = +45; end
		12856: begin l_1 = +34;
				 l_2 = -45; end
		5757: begin l_1 = -34;
				 l_2 = +45; end
		17124: begin l_1 = -34;
				 l_2 = -45; end
		5809: begin l_1 = -35;
				 l_2 = +37; end
		12804: begin l_1 = -35;
				 l_2 = -36; end
		15886: begin l_1 = +35;
				 l_2 = +37; end
		2727: begin l_1 = -35;
				 l_2 = -37; end
		17427: begin l_1 = +35;
				 l_2 = +38; end
		11263: begin l_1 = +35;
				 l_2 = -38; end
		7350: begin l_1 = -35;
				 l_2 = +38; end
		1186: begin l_1 = -35;
				 l_2 = -38; end
		1896: begin l_1 = +35;
				 l_2 = +39; end
		8181: begin l_1 = +35;
				 l_2 = -39; end
		10432: begin l_1 = -35;
				 l_2 = +39; end
		16717: begin l_1 = -35;
				 l_2 = -39; end
		8060: begin l_1 = +35;
				 l_2 = +40; end
		2017: begin l_1 = +35;
				 l_2 = -40; end
		16596: begin l_1 = -35;
				 l_2 = +40; end
		10553: begin l_1 = -35;
				 l_2 = -40; end
		1775: begin l_1 = +35;
				 l_2 = +41; end
		8302: begin l_1 = +35;
				 l_2 = -41; end
		10311: begin l_1 = -35;
				 l_2 = +41; end
		16838: begin l_1 = -35;
				 l_2 = -41; end
		7818: begin l_1 = +35;
				 l_2 = +42; end
		2259: begin l_1 = +35;
				 l_2 = -42; end
		16354: begin l_1 = -35;
				 l_2 = +42; end
		10795: begin l_1 = -35;
				 l_2 = -42; end
		1291: begin l_1 = +35;
				 l_2 = +43; end
		8786: begin l_1 = +35;
				 l_2 = -43; end
		9827: begin l_1 = -35;
				 l_2 = +43; end
		17322: begin l_1 = -35;
				 l_2 = -43; end
		6850: begin l_1 = +35;
				 l_2 = +44; end
		3227: begin l_1 = +35;
				 l_2 = -44; end
		15386: begin l_1 = -35;
				 l_2 = +44; end
		11763: begin l_1 = -35;
				 l_2 = -44; end
		17968: begin l_1 = +35;
				 l_2 = +45; end
		10722: begin l_1 = +35;
				 l_2 = -45; end
		7891: begin l_1 = -35;
				 l_2 = +45; end
		645: begin l_1 = -35;
				 l_2 = -45; end
		11618: begin l_1 = -36;
				 l_2 = +38; end
		6995: begin l_1 = -36;
				 l_2 = -37; end
		13159: begin l_1 = +36;
				 l_2 = +38; end
		5454: begin l_1 = -36;
				 l_2 = -38; end
		16241: begin l_1 = +36;
				 l_2 = +39; end
		3913: begin l_1 = +36;
				 l_2 = -39; end
		14700: begin l_1 = -36;
				 l_2 = +39; end
		2372: begin l_1 = -36;
				 l_2 = -39; end
		3792: begin l_1 = +36;
				 l_2 = +40; end
		16362: begin l_1 = +36;
				 l_2 = -40; end
		2251: begin l_1 = -36;
				 l_2 = +40; end
		14821: begin l_1 = -36;
				 l_2 = -40; end
		16120: begin l_1 = +36;
				 l_2 = +41; end
		4034: begin l_1 = +36;
				 l_2 = -41; end
		14579: begin l_1 = -36;
				 l_2 = +41; end
		2493: begin l_1 = -36;
				 l_2 = -41; end
		3550: begin l_1 = +36;
				 l_2 = +42; end
		16604: begin l_1 = +36;
				 l_2 = -42; end
		2009: begin l_1 = -36;
				 l_2 = +42; end
		15063: begin l_1 = -36;
				 l_2 = -42; end
		15636: begin l_1 = +36;
				 l_2 = +43; end
		4518: begin l_1 = +36;
				 l_2 = -43; end
		14095: begin l_1 = -36;
				 l_2 = +43; end
		2977: begin l_1 = -36;
				 l_2 = -43; end
		2582: begin l_1 = +36;
				 l_2 = +44; end
		17572: begin l_1 = +36;
				 l_2 = -44; end
		1041: begin l_1 = -36;
				 l_2 = +44; end
		16031: begin l_1 = -36;
				 l_2 = -44; end
		13700: begin l_1 = +36;
				 l_2 = +45; end
		6454: begin l_1 = +36;
				 l_2 = -45; end
		12159: begin l_1 = -36;
				 l_2 = +45; end
		4913: begin l_1 = -36;
				 l_2 = -45; end
		4623: begin l_1 = -37;
				 l_2 = +39; end
		13990: begin l_1 = -37;
				 l_2 = -38; end
		7705: begin l_1 = +37;
				 l_2 = +39; end
		10908: begin l_1 = -37;
				 l_2 = -39; end
		13869: begin l_1 = +37;
				 l_2 = +40; end
		7826: begin l_1 = +37;
				 l_2 = -40; end
		10787: begin l_1 = -37;
				 l_2 = +40; end
		4744: begin l_1 = -37;
				 l_2 = -40; end
		7584: begin l_1 = +37;
				 l_2 = +41; end
		14111: begin l_1 = +37;
				 l_2 = -41; end
		4502: begin l_1 = -37;
				 l_2 = +41; end
		11029: begin l_1 = -37;
				 l_2 = -41; end
		13627: begin l_1 = +37;
				 l_2 = +42; end
		8068: begin l_1 = +37;
				 l_2 = -42; end
		10545: begin l_1 = -37;
				 l_2 = +42; end
		4986: begin l_1 = -37;
				 l_2 = -42; end
		7100: begin l_1 = +37;
				 l_2 = +43; end
		14595: begin l_1 = +37;
				 l_2 = -43; end
		4018: begin l_1 = -37;
				 l_2 = +43; end
		11513: begin l_1 = -37;
				 l_2 = -43; end
		12659: begin l_1 = +37;
				 l_2 = +44; end
		9036: begin l_1 = +37;
				 l_2 = -44; end
		9577: begin l_1 = -37;
				 l_2 = +44; end
		5954: begin l_1 = -37;
				 l_2 = -44; end
		5164: begin l_1 = +37;
				 l_2 = +45; end
		16531: begin l_1 = +37;
				 l_2 = -45; end
		2082: begin l_1 = -37;
				 l_2 = +45; end
		13449: begin l_1 = -37;
				 l_2 = -45; end
		9246: begin l_1 = -38;
				 l_2 = +40; end
		9367: begin l_1 = -38;
				 l_2 = -39; end
		15410: begin l_1 = +38;
				 l_2 = +40; end
		3203: begin l_1 = -38;
				 l_2 = -40; end
		9125: begin l_1 = +38;
				 l_2 = +41; end
		15652: begin l_1 = +38;
				 l_2 = -41; end
		2961: begin l_1 = -38;
				 l_2 = +41; end
		9488: begin l_1 = -38;
				 l_2 = -41; end
		15168: begin l_1 = +38;
				 l_2 = +42; end
		9609: begin l_1 = +38;
				 l_2 = -42; end
		9004: begin l_1 = -38;
				 l_2 = +42; end
		3445: begin l_1 = -38;
				 l_2 = -42; end
		8641: begin l_1 = +38;
				 l_2 = +43; end
		16136: begin l_1 = +38;
				 l_2 = -43; end
		2477: begin l_1 = -38;
				 l_2 = +43; end
		9972: begin l_1 = -38;
				 l_2 = -43; end
		14200: begin l_1 = +38;
				 l_2 = +44; end
		10577: begin l_1 = +38;
				 l_2 = -44; end
		8036: begin l_1 = -38;
				 l_2 = +44; end
		4413: begin l_1 = -38;
				 l_2 = -44; end
		6705: begin l_1 = +38;
				 l_2 = +45; end
		18072: begin l_1 = +38;
				 l_2 = -45; end
		541: begin l_1 = -38;
				 l_2 = +45; end
		11908: begin l_1 = -38;
				 l_2 = -45; end
		18492: begin l_1 = -39;
				 l_2 = +41; end
		121: begin l_1 = -39;
				 l_2 = -40; end
		12207: begin l_1 = +39;
				 l_2 = +41; end
		6406: begin l_1 = -39;
				 l_2 = -41; end
		18250: begin l_1 = +39;
				 l_2 = +42; end
		12691: begin l_1 = +39;
				 l_2 = -42; end
		5922: begin l_1 = -39;
				 l_2 = +42; end
		363: begin l_1 = -39;
				 l_2 = -42; end
		11723: begin l_1 = +39;
				 l_2 = +43; end
		605: begin l_1 = +39;
				 l_2 = -43; end
		18008: begin l_1 = -39;
				 l_2 = +43; end
		6890: begin l_1 = -39;
				 l_2 = -43; end
		17282: begin l_1 = +39;
				 l_2 = +44; end
		13659: begin l_1 = +39;
				 l_2 = -44; end
		4954: begin l_1 = -39;
				 l_2 = +44; end
		1331: begin l_1 = -39;
				 l_2 = -44; end
		9787: begin l_1 = +39;
				 l_2 = +45; end
		2541: begin l_1 = +39;
				 l_2 = -45; end
		16072: begin l_1 = -39;
				 l_2 = +45; end
		8826: begin l_1 = -39;
				 l_2 = -45; end
		18371: begin l_1 = -40;
				 l_2 = +42; end
		242: begin l_1 = -40;
				 l_2 = -41; end
		5801: begin l_1 = +40;
				 l_2 = +42; end
		12812: begin l_1 = -40;
				 l_2 = -42; end
		17887: begin l_1 = +40;
				 l_2 = +43; end
		6769: begin l_1 = +40;
				 l_2 = -43; end
		11844: begin l_1 = -40;
				 l_2 = +43; end
		726: begin l_1 = -40;
				 l_2 = -43; end
		4833: begin l_1 = +40;
				 l_2 = +44; end
		1210: begin l_1 = +40;
				 l_2 = -44; end
		17403: begin l_1 = -40;
				 l_2 = +44; end
		13780: begin l_1 = -40;
				 l_2 = -44; end
		15951: begin l_1 = +40;
				 l_2 = +45; end
		8705: begin l_1 = +40;
				 l_2 = -45; end
		9908: begin l_1 = -40;
				 l_2 = +45; end
		2662: begin l_1 = -40;
				 l_2 = -45; end
		18129: begin l_1 = -41;
				 l_2 = +43; end
		484: begin l_1 = -41;
				 l_2 = -42; end
		11602: begin l_1 = +41;
				 l_2 = +43; end
		7011: begin l_1 = -41;
				 l_2 = -43; end
		17161: begin l_1 = +41;
				 l_2 = +44; end
		13538: begin l_1 = +41;
				 l_2 = -44; end
		5075: begin l_1 = -41;
				 l_2 = +44; end
		1452: begin l_1 = -41;
				 l_2 = -44; end
		9666: begin l_1 = +41;
				 l_2 = +45; end
		2420: begin l_1 = +41;
				 l_2 = -45; end
		16193: begin l_1 = -41;
				 l_2 = +45; end
		8947: begin l_1 = -41;
				 l_2 = -45; end
		17645: begin l_1 = -42;
				 l_2 = +44; end
		968: begin l_1 = -42;
				 l_2 = -43; end
		4591: begin l_1 = +42;
				 l_2 = +44; end
		14022: begin l_1 = -42;
				 l_2 = -44; end
		15709: begin l_1 = +42;
				 l_2 = +45; end
		8463: begin l_1 = +42;
				 l_2 = -45; end
		10150: begin l_1 = -42;
				 l_2 = +45; end
		2904: begin l_1 = -42;
				 l_2 = -45; end
		16677: begin l_1 = -43;
				 l_2 = +45; end
		1936: begin l_1 = -43;
				 l_2 = -44; end
		9182: begin l_1 = +43;
				 l_2 = +45; end
		9431: begin l_1 = -43;
				 l_2 = -45; end
		14741: begin l_1 = +44;
				 l_2 = +45; end
		3872: begin l_1 = -44;
				 l_2 = -45; end
		default: begin l_1 = 0;
					   l_2 = 0; end
	endcase
end

endmodule

// Product (AN) Code SEC_LUT_Decoder
// SEC_LUT_Decoder28bits.v
// Received codeword W = AN + e, e is single arithmetic weight error (AWE), +2^i or -2^i.
module SEC_LUT_Decoder28bits(W, N);
input 	[42:0]	W;
output	[27:0]	N;
parameter A = 17619;

wire 	[27:0]	Q;
wire 	[14:0]	R;
assign Q = W / A;
assign R = W - (A * Q);

reg	signed	[43:0]	Delta;
always@(*) begin
	case(R)
		1: Delta = 44'sb00000000000000000000000000000000000000000001;
		17618: Delta = 44'sb11111111111111111111111111111111111111111111;
		2: Delta = 44'sb00000000000000000000000000000000000000000010;
		17617: Delta = 44'sb11111111111111111111111111111111111111111110;
		4: Delta = 44'sb00000000000000000000000000000000000000000100;
		17615: Delta = 44'sb11111111111111111111111111111111111111111100;
		8: Delta = 44'sb00000000000000000000000000000000000000001000;
		17611: Delta = 44'sb11111111111111111111111111111111111111111000;
		16: Delta = 44'sb00000000000000000000000000000000000000010000;
		17603: Delta = 44'sb11111111111111111111111111111111111111110000;
		32: Delta = 44'sb00000000000000000000000000000000000000100000;
		17587: Delta = 44'sb11111111111111111111111111111111111111100000;
		64: Delta = 44'sb00000000000000000000000000000000000001000000;
		17555: Delta = 44'sb11111111111111111111111111111111111111000000;
		128: Delta = 44'sb00000000000000000000000000000000000010000000;
		17491: Delta = 44'sb11111111111111111111111111111111111110000000;
		256: Delta = 44'sb00000000000000000000000000000000000100000000;
		17363: Delta = 44'sb11111111111111111111111111111111111100000000;
		512: Delta = 44'sb00000000000000000000000000000000001000000000;
		17107: Delta = 44'sb11111111111111111111111111111111111000000000;
		1024: Delta = 44'sb00000000000000000000000000000000010000000000;
		16595: Delta = 44'sb11111111111111111111111111111111110000000000;
		2048: Delta = 44'sb00000000000000000000000000000000100000000000;
		15571: Delta = 44'sb11111111111111111111111111111111100000000000;
		4096: Delta = 44'sb00000000000000000000000000000001000000000000;
		13523: Delta = 44'sb11111111111111111111111111111111000000000000;
		8192: Delta = 44'sb00000000000000000000000000000010000000000000;
		9427: Delta = 44'sb11111111111111111111111111111110000000000000;
		16384: Delta = 44'sb00000000000000000000000000000100000000000000;
		1235: Delta = 44'sb11111111111111111111111111111100000000000000;
		15149: Delta = 44'sb00000000000000000000000000001000000000000000;
		2470: Delta = 44'sb11111111111111111111111111111000000000000000;
		12679: Delta = 44'sb00000000000000000000000000010000000000000000;
		4940: Delta = 44'sb11111111111111111111111111110000000000000000;
		7739: Delta = 44'sb00000000000000000000000000100000000000000000;
		9880: Delta = 44'sb11111111111111111111111111100000000000000000;
		15478: Delta = 44'sb00000000000000000000000001000000000000000000;
		2141: Delta = 44'sb11111111111111111111111111000000000000000000;
		13337: Delta = 44'sb00000000000000000000000010000000000000000000;
		4282: Delta = 44'sb11111111111111111111111110000000000000000000;
		9055: Delta = 44'sb00000000000000000000000100000000000000000000;
		8564: Delta = 44'sb11111111111111111111111100000000000000000000;
		491: Delta = 44'sb00000000000000000000001000000000000000000000;
		17128: Delta = 44'sb11111111111111111111111000000000000000000000;
		982: Delta = 44'sb00000000000000000000010000000000000000000000;
		16637: Delta = 44'sb11111111111111111111110000000000000000000000;
		1964: Delta = 44'sb00000000000000000000100000000000000000000000;
		15655: Delta = 44'sb11111111111111111111100000000000000000000000;
		3928: Delta = 44'sb00000000000000000001000000000000000000000000;
		13691: Delta = 44'sb11111111111111111111000000000000000000000000;
		7856: Delta = 44'sb00000000000000000010000000000000000000000000;
		9763: Delta = 44'sb11111111111111111110000000000000000000000000;
		15712: Delta = 44'sb00000000000000000100000000000000000000000000;
		1907: Delta = 44'sb11111111111111111100000000000000000000000000;
		13805: Delta = 44'sb00000000000000001000000000000000000000000000;
		3814: Delta = 44'sb11111111111111111000000000000000000000000000;
		9991: Delta = 44'sb00000000000000010000000000000000000000000000;
		7628: Delta = 44'sb11111111111111110000000000000000000000000000;
		2363: Delta = 44'sb00000000000000100000000000000000000000000000;
		15256: Delta = 44'sb11111111111111100000000000000000000000000000;
		4726: Delta = 44'sb00000000000001000000000000000000000000000000;
		12893: Delta = 44'sb11111111111111000000000000000000000000000000;
		9452: Delta = 44'sb00000000000010000000000000000000000000000000;
		8167: Delta = 44'sb11111111111110000000000000000000000000000000;
		1285: Delta = 44'sb00000000000100000000000000000000000000000000;
		16334: Delta = 44'sb11111111111100000000000000000000000000000000;
		2570: Delta = 44'sb00000000001000000000000000000000000000000000;
		15049: Delta = 44'sb11111111111000000000000000000000000000000000;
		5140: Delta = 44'sb00000000010000000000000000000000000000000000;
		12479: Delta = 44'sb11111111110000000000000000000000000000000000;
		10280: Delta = 44'sb00000000100000000000000000000000000000000000;
		7339: Delta = 44'sb11111111100000000000000000000000000000000000;
		2941: Delta = 44'sb00000001000000000000000000000000000000000000;
		14678: Delta = 44'sb11111111000000000000000000000000000000000000;
		5882: Delta = 44'sb00000010000000000000000000000000000000000000;
		11737: Delta = 44'sb11111110000000000000000000000000000000000000;
		11764: Delta = 44'sb00000100000000000000000000000000000000000000;
		5855: Delta = 44'sb11111100000000000000000000000000000000000000;
		5909: Delta = 44'sb00001000000000000000000000000000000000000000;
		11710: Delta = 44'sb11111000000000000000000000000000000000000000;
		11818: Delta = 44'sb00010000000000000000000000000000000000000000;
		5801: Delta = 44'sb11110000000000000000000000000000000000000000;
		6017: Delta = 44'sb00100000000000000000000000000000000000000000;
		11602: Delta = 44'sb11100000000000000000000000000000000000000000;
		12034: Delta = 44'sb01000000000000000000000000000000000000000000;
		5585: Delta = 44'sb11000000000000000000000000000000000000000000;
		default: Delta =44'sb0;
	endcase
end

assign N = (W - Delta) / A;

endmodule

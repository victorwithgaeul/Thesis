// Product (AN) Code DEC r-LUT
// DEC_rLUT16bits.v
// Used to do DEC, but corrected errors by locations, not AWE
// Received remainder r, output two error locations.
module DEC_rLUT16bits(r, l_1, l_2);
input 	[12:0]	r;
output	reg	signed	[5:0]	l_1;
output	reg	signed	[5:0]	l_2;
always@(*) begin
	case(r)
		1: begin l_1 = -1;
				 l_2 = +2; end
		4546: begin l_1 = +1;
				 l_2 = -2; end
		2: begin l_1 = +1;
				 l_2 = +1; end
		4545: begin l_1 = -1;
				 l_2 = -1; end
		4: begin l_1 = +2;
				 l_2 = +2; end
		4543: begin l_1 = -2;
				 l_2 = -2; end
		8: begin l_1 = +3;
				 l_2 = +3; end
		4539: begin l_1 = -3;
				 l_2 = -3; end
		16: begin l_1 = +4;
				 l_2 = +4; end
		4531: begin l_1 = -4;
				 l_2 = -4; end
		32: begin l_1 = +5;
				 l_2 = +5; end
		4515: begin l_1 = -5;
				 l_2 = -5; end
		64: begin l_1 = +6;
				 l_2 = +6; end
		4483: begin l_1 = -6;
				 l_2 = -6; end
		128: begin l_1 = +7;
				 l_2 = +7; end
		4419: begin l_1 = -7;
				 l_2 = -7; end
		256: begin l_1 = +8;
				 l_2 = +8; end
		4291: begin l_1 = -8;
				 l_2 = -8; end
		512: begin l_1 = +9;
				 l_2 = +9; end
		4035: begin l_1 = -9;
				 l_2 = -9; end
		1024: begin l_1 = +10;
				 l_2 = +10; end
		3523: begin l_1 = -10;
				 l_2 = -10; end
		2048: begin l_1 = +11;
				 l_2 = +11; end
		2499: begin l_1 = -11;
				 l_2 = -11; end
		4096: begin l_1 = +12;
				 l_2 = +12; end
		451: begin l_1 = -12;
				 l_2 = -12; end
		3645: begin l_1 = +13;
				 l_2 = +13; end
		902: begin l_1 = -13;
				 l_2 = -13; end
		2743: begin l_1 = +14;
				 l_2 = +14; end
		1804: begin l_1 = -14;
				 l_2 = -14; end
		939: begin l_1 = +15;
				 l_2 = +15; end
		3608: begin l_1 = -15;
				 l_2 = -15; end
		1878: begin l_1 = +16;
				 l_2 = +16; end
		2669: begin l_1 = -16;
				 l_2 = -16; end
		3756: begin l_1 = +17;
				 l_2 = +17; end
		791: begin l_1 = -17;
				 l_2 = -17; end
		2965: begin l_1 = +18;
				 l_2 = +18; end
		1582: begin l_1 = -18;
				 l_2 = -18; end
		1383: begin l_1 = +19;
				 l_2 = +19; end
		3164: begin l_1 = -19;
				 l_2 = -19; end
		2766: begin l_1 = +20;
				 l_2 = +20; end
		1781: begin l_1 = -20;
				 l_2 = -20; end
		985: begin l_1 = +21;
				 l_2 = +21; end
		3562: begin l_1 = -21;
				 l_2 = -21; end
		1970: begin l_1 = +22;
				 l_2 = +22; end
		2577: begin l_1 = -22;
				 l_2 = -22; end
		3940: begin l_1 = +23;
				 l_2 = +23; end
		607: begin l_1 = -23;
				 l_2 = -23; end
		3333: begin l_1 = +24;
				 l_2 = +24; end
		1214: begin l_1 = -24;
				 l_2 = -24; end
		2119: begin l_1 = +25;
				 l_2 = +25; end
		2428: begin l_1 = -25;
				 l_2 = -25; end
		4238: begin l_1 = +26;
				 l_2 = +26; end
		309: begin l_1 = -26;
				 l_2 = -26; end
		3929: begin l_1 = +27;
				 l_2 = +27; end
		618: begin l_1 = -27;
				 l_2 = -27; end
		3311: begin l_1 = +28;
				 l_2 = +28; end
		1236: begin l_1 = -28;
				 l_2 = -28; end
		3: begin l_1 = -1;
				 l_2 = +3; end
		4544: begin l_1 = -1;
				 l_2 = -2; end
		5: begin l_1 = +1;
				 l_2 = +3; end
		4542: begin l_1 = -1;
				 l_2 = -3; end
		9: begin l_1 = +1;
				 l_2 = +4; end
		4540: begin l_1 = +1;
				 l_2 = -4; end
		7: begin l_1 = -1;
				 l_2 = +4; end
		4538: begin l_1 = -1;
				 l_2 = -4; end
		17: begin l_1 = +1;
				 l_2 = +5; end
		4532: begin l_1 = +1;
				 l_2 = -5; end
		15: begin l_1 = -1;
				 l_2 = +5; end
		4530: begin l_1 = -1;
				 l_2 = -5; end
		33: begin l_1 = +1;
				 l_2 = +6; end
		4516: begin l_1 = +1;
				 l_2 = -6; end
		31: begin l_1 = -1;
				 l_2 = +6; end
		4514: begin l_1 = -1;
				 l_2 = -6; end
		65: begin l_1 = +1;
				 l_2 = +7; end
		4484: begin l_1 = +1;
				 l_2 = -7; end
		63: begin l_1 = -1;
				 l_2 = +7; end
		4482: begin l_1 = -1;
				 l_2 = -7; end
		129: begin l_1 = +1;
				 l_2 = +8; end
		4420: begin l_1 = +1;
				 l_2 = -8; end
		127: begin l_1 = -1;
				 l_2 = +8; end
		4418: begin l_1 = -1;
				 l_2 = -8; end
		257: begin l_1 = +1;
				 l_2 = +9; end
		4292: begin l_1 = +1;
				 l_2 = -9; end
		255: begin l_1 = -1;
				 l_2 = +9; end
		4290: begin l_1 = -1;
				 l_2 = -9; end
		513: begin l_1 = +1;
				 l_2 = +10; end
		4036: begin l_1 = +1;
				 l_2 = -10; end
		511: begin l_1 = -1;
				 l_2 = +10; end
		4034: begin l_1 = -1;
				 l_2 = -10; end
		1025: begin l_1 = +1;
				 l_2 = +11; end
		3524: begin l_1 = +1;
				 l_2 = -11; end
		1023: begin l_1 = -1;
				 l_2 = +11; end
		3522: begin l_1 = -1;
				 l_2 = -11; end
		2049: begin l_1 = +1;
				 l_2 = +12; end
		2500: begin l_1 = +1;
				 l_2 = -12; end
		2047: begin l_1 = -1;
				 l_2 = +12; end
		2498: begin l_1 = -1;
				 l_2 = -12; end
		4097: begin l_1 = +1;
				 l_2 = +13; end
		452: begin l_1 = +1;
				 l_2 = -13; end
		4095: begin l_1 = -1;
				 l_2 = +13; end
		450: begin l_1 = -1;
				 l_2 = -13; end
		3646: begin l_1 = +1;
				 l_2 = +14; end
		903: begin l_1 = +1;
				 l_2 = -14; end
		3644: begin l_1 = -1;
				 l_2 = +14; end
		901: begin l_1 = -1;
				 l_2 = -14; end
		2744: begin l_1 = +1;
				 l_2 = +15; end
		1805: begin l_1 = +1;
				 l_2 = -15; end
		2742: begin l_1 = -1;
				 l_2 = +15; end
		1803: begin l_1 = -1;
				 l_2 = -15; end
		940: begin l_1 = +1;
				 l_2 = +16; end
		3609: begin l_1 = +1;
				 l_2 = -16; end
		938: begin l_1 = -1;
				 l_2 = +16; end
		3607: begin l_1 = -1;
				 l_2 = -16; end
		1879: begin l_1 = +1;
				 l_2 = +17; end
		2670: begin l_1 = +1;
				 l_2 = -17; end
		1877: begin l_1 = -1;
				 l_2 = +17; end
		2668: begin l_1 = -1;
				 l_2 = -17; end
		3757: begin l_1 = +1;
				 l_2 = +18; end
		792: begin l_1 = +1;
				 l_2 = -18; end
		3755: begin l_1 = -1;
				 l_2 = +18; end
		790: begin l_1 = -1;
				 l_2 = -18; end
		2966: begin l_1 = +1;
				 l_2 = +19; end
		1583: begin l_1 = +1;
				 l_2 = -19; end
		2964: begin l_1 = -1;
				 l_2 = +19; end
		1581: begin l_1 = -1;
				 l_2 = -19; end
		1384: begin l_1 = +1;
				 l_2 = +20; end
		3165: begin l_1 = +1;
				 l_2 = -20; end
		1382: begin l_1 = -1;
				 l_2 = +20; end
		3163: begin l_1 = -1;
				 l_2 = -20; end
		2767: begin l_1 = +1;
				 l_2 = +21; end
		1782: begin l_1 = +1;
				 l_2 = -21; end
		2765: begin l_1 = -1;
				 l_2 = +21; end
		1780: begin l_1 = -1;
				 l_2 = -21; end
		986: begin l_1 = +1;
				 l_2 = +22; end
		3563: begin l_1 = +1;
				 l_2 = -22; end
		984: begin l_1 = -1;
				 l_2 = +22; end
		3561: begin l_1 = -1;
				 l_2 = -22; end
		1971: begin l_1 = +1;
				 l_2 = +23; end
		2578: begin l_1 = +1;
				 l_2 = -23; end
		1969: begin l_1 = -1;
				 l_2 = +23; end
		2576: begin l_1 = -1;
				 l_2 = -23; end
		3941: begin l_1 = +1;
				 l_2 = +24; end
		608: begin l_1 = +1;
				 l_2 = -24; end
		3939: begin l_1 = -1;
				 l_2 = +24; end
		606: begin l_1 = -1;
				 l_2 = -24; end
		3334: begin l_1 = +1;
				 l_2 = +25; end
		1215: begin l_1 = +1;
				 l_2 = -25; end
		3332: begin l_1 = -1;
				 l_2 = +25; end
		1213: begin l_1 = -1;
				 l_2 = -25; end
		2120: begin l_1 = +1;
				 l_2 = +26; end
		2429: begin l_1 = +1;
				 l_2 = -26; end
		2118: begin l_1 = -1;
				 l_2 = +26; end
		2427: begin l_1 = -1;
				 l_2 = -26; end
		4239: begin l_1 = +1;
				 l_2 = +27; end
		310: begin l_1 = +1;
				 l_2 = -27; end
		4237: begin l_1 = -1;
				 l_2 = +27; end
		308: begin l_1 = -1;
				 l_2 = -27; end
		3930: begin l_1 = +1;
				 l_2 = +28; end
		619: begin l_1 = +1;
				 l_2 = -28; end
		3928: begin l_1 = -1;
				 l_2 = +28; end
		617: begin l_1 = -1;
				 l_2 = -28; end
		3312: begin l_1 = +1;
				 l_2 = +29; end
		1237: begin l_1 = +1;
				 l_2 = -29; end
		3310: begin l_1 = -1;
				 l_2 = +29; end
		1235: begin l_1 = -1;
				 l_2 = -29; end
		6: begin l_1 = -2;
				 l_2 = +4; end
		4541: begin l_1 = -2;
				 l_2 = -3; end
		10: begin l_1 = +2;
				 l_2 = +4; end
		4537: begin l_1 = -2;
				 l_2 = -4; end
		18: begin l_1 = +2;
				 l_2 = +5; end
		4533: begin l_1 = +2;
				 l_2 = -5; end
		14: begin l_1 = -2;
				 l_2 = +5; end
		4529: begin l_1 = -2;
				 l_2 = -5; end
		34: begin l_1 = +2;
				 l_2 = +6; end
		4517: begin l_1 = +2;
				 l_2 = -6; end
		30: begin l_1 = -2;
				 l_2 = +6; end
		4513: begin l_1 = -2;
				 l_2 = -6; end
		66: begin l_1 = +2;
				 l_2 = +7; end
		4485: begin l_1 = +2;
				 l_2 = -7; end
		62: begin l_1 = -2;
				 l_2 = +7; end
		4481: begin l_1 = -2;
				 l_2 = -7; end
		130: begin l_1 = +2;
				 l_2 = +8; end
		4421: begin l_1 = +2;
				 l_2 = -8; end
		126: begin l_1 = -2;
				 l_2 = +8; end
		4417: begin l_1 = -2;
				 l_2 = -8; end
		258: begin l_1 = +2;
				 l_2 = +9; end
		4293: begin l_1 = +2;
				 l_2 = -9; end
		254: begin l_1 = -2;
				 l_2 = +9; end
		4289: begin l_1 = -2;
				 l_2 = -9; end
		514: begin l_1 = +2;
				 l_2 = +10; end
		4037: begin l_1 = +2;
				 l_2 = -10; end
		510: begin l_1 = -2;
				 l_2 = +10; end
		4033: begin l_1 = -2;
				 l_2 = -10; end
		1026: begin l_1 = +2;
				 l_2 = +11; end
		3525: begin l_1 = +2;
				 l_2 = -11; end
		1022: begin l_1 = -2;
				 l_2 = +11; end
		3521: begin l_1 = -2;
				 l_2 = -11; end
		2050: begin l_1 = +2;
				 l_2 = +12; end
		2501: begin l_1 = +2;
				 l_2 = -12; end
		2046: begin l_1 = -2;
				 l_2 = +12; end
		2497: begin l_1 = -2;
				 l_2 = -12; end
		4098: begin l_1 = +2;
				 l_2 = +13; end
		453: begin l_1 = +2;
				 l_2 = -13; end
		4094: begin l_1 = -2;
				 l_2 = +13; end
		449: begin l_1 = -2;
				 l_2 = -13; end
		3647: begin l_1 = +2;
				 l_2 = +14; end
		904: begin l_1 = +2;
				 l_2 = -14; end
		3643: begin l_1 = -2;
				 l_2 = +14; end
		900: begin l_1 = -2;
				 l_2 = -14; end
		2745: begin l_1 = +2;
				 l_2 = +15; end
		1806: begin l_1 = +2;
				 l_2 = -15; end
		2741: begin l_1 = -2;
				 l_2 = +15; end
		1802: begin l_1 = -2;
				 l_2 = -15; end
		941: begin l_1 = +2;
				 l_2 = +16; end
		3610: begin l_1 = +2;
				 l_2 = -16; end
		937: begin l_1 = -2;
				 l_2 = +16; end
		3606: begin l_1 = -2;
				 l_2 = -16; end
		1880: begin l_1 = +2;
				 l_2 = +17; end
		2671: begin l_1 = +2;
				 l_2 = -17; end
		1876: begin l_1 = -2;
				 l_2 = +17; end
		2667: begin l_1 = -2;
				 l_2 = -17; end
		3758: begin l_1 = +2;
				 l_2 = +18; end
		793: begin l_1 = +2;
				 l_2 = -18; end
		3754: begin l_1 = -2;
				 l_2 = +18; end
		789: begin l_1 = -2;
				 l_2 = -18; end
		2967: begin l_1 = +2;
				 l_2 = +19; end
		1584: begin l_1 = +2;
				 l_2 = -19; end
		2963: begin l_1 = -2;
				 l_2 = +19; end
		1580: begin l_1 = -2;
				 l_2 = -19; end
		1385: begin l_1 = +2;
				 l_2 = +20; end
		3166: begin l_1 = +2;
				 l_2 = -20; end
		1381: begin l_1 = -2;
				 l_2 = +20; end
		3162: begin l_1 = -2;
				 l_2 = -20; end
		2768: begin l_1 = +2;
				 l_2 = +21; end
		1783: begin l_1 = +2;
				 l_2 = -21; end
		2764: begin l_1 = -2;
				 l_2 = +21; end
		1779: begin l_1 = -2;
				 l_2 = -21; end
		987: begin l_1 = +2;
				 l_2 = +22; end
		3564: begin l_1 = +2;
				 l_2 = -22; end
		983: begin l_1 = -2;
				 l_2 = +22; end
		3560: begin l_1 = -2;
				 l_2 = -22; end
		1972: begin l_1 = +2;
				 l_2 = +23; end
		2579: begin l_1 = +2;
				 l_2 = -23; end
		1968: begin l_1 = -2;
				 l_2 = +23; end
		2575: begin l_1 = -2;
				 l_2 = -23; end
		3942: begin l_1 = +2;
				 l_2 = +24; end
		609: begin l_1 = +2;
				 l_2 = -24; end
		3938: begin l_1 = -2;
				 l_2 = +24; end
		605: begin l_1 = -2;
				 l_2 = -24; end
		3335: begin l_1 = +2;
				 l_2 = +25; end
		1216: begin l_1 = +2;
				 l_2 = -25; end
		3331: begin l_1 = -2;
				 l_2 = +25; end
		1212: begin l_1 = -2;
				 l_2 = -25; end
		2121: begin l_1 = +2;
				 l_2 = +26; end
		2430: begin l_1 = +2;
				 l_2 = -26; end
		2117: begin l_1 = -2;
				 l_2 = +26; end
		2426: begin l_1 = -2;
				 l_2 = -26; end
		4240: begin l_1 = +2;
				 l_2 = +27; end
		311: begin l_1 = +2;
				 l_2 = -27; end
		4236: begin l_1 = -2;
				 l_2 = +27; end
		307: begin l_1 = -2;
				 l_2 = -27; end
		3931: begin l_1 = +2;
				 l_2 = +28; end
		620: begin l_1 = +2;
				 l_2 = -28; end
		3927: begin l_1 = -2;
				 l_2 = +28; end
		616: begin l_1 = -2;
				 l_2 = -28; end
		3313: begin l_1 = +2;
				 l_2 = +29; end
		1238: begin l_1 = +2;
				 l_2 = -29; end
		3309: begin l_1 = -2;
				 l_2 = +29; end
		1234: begin l_1 = -2;
				 l_2 = -29; end
		12: begin l_1 = -3;
				 l_2 = +5; end
		4535: begin l_1 = -3;
				 l_2 = -4; end
		20: begin l_1 = +3;
				 l_2 = +5; end
		4527: begin l_1 = -3;
				 l_2 = -5; end
		36: begin l_1 = +3;
				 l_2 = +6; end
		4519: begin l_1 = +3;
				 l_2 = -6; end
		28: begin l_1 = -3;
				 l_2 = +6; end
		4511: begin l_1 = -3;
				 l_2 = -6; end
		68: begin l_1 = +3;
				 l_2 = +7; end
		4487: begin l_1 = +3;
				 l_2 = -7; end
		60: begin l_1 = -3;
				 l_2 = +7; end
		4479: begin l_1 = -3;
				 l_2 = -7; end
		132: begin l_1 = +3;
				 l_2 = +8; end
		4423: begin l_1 = +3;
				 l_2 = -8; end
		124: begin l_1 = -3;
				 l_2 = +8; end
		4415: begin l_1 = -3;
				 l_2 = -8; end
		260: begin l_1 = +3;
				 l_2 = +9; end
		4295: begin l_1 = +3;
				 l_2 = -9; end
		252: begin l_1 = -3;
				 l_2 = +9; end
		4287: begin l_1 = -3;
				 l_2 = -9; end
		516: begin l_1 = +3;
				 l_2 = +10; end
		4039: begin l_1 = +3;
				 l_2 = -10; end
		508: begin l_1 = -3;
				 l_2 = +10; end
		4031: begin l_1 = -3;
				 l_2 = -10; end
		1028: begin l_1 = +3;
				 l_2 = +11; end
		3527: begin l_1 = +3;
				 l_2 = -11; end
		1020: begin l_1 = -3;
				 l_2 = +11; end
		3519: begin l_1 = -3;
				 l_2 = -11; end
		2052: begin l_1 = +3;
				 l_2 = +12; end
		2503: begin l_1 = +3;
				 l_2 = -12; end
		2044: begin l_1 = -3;
				 l_2 = +12; end
		2495: begin l_1 = -3;
				 l_2 = -12; end
		4100: begin l_1 = +3;
				 l_2 = +13; end
		455: begin l_1 = +3;
				 l_2 = -13; end
		4092: begin l_1 = -3;
				 l_2 = +13; end
		447: begin l_1 = -3;
				 l_2 = -13; end
		3649: begin l_1 = +3;
				 l_2 = +14; end
		906: begin l_1 = +3;
				 l_2 = -14; end
		3641: begin l_1 = -3;
				 l_2 = +14; end
		898: begin l_1 = -3;
				 l_2 = -14; end
		2747: begin l_1 = +3;
				 l_2 = +15; end
		1808: begin l_1 = +3;
				 l_2 = -15; end
		2739: begin l_1 = -3;
				 l_2 = +15; end
		1800: begin l_1 = -3;
				 l_2 = -15; end
		943: begin l_1 = +3;
				 l_2 = +16; end
		3612: begin l_1 = +3;
				 l_2 = -16; end
		935: begin l_1 = -3;
				 l_2 = +16; end
		3604: begin l_1 = -3;
				 l_2 = -16; end
		1882: begin l_1 = +3;
				 l_2 = +17; end
		2673: begin l_1 = +3;
				 l_2 = -17; end
		1874: begin l_1 = -3;
				 l_2 = +17; end
		2665: begin l_1 = -3;
				 l_2 = -17; end
		3760: begin l_1 = +3;
				 l_2 = +18; end
		795: begin l_1 = +3;
				 l_2 = -18; end
		3752: begin l_1 = -3;
				 l_2 = +18; end
		787: begin l_1 = -3;
				 l_2 = -18; end
		2969: begin l_1 = +3;
				 l_2 = +19; end
		1586: begin l_1 = +3;
				 l_2 = -19; end
		2961: begin l_1 = -3;
				 l_2 = +19; end
		1578: begin l_1 = -3;
				 l_2 = -19; end
		1387: begin l_1 = +3;
				 l_2 = +20; end
		3168: begin l_1 = +3;
				 l_2 = -20; end
		1379: begin l_1 = -3;
				 l_2 = +20; end
		3160: begin l_1 = -3;
				 l_2 = -20; end
		2770: begin l_1 = +3;
				 l_2 = +21; end
		1785: begin l_1 = +3;
				 l_2 = -21; end
		2762: begin l_1 = -3;
				 l_2 = +21; end
		1777: begin l_1 = -3;
				 l_2 = -21; end
		989: begin l_1 = +3;
				 l_2 = +22; end
		3566: begin l_1 = +3;
				 l_2 = -22; end
		981: begin l_1 = -3;
				 l_2 = +22; end
		3558: begin l_1 = -3;
				 l_2 = -22; end
		1974: begin l_1 = +3;
				 l_2 = +23; end
		2581: begin l_1 = +3;
				 l_2 = -23; end
		1966: begin l_1 = -3;
				 l_2 = +23; end
		2573: begin l_1 = -3;
				 l_2 = -23; end
		3944: begin l_1 = +3;
				 l_2 = +24; end
		611: begin l_1 = +3;
				 l_2 = -24; end
		3936: begin l_1 = -3;
				 l_2 = +24; end
		603: begin l_1 = -3;
				 l_2 = -24; end
		3337: begin l_1 = +3;
				 l_2 = +25; end
		1218: begin l_1 = +3;
				 l_2 = -25; end
		3329: begin l_1 = -3;
				 l_2 = +25; end
		1210: begin l_1 = -3;
				 l_2 = -25; end
		2123: begin l_1 = +3;
				 l_2 = +26; end
		2432: begin l_1 = +3;
				 l_2 = -26; end
		2115: begin l_1 = -3;
				 l_2 = +26; end
		2424: begin l_1 = -3;
				 l_2 = -26; end
		4242: begin l_1 = +3;
				 l_2 = +27; end
		313: begin l_1 = +3;
				 l_2 = -27; end
		4234: begin l_1 = -3;
				 l_2 = +27; end
		305: begin l_1 = -3;
				 l_2 = -27; end
		3933: begin l_1 = +3;
				 l_2 = +28; end
		622: begin l_1 = +3;
				 l_2 = -28; end
		3925: begin l_1 = -3;
				 l_2 = +28; end
		614: begin l_1 = -3;
				 l_2 = -28; end
		3315: begin l_1 = +3;
				 l_2 = +29; end
		1240: begin l_1 = +3;
				 l_2 = -29; end
		3307: begin l_1 = -3;
				 l_2 = +29; end
		1232: begin l_1 = -3;
				 l_2 = -29; end
		24: begin l_1 = -4;
				 l_2 = +6; end
		4523: begin l_1 = -4;
				 l_2 = -5; end
		40: begin l_1 = +4;
				 l_2 = +6; end
		4507: begin l_1 = -4;
				 l_2 = -6; end
		72: begin l_1 = +4;
				 l_2 = +7; end
		4491: begin l_1 = +4;
				 l_2 = -7; end
		56: begin l_1 = -4;
				 l_2 = +7; end
		4475: begin l_1 = -4;
				 l_2 = -7; end
		136: begin l_1 = +4;
				 l_2 = +8; end
		4427: begin l_1 = +4;
				 l_2 = -8; end
		120: begin l_1 = -4;
				 l_2 = +8; end
		4411: begin l_1 = -4;
				 l_2 = -8; end
		264: begin l_1 = +4;
				 l_2 = +9; end
		4299: begin l_1 = +4;
				 l_2 = -9; end
		248: begin l_1 = -4;
				 l_2 = +9; end
		4283: begin l_1 = -4;
				 l_2 = -9; end
		520: begin l_1 = +4;
				 l_2 = +10; end
		4043: begin l_1 = +4;
				 l_2 = -10; end
		504: begin l_1 = -4;
				 l_2 = +10; end
		4027: begin l_1 = -4;
				 l_2 = -10; end
		1032: begin l_1 = +4;
				 l_2 = +11; end
		3531: begin l_1 = +4;
				 l_2 = -11; end
		1016: begin l_1 = -4;
				 l_2 = +11; end
		3515: begin l_1 = -4;
				 l_2 = -11; end
		2056: begin l_1 = +4;
				 l_2 = +12; end
		2507: begin l_1 = +4;
				 l_2 = -12; end
		2040: begin l_1 = -4;
				 l_2 = +12; end
		2491: begin l_1 = -4;
				 l_2 = -12; end
		4104: begin l_1 = +4;
				 l_2 = +13; end
		459: begin l_1 = +4;
				 l_2 = -13; end
		4088: begin l_1 = -4;
				 l_2 = +13; end
		443: begin l_1 = -4;
				 l_2 = -13; end
		3653: begin l_1 = +4;
				 l_2 = +14; end
		910: begin l_1 = +4;
				 l_2 = -14; end
		3637: begin l_1 = -4;
				 l_2 = +14; end
		894: begin l_1 = -4;
				 l_2 = -14; end
		2751: begin l_1 = +4;
				 l_2 = +15; end
		1812: begin l_1 = +4;
				 l_2 = -15; end
		2735: begin l_1 = -4;
				 l_2 = +15; end
		1796: begin l_1 = -4;
				 l_2 = -15; end
		947: begin l_1 = +4;
				 l_2 = +16; end
		3616: begin l_1 = +4;
				 l_2 = -16; end
		931: begin l_1 = -4;
				 l_2 = +16; end
		3600: begin l_1 = -4;
				 l_2 = -16; end
		1886: begin l_1 = +4;
				 l_2 = +17; end
		2677: begin l_1 = +4;
				 l_2 = -17; end
		1870: begin l_1 = -4;
				 l_2 = +17; end
		2661: begin l_1 = -4;
				 l_2 = -17; end
		3764: begin l_1 = +4;
				 l_2 = +18; end
		799: begin l_1 = +4;
				 l_2 = -18; end
		3748: begin l_1 = -4;
				 l_2 = +18; end
		783: begin l_1 = -4;
				 l_2 = -18; end
		2973: begin l_1 = +4;
				 l_2 = +19; end
		1590: begin l_1 = +4;
				 l_2 = -19; end
		2957: begin l_1 = -4;
				 l_2 = +19; end
		1574: begin l_1 = -4;
				 l_2 = -19; end
		1391: begin l_1 = +4;
				 l_2 = +20; end
		3172: begin l_1 = +4;
				 l_2 = -20; end
		1375: begin l_1 = -4;
				 l_2 = +20; end
		3156: begin l_1 = -4;
				 l_2 = -20; end
		2774: begin l_1 = +4;
				 l_2 = +21; end
		1789: begin l_1 = +4;
				 l_2 = -21; end
		2758: begin l_1 = -4;
				 l_2 = +21; end
		1773: begin l_1 = -4;
				 l_2 = -21; end
		993: begin l_1 = +4;
				 l_2 = +22; end
		3570: begin l_1 = +4;
				 l_2 = -22; end
		977: begin l_1 = -4;
				 l_2 = +22; end
		3554: begin l_1 = -4;
				 l_2 = -22; end
		1978: begin l_1 = +4;
				 l_2 = +23; end
		2585: begin l_1 = +4;
				 l_2 = -23; end
		1962: begin l_1 = -4;
				 l_2 = +23; end
		2569: begin l_1 = -4;
				 l_2 = -23; end
		3948: begin l_1 = +4;
				 l_2 = +24; end
		615: begin l_1 = +4;
				 l_2 = -24; end
		3932: begin l_1 = -4;
				 l_2 = +24; end
		599: begin l_1 = -4;
				 l_2 = -24; end
		3341: begin l_1 = +4;
				 l_2 = +25; end
		1222: begin l_1 = +4;
				 l_2 = -25; end
		3325: begin l_1 = -4;
				 l_2 = +25; end
		1206: begin l_1 = -4;
				 l_2 = -25; end
		2127: begin l_1 = +4;
				 l_2 = +26; end
		2436: begin l_1 = +4;
				 l_2 = -26; end
		2111: begin l_1 = -4;
				 l_2 = +26; end
		2420: begin l_1 = -4;
				 l_2 = -26; end
		4246: begin l_1 = +4;
				 l_2 = +27; end
		317: begin l_1 = +4;
				 l_2 = -27; end
		4230: begin l_1 = -4;
				 l_2 = +27; end
		301: begin l_1 = -4;
				 l_2 = -27; end
		3937: begin l_1 = +4;
				 l_2 = +28; end
		626: begin l_1 = +4;
				 l_2 = -28; end
		3921: begin l_1 = -4;
				 l_2 = +28; end
		610: begin l_1 = -4;
				 l_2 = -28; end
		3319: begin l_1 = +4;
				 l_2 = +29; end
		1244: begin l_1 = +4;
				 l_2 = -29; end
		3303: begin l_1 = -4;
				 l_2 = +29; end
		1228: begin l_1 = -4;
				 l_2 = -29; end
		48: begin l_1 = -5;
				 l_2 = +7; end
		4499: begin l_1 = -5;
				 l_2 = -6; end
		80: begin l_1 = +5;
				 l_2 = +7; end
		4467: begin l_1 = -5;
				 l_2 = -7; end
		144: begin l_1 = +5;
				 l_2 = +8; end
		4435: begin l_1 = +5;
				 l_2 = -8; end
		112: begin l_1 = -5;
				 l_2 = +8; end
		4403: begin l_1 = -5;
				 l_2 = -8; end
		272: begin l_1 = +5;
				 l_2 = +9; end
		4307: begin l_1 = +5;
				 l_2 = -9; end
		240: begin l_1 = -5;
				 l_2 = +9; end
		4275: begin l_1 = -5;
				 l_2 = -9; end
		528: begin l_1 = +5;
				 l_2 = +10; end
		4051: begin l_1 = +5;
				 l_2 = -10; end
		496: begin l_1 = -5;
				 l_2 = +10; end
		4019: begin l_1 = -5;
				 l_2 = -10; end
		1040: begin l_1 = +5;
				 l_2 = +11; end
		3539: begin l_1 = +5;
				 l_2 = -11; end
		1008: begin l_1 = -5;
				 l_2 = +11; end
		3507: begin l_1 = -5;
				 l_2 = -11; end
		2064: begin l_1 = +5;
				 l_2 = +12; end
		2515: begin l_1 = +5;
				 l_2 = -12; end
		2032: begin l_1 = -5;
				 l_2 = +12; end
		2483: begin l_1 = -5;
				 l_2 = -12; end
		4112: begin l_1 = +5;
				 l_2 = +13; end
		467: begin l_1 = +5;
				 l_2 = -13; end
		4080: begin l_1 = -5;
				 l_2 = +13; end
		435: begin l_1 = -5;
				 l_2 = -13; end
		3661: begin l_1 = +5;
				 l_2 = +14; end
		918: begin l_1 = +5;
				 l_2 = -14; end
		3629: begin l_1 = -5;
				 l_2 = +14; end
		886: begin l_1 = -5;
				 l_2 = -14; end
		2759: begin l_1 = +5;
				 l_2 = +15; end
		1820: begin l_1 = +5;
				 l_2 = -15; end
		2727: begin l_1 = -5;
				 l_2 = +15; end
		1788: begin l_1 = -5;
				 l_2 = -15; end
		955: begin l_1 = +5;
				 l_2 = +16; end
		3624: begin l_1 = +5;
				 l_2 = -16; end
		923: begin l_1 = -5;
				 l_2 = +16; end
		3592: begin l_1 = -5;
				 l_2 = -16; end
		1894: begin l_1 = +5;
				 l_2 = +17; end
		2685: begin l_1 = +5;
				 l_2 = -17; end
		1862: begin l_1 = -5;
				 l_2 = +17; end
		2653: begin l_1 = -5;
				 l_2 = -17; end
		3772: begin l_1 = +5;
				 l_2 = +18; end
		807: begin l_1 = +5;
				 l_2 = -18; end
		3740: begin l_1 = -5;
				 l_2 = +18; end
		775: begin l_1 = -5;
				 l_2 = -18; end
		2981: begin l_1 = +5;
				 l_2 = +19; end
		1598: begin l_1 = +5;
				 l_2 = -19; end
		2949: begin l_1 = -5;
				 l_2 = +19; end
		1566: begin l_1 = -5;
				 l_2 = -19; end
		1399: begin l_1 = +5;
				 l_2 = +20; end
		3180: begin l_1 = +5;
				 l_2 = -20; end
		1367: begin l_1 = -5;
				 l_2 = +20; end
		3148: begin l_1 = -5;
				 l_2 = -20; end
		2782: begin l_1 = +5;
				 l_2 = +21; end
		1797: begin l_1 = +5;
				 l_2 = -21; end
		2750: begin l_1 = -5;
				 l_2 = +21; end
		1765: begin l_1 = -5;
				 l_2 = -21; end
		1001: begin l_1 = +5;
				 l_2 = +22; end
		3578: begin l_1 = +5;
				 l_2 = -22; end
		969: begin l_1 = -5;
				 l_2 = +22; end
		3546: begin l_1 = -5;
				 l_2 = -22; end
		1986: begin l_1 = +5;
				 l_2 = +23; end
		2593: begin l_1 = +5;
				 l_2 = -23; end
		1954: begin l_1 = -5;
				 l_2 = +23; end
		2561: begin l_1 = -5;
				 l_2 = -23; end
		3956: begin l_1 = +5;
				 l_2 = +24; end
		623: begin l_1 = +5;
				 l_2 = -24; end
		3924: begin l_1 = -5;
				 l_2 = +24; end
		591: begin l_1 = -5;
				 l_2 = -24; end
		3349: begin l_1 = +5;
				 l_2 = +25; end
		1230: begin l_1 = +5;
				 l_2 = -25; end
		3317: begin l_1 = -5;
				 l_2 = +25; end
		1198: begin l_1 = -5;
				 l_2 = -25; end
		2135: begin l_1 = +5;
				 l_2 = +26; end
		2444: begin l_1 = +5;
				 l_2 = -26; end
		2103: begin l_1 = -5;
				 l_2 = +26; end
		2412: begin l_1 = -5;
				 l_2 = -26; end
		4254: begin l_1 = +5;
				 l_2 = +27; end
		325: begin l_1 = +5;
				 l_2 = -27; end
		4222: begin l_1 = -5;
				 l_2 = +27; end
		293: begin l_1 = -5;
				 l_2 = -27; end
		3945: begin l_1 = +5;
				 l_2 = +28; end
		634: begin l_1 = +5;
				 l_2 = -28; end
		3913: begin l_1 = -5;
				 l_2 = +28; end
		602: begin l_1 = -5;
				 l_2 = -28; end
		3327: begin l_1 = +5;
				 l_2 = +29; end
		1252: begin l_1 = +5;
				 l_2 = -29; end
		3295: begin l_1 = -5;
				 l_2 = +29; end
		1220: begin l_1 = -5;
				 l_2 = -29; end
		96: begin l_1 = -6;
				 l_2 = +8; end
		4451: begin l_1 = -6;
				 l_2 = -7; end
		160: begin l_1 = +6;
				 l_2 = +8; end
		4387: begin l_1 = -6;
				 l_2 = -8; end
		288: begin l_1 = +6;
				 l_2 = +9; end
		4323: begin l_1 = +6;
				 l_2 = -9; end
		224: begin l_1 = -6;
				 l_2 = +9; end
		4259: begin l_1 = -6;
				 l_2 = -9; end
		544: begin l_1 = +6;
				 l_2 = +10; end
		4067: begin l_1 = +6;
				 l_2 = -10; end
		480: begin l_1 = -6;
				 l_2 = +10; end
		4003: begin l_1 = -6;
				 l_2 = -10; end
		1056: begin l_1 = +6;
				 l_2 = +11; end
		3555: begin l_1 = +6;
				 l_2 = -11; end
		992: begin l_1 = -6;
				 l_2 = +11; end
		3491: begin l_1 = -6;
				 l_2 = -11; end
		2080: begin l_1 = +6;
				 l_2 = +12; end
		2531: begin l_1 = +6;
				 l_2 = -12; end
		2016: begin l_1 = -6;
				 l_2 = +12; end
		2467: begin l_1 = -6;
				 l_2 = -12; end
		4128: begin l_1 = +6;
				 l_2 = +13; end
		483: begin l_1 = +6;
				 l_2 = -13; end
		4064: begin l_1 = -6;
				 l_2 = +13; end
		419: begin l_1 = -6;
				 l_2 = -13; end
		3677: begin l_1 = +6;
				 l_2 = +14; end
		934: begin l_1 = +6;
				 l_2 = -14; end
		3613: begin l_1 = -6;
				 l_2 = +14; end
		870: begin l_1 = -6;
				 l_2 = -14; end
		2775: begin l_1 = +6;
				 l_2 = +15; end
		1836: begin l_1 = +6;
				 l_2 = -15; end
		2711: begin l_1 = -6;
				 l_2 = +15; end
		1772: begin l_1 = -6;
				 l_2 = -15; end
		971: begin l_1 = +6;
				 l_2 = +16; end
		3640: begin l_1 = +6;
				 l_2 = -16; end
		907: begin l_1 = -6;
				 l_2 = +16; end
		3576: begin l_1 = -6;
				 l_2 = -16; end
		1910: begin l_1 = +6;
				 l_2 = +17; end
		2701: begin l_1 = +6;
				 l_2 = -17; end
		1846: begin l_1 = -6;
				 l_2 = +17; end
		2637: begin l_1 = -6;
				 l_2 = -17; end
		3788: begin l_1 = +6;
				 l_2 = +18; end
		823: begin l_1 = +6;
				 l_2 = -18; end
		3724: begin l_1 = -6;
				 l_2 = +18; end
		759: begin l_1 = -6;
				 l_2 = -18; end
		2997: begin l_1 = +6;
				 l_2 = +19; end
		1614: begin l_1 = +6;
				 l_2 = -19; end
		2933: begin l_1 = -6;
				 l_2 = +19; end
		1550: begin l_1 = -6;
				 l_2 = -19; end
		1415: begin l_1 = +6;
				 l_2 = +20; end
		3196: begin l_1 = +6;
				 l_2 = -20; end
		1351: begin l_1 = -6;
				 l_2 = +20; end
		3132: begin l_1 = -6;
				 l_2 = -20; end
		2798: begin l_1 = +6;
				 l_2 = +21; end
		1813: begin l_1 = +6;
				 l_2 = -21; end
		2734: begin l_1 = -6;
				 l_2 = +21; end
		1749: begin l_1 = -6;
				 l_2 = -21; end
		1017: begin l_1 = +6;
				 l_2 = +22; end
		3594: begin l_1 = +6;
				 l_2 = -22; end
		953: begin l_1 = -6;
				 l_2 = +22; end
		3530: begin l_1 = -6;
				 l_2 = -22; end
		2002: begin l_1 = +6;
				 l_2 = +23; end
		2609: begin l_1 = +6;
				 l_2 = -23; end
		1938: begin l_1 = -6;
				 l_2 = +23; end
		2545: begin l_1 = -6;
				 l_2 = -23; end
		3972: begin l_1 = +6;
				 l_2 = +24; end
		639: begin l_1 = +6;
				 l_2 = -24; end
		3908: begin l_1 = -6;
				 l_2 = +24; end
		575: begin l_1 = -6;
				 l_2 = -24; end
		3365: begin l_1 = +6;
				 l_2 = +25; end
		1246: begin l_1 = +6;
				 l_2 = -25; end
		3301: begin l_1 = -6;
				 l_2 = +25; end
		1182: begin l_1 = -6;
				 l_2 = -25; end
		2151: begin l_1 = +6;
				 l_2 = +26; end
		2460: begin l_1 = +6;
				 l_2 = -26; end
		2087: begin l_1 = -6;
				 l_2 = +26; end
		2396: begin l_1 = -6;
				 l_2 = -26; end
		4270: begin l_1 = +6;
				 l_2 = +27; end
		341: begin l_1 = +6;
				 l_2 = -27; end
		4206: begin l_1 = -6;
				 l_2 = +27; end
		277: begin l_1 = -6;
				 l_2 = -27; end
		3961: begin l_1 = +6;
				 l_2 = +28; end
		650: begin l_1 = +6;
				 l_2 = -28; end
		3897: begin l_1 = -6;
				 l_2 = +28; end
		586: begin l_1 = -6;
				 l_2 = -28; end
		3343: begin l_1 = +6;
				 l_2 = +29; end
		1268: begin l_1 = +6;
				 l_2 = -29; end
		3279: begin l_1 = -6;
				 l_2 = +29; end
		1204: begin l_1 = -6;
				 l_2 = -29; end
		192: begin l_1 = -7;
				 l_2 = +9; end
		4355: begin l_1 = -7;
				 l_2 = -8; end
		320: begin l_1 = +7;
				 l_2 = +9; end
		4227: begin l_1 = -7;
				 l_2 = -9; end
		576: begin l_1 = +7;
				 l_2 = +10; end
		4099: begin l_1 = +7;
				 l_2 = -10; end
		448: begin l_1 = -7;
				 l_2 = +10; end
		3971: begin l_1 = -7;
				 l_2 = -10; end
		1088: begin l_1 = +7;
				 l_2 = +11; end
		3587: begin l_1 = +7;
				 l_2 = -11; end
		960: begin l_1 = -7;
				 l_2 = +11; end
		3459: begin l_1 = -7;
				 l_2 = -11; end
		2112: begin l_1 = +7;
				 l_2 = +12; end
		2563: begin l_1 = +7;
				 l_2 = -12; end
		1984: begin l_1 = -7;
				 l_2 = +12; end
		2435: begin l_1 = -7;
				 l_2 = -12; end
		4160: begin l_1 = +7;
				 l_2 = +13; end
		515: begin l_1 = +7;
				 l_2 = -13; end
		4032: begin l_1 = -7;
				 l_2 = +13; end
		387: begin l_1 = -7;
				 l_2 = -13; end
		3709: begin l_1 = +7;
				 l_2 = +14; end
		966: begin l_1 = +7;
				 l_2 = -14; end
		3581: begin l_1 = -7;
				 l_2 = +14; end
		838: begin l_1 = -7;
				 l_2 = -14; end
		2807: begin l_1 = +7;
				 l_2 = +15; end
		1868: begin l_1 = +7;
				 l_2 = -15; end
		2679: begin l_1 = -7;
				 l_2 = +15; end
		1740: begin l_1 = -7;
				 l_2 = -15; end
		1003: begin l_1 = +7;
				 l_2 = +16; end
		3672: begin l_1 = +7;
				 l_2 = -16; end
		875: begin l_1 = -7;
				 l_2 = +16; end
		3544: begin l_1 = -7;
				 l_2 = -16; end
		1942: begin l_1 = +7;
				 l_2 = +17; end
		2733: begin l_1 = +7;
				 l_2 = -17; end
		1814: begin l_1 = -7;
				 l_2 = +17; end
		2605: begin l_1 = -7;
				 l_2 = -17; end
		3820: begin l_1 = +7;
				 l_2 = +18; end
		855: begin l_1 = +7;
				 l_2 = -18; end
		3692: begin l_1 = -7;
				 l_2 = +18; end
		727: begin l_1 = -7;
				 l_2 = -18; end
		3029: begin l_1 = +7;
				 l_2 = +19; end
		1646: begin l_1 = +7;
				 l_2 = -19; end
		2901: begin l_1 = -7;
				 l_2 = +19; end
		1518: begin l_1 = -7;
				 l_2 = -19; end
		1447: begin l_1 = +7;
				 l_2 = +20; end
		3228: begin l_1 = +7;
				 l_2 = -20; end
		1319: begin l_1 = -7;
				 l_2 = +20; end
		3100: begin l_1 = -7;
				 l_2 = -20; end
		2830: begin l_1 = +7;
				 l_2 = +21; end
		1845: begin l_1 = +7;
				 l_2 = -21; end
		2702: begin l_1 = -7;
				 l_2 = +21; end
		1717: begin l_1 = -7;
				 l_2 = -21; end
		1049: begin l_1 = +7;
				 l_2 = +22; end
		3626: begin l_1 = +7;
				 l_2 = -22; end
		921: begin l_1 = -7;
				 l_2 = +22; end
		3498: begin l_1 = -7;
				 l_2 = -22; end
		2034: begin l_1 = +7;
				 l_2 = +23; end
		2641: begin l_1 = +7;
				 l_2 = -23; end
		1906: begin l_1 = -7;
				 l_2 = +23; end
		2513: begin l_1 = -7;
				 l_2 = -23; end
		4004: begin l_1 = +7;
				 l_2 = +24; end
		671: begin l_1 = +7;
				 l_2 = -24; end
		3876: begin l_1 = -7;
				 l_2 = +24; end
		543: begin l_1 = -7;
				 l_2 = -24; end
		3397: begin l_1 = +7;
				 l_2 = +25; end
		1278: begin l_1 = +7;
				 l_2 = -25; end
		3269: begin l_1 = -7;
				 l_2 = +25; end
		1150: begin l_1 = -7;
				 l_2 = -25; end
		2183: begin l_1 = +7;
				 l_2 = +26; end
		2492: begin l_1 = +7;
				 l_2 = -26; end
		2055: begin l_1 = -7;
				 l_2 = +26; end
		2364: begin l_1 = -7;
				 l_2 = -26; end
		4302: begin l_1 = +7;
				 l_2 = +27; end
		373: begin l_1 = +7;
				 l_2 = -27; end
		4174: begin l_1 = -7;
				 l_2 = +27; end
		245: begin l_1 = -7;
				 l_2 = -27; end
		3993: begin l_1 = +7;
				 l_2 = +28; end
		682: begin l_1 = +7;
				 l_2 = -28; end
		3865: begin l_1 = -7;
				 l_2 = +28; end
		554: begin l_1 = -7;
				 l_2 = -28; end
		3375: begin l_1 = +7;
				 l_2 = +29; end
		1300: begin l_1 = +7;
				 l_2 = -29; end
		3247: begin l_1 = -7;
				 l_2 = +29; end
		1172: begin l_1 = -7;
				 l_2 = -29; end
		384: begin l_1 = -8;
				 l_2 = +10; end
		4163: begin l_1 = -8;
				 l_2 = -9; end
		640: begin l_1 = +8;
				 l_2 = +10; end
		3907: begin l_1 = -8;
				 l_2 = -10; end
		1152: begin l_1 = +8;
				 l_2 = +11; end
		3651: begin l_1 = +8;
				 l_2 = -11; end
		896: begin l_1 = -8;
				 l_2 = +11; end
		3395: begin l_1 = -8;
				 l_2 = -11; end
		2176: begin l_1 = +8;
				 l_2 = +12; end
		2627: begin l_1 = +8;
				 l_2 = -12; end
		1920: begin l_1 = -8;
				 l_2 = +12; end
		2371: begin l_1 = -8;
				 l_2 = -12; end
		4224: begin l_1 = +8;
				 l_2 = +13; end
		579: begin l_1 = +8;
				 l_2 = -13; end
		3968: begin l_1 = -8;
				 l_2 = +13; end
		323: begin l_1 = -8;
				 l_2 = -13; end
		3773: begin l_1 = +8;
				 l_2 = +14; end
		1030: begin l_1 = +8;
				 l_2 = -14; end
		3517: begin l_1 = -8;
				 l_2 = +14; end
		774: begin l_1 = -8;
				 l_2 = -14; end
		2871: begin l_1 = +8;
				 l_2 = +15; end
		1932: begin l_1 = +8;
				 l_2 = -15; end
		2615: begin l_1 = -8;
				 l_2 = +15; end
		1676: begin l_1 = -8;
				 l_2 = -15; end
		1067: begin l_1 = +8;
				 l_2 = +16; end
		3736: begin l_1 = +8;
				 l_2 = -16; end
		811: begin l_1 = -8;
				 l_2 = +16; end
		3480: begin l_1 = -8;
				 l_2 = -16; end
		2006: begin l_1 = +8;
				 l_2 = +17; end
		2797: begin l_1 = +8;
				 l_2 = -17; end
		1750: begin l_1 = -8;
				 l_2 = +17; end
		2541: begin l_1 = -8;
				 l_2 = -17; end
		3884: begin l_1 = +8;
				 l_2 = +18; end
		919: begin l_1 = +8;
				 l_2 = -18; end
		3628: begin l_1 = -8;
				 l_2 = +18; end
		663: begin l_1 = -8;
				 l_2 = -18; end
		3093: begin l_1 = +8;
				 l_2 = +19; end
		1710: begin l_1 = +8;
				 l_2 = -19; end
		2837: begin l_1 = -8;
				 l_2 = +19; end
		1454: begin l_1 = -8;
				 l_2 = -19; end
		1511: begin l_1 = +8;
				 l_2 = +20; end
		3292: begin l_1 = +8;
				 l_2 = -20; end
		1255: begin l_1 = -8;
				 l_2 = +20; end
		3036: begin l_1 = -8;
				 l_2 = -20; end
		2894: begin l_1 = +8;
				 l_2 = +21; end
		1909: begin l_1 = +8;
				 l_2 = -21; end
		2638: begin l_1 = -8;
				 l_2 = +21; end
		1653: begin l_1 = -8;
				 l_2 = -21; end
		1113: begin l_1 = +8;
				 l_2 = +22; end
		3690: begin l_1 = +8;
				 l_2 = -22; end
		857: begin l_1 = -8;
				 l_2 = +22; end
		3434: begin l_1 = -8;
				 l_2 = -22; end
		2098: begin l_1 = +8;
				 l_2 = +23; end
		2705: begin l_1 = +8;
				 l_2 = -23; end
		1842: begin l_1 = -8;
				 l_2 = +23; end
		2449: begin l_1 = -8;
				 l_2 = -23; end
		4068: begin l_1 = +8;
				 l_2 = +24; end
		735: begin l_1 = +8;
				 l_2 = -24; end
		3812: begin l_1 = -8;
				 l_2 = +24; end
		479: begin l_1 = -8;
				 l_2 = -24; end
		3461: begin l_1 = +8;
				 l_2 = +25; end
		1342: begin l_1 = +8;
				 l_2 = -25; end
		3205: begin l_1 = -8;
				 l_2 = +25; end
		1086: begin l_1 = -8;
				 l_2 = -25; end
		2247: begin l_1 = +8;
				 l_2 = +26; end
		2556: begin l_1 = +8;
				 l_2 = -26; end
		1991: begin l_1 = -8;
				 l_2 = +26; end
		2300: begin l_1 = -8;
				 l_2 = -26; end
		4366: begin l_1 = +8;
				 l_2 = +27; end
		437: begin l_1 = +8;
				 l_2 = -27; end
		4110: begin l_1 = -8;
				 l_2 = +27; end
		181: begin l_1 = -8;
				 l_2 = -27; end
		4057: begin l_1 = +8;
				 l_2 = +28; end
		746: begin l_1 = +8;
				 l_2 = -28; end
		3801: begin l_1 = -8;
				 l_2 = +28; end
		490: begin l_1 = -8;
				 l_2 = -28; end
		3439: begin l_1 = +8;
				 l_2 = +29; end
		1364: begin l_1 = +8;
				 l_2 = -29; end
		3183: begin l_1 = -8;
				 l_2 = +29; end
		1108: begin l_1 = -8;
				 l_2 = -29; end
		768: begin l_1 = -9;
				 l_2 = +11; end
		3779: begin l_1 = -9;
				 l_2 = -10; end
		1280: begin l_1 = +9;
				 l_2 = +11; end
		3267: begin l_1 = -9;
				 l_2 = -11; end
		2304: begin l_1 = +9;
				 l_2 = +12; end
		2755: begin l_1 = +9;
				 l_2 = -12; end
		1792: begin l_1 = -9;
				 l_2 = +12; end
		2243: begin l_1 = -9;
				 l_2 = -12; end
		4352: begin l_1 = +9;
				 l_2 = +13; end
		707: begin l_1 = +9;
				 l_2 = -13; end
		3840: begin l_1 = -9;
				 l_2 = +13; end
		195: begin l_1 = -9;
				 l_2 = -13; end
		3901: begin l_1 = +9;
				 l_2 = +14; end
		1158: begin l_1 = +9;
				 l_2 = -14; end
		3389: begin l_1 = -9;
				 l_2 = +14; end
		646: begin l_1 = -9;
				 l_2 = -14; end
		2999: begin l_1 = +9;
				 l_2 = +15; end
		2060: begin l_1 = +9;
				 l_2 = -15; end
		2487: begin l_1 = -9;
				 l_2 = +15; end
		1548: begin l_1 = -9;
				 l_2 = -15; end
		1195: begin l_1 = +9;
				 l_2 = +16; end
		3864: begin l_1 = +9;
				 l_2 = -16; end
		683: begin l_1 = -9;
				 l_2 = +16; end
		3352: begin l_1 = -9;
				 l_2 = -16; end
		2134: begin l_1 = +9;
				 l_2 = +17; end
		2925: begin l_1 = +9;
				 l_2 = -17; end
		1622: begin l_1 = -9;
				 l_2 = +17; end
		2413: begin l_1 = -9;
				 l_2 = -17; end
		4012: begin l_1 = +9;
				 l_2 = +18; end
		1047: begin l_1 = +9;
				 l_2 = -18; end
		3500: begin l_1 = -9;
				 l_2 = +18; end
		535: begin l_1 = -9;
				 l_2 = -18; end
		3221: begin l_1 = +9;
				 l_2 = +19; end
		1838: begin l_1 = +9;
				 l_2 = -19; end
		2709: begin l_1 = -9;
				 l_2 = +19; end
		1326: begin l_1 = -9;
				 l_2 = -19; end
		1639: begin l_1 = +9;
				 l_2 = +20; end
		3420: begin l_1 = +9;
				 l_2 = -20; end
		1127: begin l_1 = -9;
				 l_2 = +20; end
		2908: begin l_1 = -9;
				 l_2 = -20; end
		3022: begin l_1 = +9;
				 l_2 = +21; end
		2037: begin l_1 = +9;
				 l_2 = -21; end
		2510: begin l_1 = -9;
				 l_2 = +21; end
		1525: begin l_1 = -9;
				 l_2 = -21; end
		1241: begin l_1 = +9;
				 l_2 = +22; end
		3818: begin l_1 = +9;
				 l_2 = -22; end
		729: begin l_1 = -9;
				 l_2 = +22; end
		3306: begin l_1 = -9;
				 l_2 = -22; end
		2226: begin l_1 = +9;
				 l_2 = +23; end
		2833: begin l_1 = +9;
				 l_2 = -23; end
		1714: begin l_1 = -9;
				 l_2 = +23; end
		2321: begin l_1 = -9;
				 l_2 = -23; end
		4196: begin l_1 = +9;
				 l_2 = +24; end
		863: begin l_1 = +9;
				 l_2 = -24; end
		3684: begin l_1 = -9;
				 l_2 = +24; end
		351: begin l_1 = -9;
				 l_2 = -24; end
		3589: begin l_1 = +9;
				 l_2 = +25; end
		1470: begin l_1 = +9;
				 l_2 = -25; end
		3077: begin l_1 = -9;
				 l_2 = +25; end
		958: begin l_1 = -9;
				 l_2 = -25; end
		2375: begin l_1 = +9;
				 l_2 = +26; end
		2684: begin l_1 = +9;
				 l_2 = -26; end
		1863: begin l_1 = -9;
				 l_2 = +26; end
		2172: begin l_1 = -9;
				 l_2 = -26; end
		4494: begin l_1 = +9;
				 l_2 = +27; end
		565: begin l_1 = +9;
				 l_2 = -27; end
		3982: begin l_1 = -9;
				 l_2 = +27; end
		53: begin l_1 = -9;
				 l_2 = -27; end
		4185: begin l_1 = +9;
				 l_2 = +28; end
		874: begin l_1 = +9;
				 l_2 = -28; end
		3673: begin l_1 = -9;
				 l_2 = +28; end
		362: begin l_1 = -9;
				 l_2 = -28; end
		3567: begin l_1 = +9;
				 l_2 = +29; end
		1492: begin l_1 = +9;
				 l_2 = -29; end
		3055: begin l_1 = -9;
				 l_2 = +29; end
		980: begin l_1 = -9;
				 l_2 = -29; end
		1536: begin l_1 = -10;
				 l_2 = +12; end
		3011: begin l_1 = -10;
				 l_2 = -11; end
		2560: begin l_1 = +10;
				 l_2 = +12; end
		1987: begin l_1 = -10;
				 l_2 = -12; end
		61: begin l_1 = +10;
				 l_2 = +13; end
		963: begin l_1 = +10;
				 l_2 = -13; end
		3584: begin l_1 = -10;
				 l_2 = +13; end
		4486: begin l_1 = -10;
				 l_2 = -13; end
		4157: begin l_1 = +10;
				 l_2 = +14; end
		1414: begin l_1 = +10;
				 l_2 = -14; end
		3133: begin l_1 = -10;
				 l_2 = +14; end
		390: begin l_1 = -10;
				 l_2 = -14; end
		3255: begin l_1 = +10;
				 l_2 = +15; end
		2316: begin l_1 = +10;
				 l_2 = -15; end
		2231: begin l_1 = -10;
				 l_2 = +15; end
		1292: begin l_1 = -10;
				 l_2 = -15; end
		1451: begin l_1 = +10;
				 l_2 = +16; end
		4120: begin l_1 = +10;
				 l_2 = -16; end
		427: begin l_1 = -10;
				 l_2 = +16; end
		3096: begin l_1 = -10;
				 l_2 = -16; end
		2390: begin l_1 = +10;
				 l_2 = +17; end
		3181: begin l_1 = +10;
				 l_2 = -17; end
		1366: begin l_1 = -10;
				 l_2 = +17; end
		2157: begin l_1 = -10;
				 l_2 = -17; end
		4268: begin l_1 = +10;
				 l_2 = +18; end
		1303: begin l_1 = +10;
				 l_2 = -18; end
		3244: begin l_1 = -10;
				 l_2 = +18; end
		279: begin l_1 = -10;
				 l_2 = -18; end
		3477: begin l_1 = +10;
				 l_2 = +19; end
		2094: begin l_1 = +10;
				 l_2 = -19; end
		2453: begin l_1 = -10;
				 l_2 = +19; end
		1070: begin l_1 = -10;
				 l_2 = -19; end
		1895: begin l_1 = +10;
				 l_2 = +20; end
		3676: begin l_1 = +10;
				 l_2 = -20; end
		871: begin l_1 = -10;
				 l_2 = +20; end
		2652: begin l_1 = -10;
				 l_2 = -20; end
		3278: begin l_1 = +10;
				 l_2 = +21; end
		2293: begin l_1 = +10;
				 l_2 = -21; end
		2254: begin l_1 = -10;
				 l_2 = +21; end
		1269: begin l_1 = -10;
				 l_2 = -21; end
		1497: begin l_1 = +10;
				 l_2 = +22; end
		4074: begin l_1 = +10;
				 l_2 = -22; end
		473: begin l_1 = -10;
				 l_2 = +22; end
		3050: begin l_1 = -10;
				 l_2 = -22; end
		2482: begin l_1 = +10;
				 l_2 = +23; end
		3089: begin l_1 = +10;
				 l_2 = -23; end
		1458: begin l_1 = -10;
				 l_2 = +23; end
		2065: begin l_1 = -10;
				 l_2 = -23; end
		4452: begin l_1 = +10;
				 l_2 = +24; end
		1119: begin l_1 = +10;
				 l_2 = -24; end
		3428: begin l_1 = -10;
				 l_2 = +24; end
		95: begin l_1 = -10;
				 l_2 = -24; end
		3845: begin l_1 = +10;
				 l_2 = +25; end
		1726: begin l_1 = +10;
				 l_2 = -25; end
		2821: begin l_1 = -10;
				 l_2 = +25; end
		702: begin l_1 = -10;
				 l_2 = -25; end
		2631: begin l_1 = +10;
				 l_2 = +26; end
		2940: begin l_1 = +10;
				 l_2 = -26; end
		1607: begin l_1 = -10;
				 l_2 = +26; end
		1916: begin l_1 = -10;
				 l_2 = -26; end
		203: begin l_1 = +10;
				 l_2 = +27; end
		821: begin l_1 = +10;
				 l_2 = -27; end
		3726: begin l_1 = -10;
				 l_2 = +27; end
		4344: begin l_1 = -10;
				 l_2 = -27; end
		4441: begin l_1 = +10;
				 l_2 = +28; end
		1130: begin l_1 = +10;
				 l_2 = -28; end
		3417: begin l_1 = -10;
				 l_2 = +28; end
		106: begin l_1 = -10;
				 l_2 = -28; end
		3823: begin l_1 = +10;
				 l_2 = +29; end
		1748: begin l_1 = +10;
				 l_2 = -29; end
		2799: begin l_1 = -10;
				 l_2 = +29; end
		724: begin l_1 = -10;
				 l_2 = -29; end
		3072: begin l_1 = -11;
				 l_2 = +13; end
		1475: begin l_1 = -11;
				 l_2 = -12; end
		573: begin l_1 = +11;
				 l_2 = +13; end
		3974: begin l_1 = -11;
				 l_2 = -13; end
		122: begin l_1 = +11;
				 l_2 = +14; end
		1926: begin l_1 = +11;
				 l_2 = -14; end
		2621: begin l_1 = -11;
				 l_2 = +14; end
		4425: begin l_1 = -11;
				 l_2 = -14; end
		3767: begin l_1 = +11;
				 l_2 = +15; end
		2828: begin l_1 = +11;
				 l_2 = -15; end
		1719: begin l_1 = -11;
				 l_2 = +15; end
		780: begin l_1 = -11;
				 l_2 = -15; end
		1963: begin l_1 = +11;
				 l_2 = +16; end
		85: begin l_1 = +11;
				 l_2 = -16; end
		4462: begin l_1 = -11;
				 l_2 = +16; end
		2584: begin l_1 = -11;
				 l_2 = -16; end
		2902: begin l_1 = +11;
				 l_2 = +17; end
		3693: begin l_1 = +11;
				 l_2 = -17; end
		854: begin l_1 = -11;
				 l_2 = +17; end
		1645: begin l_1 = -11;
				 l_2 = -17; end
		233: begin l_1 = +11;
				 l_2 = +18; end
		1815: begin l_1 = +11;
				 l_2 = -18; end
		2732: begin l_1 = -11;
				 l_2 = +18; end
		4314: begin l_1 = -11;
				 l_2 = -18; end
		3989: begin l_1 = +11;
				 l_2 = +19; end
		2606: begin l_1 = +11;
				 l_2 = -19; end
		1941: begin l_1 = -11;
				 l_2 = +19; end
		558: begin l_1 = -11;
				 l_2 = -19; end
		2407: begin l_1 = +11;
				 l_2 = +20; end
		4188: begin l_1 = +11;
				 l_2 = -20; end
		359: begin l_1 = -11;
				 l_2 = +20; end
		2140: begin l_1 = -11;
				 l_2 = -20; end
		3790: begin l_1 = +11;
				 l_2 = +21; end
		2805: begin l_1 = +11;
				 l_2 = -21; end
		1742: begin l_1 = -11;
				 l_2 = +21; end
		757: begin l_1 = -11;
				 l_2 = -21; end
		2009: begin l_1 = +11;
				 l_2 = +22; end
		39: begin l_1 = +11;
				 l_2 = -22; end
		4508: begin l_1 = -11;
				 l_2 = +22; end
		2538: begin l_1 = -11;
				 l_2 = -22; end
		2994: begin l_1 = +11;
				 l_2 = +23; end
		3601: begin l_1 = +11;
				 l_2 = -23; end
		946: begin l_1 = -11;
				 l_2 = +23; end
		1553: begin l_1 = -11;
				 l_2 = -23; end
		417: begin l_1 = +11;
				 l_2 = +24; end
		1631: begin l_1 = +11;
				 l_2 = -24; end
		2916: begin l_1 = -11;
				 l_2 = +24; end
		4130: begin l_1 = -11;
				 l_2 = -24; end
		4357: begin l_1 = +11;
				 l_2 = +25; end
		2238: begin l_1 = +11;
				 l_2 = -25; end
		2309: begin l_1 = -11;
				 l_2 = +25; end
		190: begin l_1 = -11;
				 l_2 = -25; end
		3143: begin l_1 = +11;
				 l_2 = +26; end
		3452: begin l_1 = +11;
				 l_2 = -26; end
		1095: begin l_1 = -11;
				 l_2 = +26; end
		1404: begin l_1 = -11;
				 l_2 = -26; end
		715: begin l_1 = +11;
				 l_2 = +27; end
		1333: begin l_1 = +11;
				 l_2 = -27; end
		3214: begin l_1 = -11;
				 l_2 = +27; end
		3832: begin l_1 = -11;
				 l_2 = -27; end
		406: begin l_1 = +11;
				 l_2 = +28; end
		1642: begin l_1 = +11;
				 l_2 = -28; end
		2905: begin l_1 = -11;
				 l_2 = +28; end
		4141: begin l_1 = -11;
				 l_2 = -28; end
		4335: begin l_1 = +11;
				 l_2 = +29; end
		2260: begin l_1 = +11;
				 l_2 = -29; end
		2287: begin l_1 = -11;
				 l_2 = +29; end
		212: begin l_1 = -11;
				 l_2 = -29; end
		1597: begin l_1 = -12;
				 l_2 = +14; end
		2950: begin l_1 = -12;
				 l_2 = -13; end
		1146: begin l_1 = +12;
				 l_2 = +14; end
		3401: begin l_1 = -12;
				 l_2 = -14; end
		244: begin l_1 = +12;
				 l_2 = +15; end
		3852: begin l_1 = +12;
				 l_2 = -15; end
		695: begin l_1 = -12;
				 l_2 = +15; end
		4303: begin l_1 = -12;
				 l_2 = -15; end
		2987: begin l_1 = +12;
				 l_2 = +16; end
		1109: begin l_1 = +12;
				 l_2 = -16; end
		3438: begin l_1 = -12;
				 l_2 = +16; end
		1560: begin l_1 = -12;
				 l_2 = -16; end
		3926: begin l_1 = +12;
				 l_2 = +17; end
		170: begin l_1 = +12;
				 l_2 = -17; end
		4377: begin l_1 = -12;
				 l_2 = +17; end
		621: begin l_1 = -12;
				 l_2 = -17; end
		1257: begin l_1 = +12;
				 l_2 = +18; end
		2839: begin l_1 = +12;
				 l_2 = -18; end
		1708: begin l_1 = -12;
				 l_2 = +18; end
		3290: begin l_1 = -12;
				 l_2 = -18; end
		466: begin l_1 = +12;
				 l_2 = +19; end
		3630: begin l_1 = +12;
				 l_2 = -19; end
		917: begin l_1 = -12;
				 l_2 = +19; end
		4081: begin l_1 = -12;
				 l_2 = -19; end
		3431: begin l_1 = +12;
				 l_2 = +20; end
		665: begin l_1 = +12;
				 l_2 = -20; end
		3882: begin l_1 = -12;
				 l_2 = +20; end
		1116: begin l_1 = -12;
				 l_2 = -20; end
		267: begin l_1 = +12;
				 l_2 = +21; end
		3829: begin l_1 = +12;
				 l_2 = -21; end
		718: begin l_1 = -12;
				 l_2 = +21; end
		4280: begin l_1 = -12;
				 l_2 = -21; end
		3033: begin l_1 = +12;
				 l_2 = +22; end
		1063: begin l_1 = +12;
				 l_2 = -22; end
		3484: begin l_1 = -12;
				 l_2 = +22; end
		1514: begin l_1 = -12;
				 l_2 = -22; end
		4018: begin l_1 = +12;
				 l_2 = +23; end
		78: begin l_1 = +12;
				 l_2 = -23; end
		4469: begin l_1 = -12;
				 l_2 = +23; end
		529: begin l_1 = -12;
				 l_2 = -23; end
		1441: begin l_1 = +12;
				 l_2 = +24; end
		2655: begin l_1 = +12;
				 l_2 = -24; end
		1892: begin l_1 = -12;
				 l_2 = +24; end
		3106: begin l_1 = -12;
				 l_2 = -24; end
		834: begin l_1 = +12;
				 l_2 = +25; end
		3262: begin l_1 = +12;
				 l_2 = -25; end
		1285: begin l_1 = -12;
				 l_2 = +25; end
		3713: begin l_1 = -12;
				 l_2 = -25; end
		4167: begin l_1 = +12;
				 l_2 = +26; end
		4476: begin l_1 = +12;
				 l_2 = -26; end
		71: begin l_1 = -12;
				 l_2 = +26; end
		380: begin l_1 = -12;
				 l_2 = -26; end
		1739: begin l_1 = +12;
				 l_2 = +27; end
		2357: begin l_1 = +12;
				 l_2 = -27; end
		2190: begin l_1 = -12;
				 l_2 = +27; end
		2808: begin l_1 = -12;
				 l_2 = -27; end
		1430: begin l_1 = +12;
				 l_2 = +28; end
		2666: begin l_1 = +12;
				 l_2 = -28; end
		1881: begin l_1 = -12;
				 l_2 = +28; end
		3117: begin l_1 = -12;
				 l_2 = -28; end
		812: begin l_1 = +12;
				 l_2 = +29; end
		3284: begin l_1 = +12;
				 l_2 = -29; end
		1263: begin l_1 = -12;
				 l_2 = +29; end
		3735: begin l_1 = -12;
				 l_2 = -29; end
		3194: begin l_1 = -13;
				 l_2 = +15; end
		1353: begin l_1 = -13;
				 l_2 = -14; end
		2292: begin l_1 = +13;
				 l_2 = +15; end
		2255: begin l_1 = -13;
				 l_2 = -15; end
		488: begin l_1 = +13;
				 l_2 = +16; end
		3157: begin l_1 = +13;
				 l_2 = -16; end
		1390: begin l_1 = -13;
				 l_2 = +16; end
		4059: begin l_1 = -13;
				 l_2 = -16; end
		1427: begin l_1 = +13;
				 l_2 = +17; end
		2218: begin l_1 = +13;
				 l_2 = -17; end
		2329: begin l_1 = -13;
				 l_2 = +17; end
		3120: begin l_1 = -13;
				 l_2 = -17; end
		3305: begin l_1 = +13;
				 l_2 = +18; end
		340: begin l_1 = +13;
				 l_2 = -18; end
		4207: begin l_1 = -13;
				 l_2 = +18; end
		1242: begin l_1 = -13;
				 l_2 = -18; end
		2514: begin l_1 = +13;
				 l_2 = +19; end
		1131: begin l_1 = +13;
				 l_2 = -19; end
		3416: begin l_1 = -13;
				 l_2 = +19; end
		2033: begin l_1 = -13;
				 l_2 = -19; end
		932: begin l_1 = +13;
				 l_2 = +20; end
		2713: begin l_1 = +13;
				 l_2 = -20; end
		1834: begin l_1 = -13;
				 l_2 = +20; end
		3615: begin l_1 = -13;
				 l_2 = -20; end
		2315: begin l_1 = +13;
				 l_2 = +21; end
		1330: begin l_1 = +13;
				 l_2 = -21; end
		3217: begin l_1 = -13;
				 l_2 = +21; end
		2232: begin l_1 = -13;
				 l_2 = -21; end
		534: begin l_1 = +13;
				 l_2 = +22; end
		3111: begin l_1 = +13;
				 l_2 = -22; end
		1436: begin l_1 = -13;
				 l_2 = +22; end
		4013: begin l_1 = -13;
				 l_2 = -22; end
		1519: begin l_1 = +13;
				 l_2 = +23; end
		2126: begin l_1 = +13;
				 l_2 = -23; end
		2421: begin l_1 = -13;
				 l_2 = +23; end
		3028: begin l_1 = -13;
				 l_2 = -23; end
		3489: begin l_1 = +13;
				 l_2 = +24; end
		156: begin l_1 = +13;
				 l_2 = -24; end
		4391: begin l_1 = -13;
				 l_2 = +24; end
		1058: begin l_1 = -13;
				 l_2 = -24; end
		2882: begin l_1 = +13;
				 l_2 = +25; end
		763: begin l_1 = +13;
				 l_2 = -25; end
		3784: begin l_1 = -13;
				 l_2 = +25; end
		1665: begin l_1 = -13;
				 l_2 = -25; end
		1668: begin l_1 = +13;
				 l_2 = +26; end
		1977: begin l_1 = +13;
				 l_2 = -26; end
		2570: begin l_1 = -13;
				 l_2 = +26; end
		2879: begin l_1 = -13;
				 l_2 = -26; end
		3787: begin l_1 = +13;
				 l_2 = +27; end
		4405: begin l_1 = +13;
				 l_2 = -27; end
		142: begin l_1 = -13;
				 l_2 = +27; end
		760: begin l_1 = -13;
				 l_2 = -27; end
		3478: begin l_1 = +13;
				 l_2 = +28; end
		167: begin l_1 = +13;
				 l_2 = -28; end
		4380: begin l_1 = -13;
				 l_2 = +28; end
		1069: begin l_1 = -13;
				 l_2 = -28; end
		2860: begin l_1 = +13;
				 l_2 = +29; end
		785: begin l_1 = +13;
				 l_2 = -29; end
		3762: begin l_1 = -13;
				 l_2 = +29; end
		1687: begin l_1 = -13;
				 l_2 = -29; end
		1841: begin l_1 = -14;
				 l_2 = +16; end
		2706: begin l_1 = -14;
				 l_2 = -15; end
		37: begin l_1 = +14;
				 l_2 = +16; end
		4510: begin l_1 = -14;
				 l_2 = -16; end
		976: begin l_1 = +14;
				 l_2 = +17; end
		1767: begin l_1 = +14;
				 l_2 = -17; end
		2780: begin l_1 = -14;
				 l_2 = +17; end
		3571: begin l_1 = -14;
				 l_2 = -17; end
		2854: begin l_1 = +14;
				 l_2 = +18; end
		4436: begin l_1 = +14;
				 l_2 = -18; end
		111: begin l_1 = -14;
				 l_2 = +18; end
		1693: begin l_1 = -14;
				 l_2 = -18; end
		2063: begin l_1 = +14;
				 l_2 = +19; end
		680: begin l_1 = +14;
				 l_2 = -19; end
		3867: begin l_1 = -14;
				 l_2 = +19; end
		2484: begin l_1 = -14;
				 l_2 = -19; end
		481: begin l_1 = +14;
				 l_2 = +20; end
		2262: begin l_1 = +14;
				 l_2 = -20; end
		2285: begin l_1 = -14;
				 l_2 = +20; end
		4066: begin l_1 = -14;
				 l_2 = -20; end
		1864: begin l_1 = +14;
				 l_2 = +21; end
		879: begin l_1 = +14;
				 l_2 = -21; end
		3668: begin l_1 = -14;
				 l_2 = +21; end
		2683: begin l_1 = -14;
				 l_2 = -21; end
		83: begin l_1 = +14;
				 l_2 = +22; end
		2660: begin l_1 = +14;
				 l_2 = -22; end
		1887: begin l_1 = -14;
				 l_2 = +22; end
		4464: begin l_1 = -14;
				 l_2 = -22; end
		1068: begin l_1 = +14;
				 l_2 = +23; end
		1675: begin l_1 = +14;
				 l_2 = -23; end
		2872: begin l_1 = -14;
				 l_2 = +23; end
		3479: begin l_1 = -14;
				 l_2 = -23; end
		3038: begin l_1 = +14;
				 l_2 = +24; end
		4252: begin l_1 = +14;
				 l_2 = -24; end
		295: begin l_1 = -14;
				 l_2 = +24; end
		1509: begin l_1 = -14;
				 l_2 = -24; end
		2431: begin l_1 = +14;
				 l_2 = +25; end
		312: begin l_1 = +14;
				 l_2 = -25; end
		4235: begin l_1 = -14;
				 l_2 = +25; end
		2116: begin l_1 = -14;
				 l_2 = -25; end
		1217: begin l_1 = +14;
				 l_2 = +26; end
		1526: begin l_1 = +14;
				 l_2 = -26; end
		3021: begin l_1 = -14;
				 l_2 = +26; end
		3330: begin l_1 = -14;
				 l_2 = -26; end
		3336: begin l_1 = +14;
				 l_2 = +27; end
		3954: begin l_1 = +14;
				 l_2 = -27; end
		593: begin l_1 = -14;
				 l_2 = +27; end
		1211: begin l_1 = -14;
				 l_2 = -27; end
		3027: begin l_1 = +14;
				 l_2 = +28; end
		4263: begin l_1 = +14;
				 l_2 = -28; end
		284: begin l_1 = -14;
				 l_2 = +28; end
		1520: begin l_1 = -14;
				 l_2 = -28; end
		2409: begin l_1 = +14;
				 l_2 = +29; end
		334: begin l_1 = +14;
				 l_2 = -29; end
		4213: begin l_1 = -14;
				 l_2 = +29; end
		2138: begin l_1 = -14;
				 l_2 = -29; end
		3682: begin l_1 = -15;
				 l_2 = +17; end
		865: begin l_1 = -15;
				 l_2 = -16; end
		74: begin l_1 = +15;
				 l_2 = +17; end
		4473: begin l_1 = -15;
				 l_2 = -17; end
		1952: begin l_1 = +15;
				 l_2 = +18; end
		3534: begin l_1 = +15;
				 l_2 = -18; end
		1013: begin l_1 = -15;
				 l_2 = +18; end
		2595: begin l_1 = -15;
				 l_2 = -18; end
		1161: begin l_1 = +15;
				 l_2 = +19; end
		4325: begin l_1 = +15;
				 l_2 = -19; end
		222: begin l_1 = -15;
				 l_2 = +19; end
		3386: begin l_1 = -15;
				 l_2 = -19; end
		4126: begin l_1 = +15;
				 l_2 = +20; end
		1360: begin l_1 = +15;
				 l_2 = -20; end
		3187: begin l_1 = -15;
				 l_2 = +20; end
		421: begin l_1 = -15;
				 l_2 = -20; end
		962: begin l_1 = +15;
				 l_2 = +21; end
		4524: begin l_1 = +15;
				 l_2 = -21; end
		23: begin l_1 = -15;
				 l_2 = +21; end
		3585: begin l_1 = -15;
				 l_2 = -21; end
		3728: begin l_1 = +15;
				 l_2 = +22; end
		1758: begin l_1 = +15;
				 l_2 = -22; end
		2789: begin l_1 = -15;
				 l_2 = +22; end
		819: begin l_1 = -15;
				 l_2 = -22; end
		166: begin l_1 = +15;
				 l_2 = +23; end
		773: begin l_1 = +15;
				 l_2 = -23; end
		3774: begin l_1 = -15;
				 l_2 = +23; end
		4381: begin l_1 = -15;
				 l_2 = -23; end
		2136: begin l_1 = +15;
				 l_2 = +24; end
		3350: begin l_1 = +15;
				 l_2 = -24; end
		1197: begin l_1 = -15;
				 l_2 = +24; end
		2411: begin l_1 = -15;
				 l_2 = -24; end
		1529: begin l_1 = +15;
				 l_2 = +25; end
		3957: begin l_1 = +15;
				 l_2 = -25; end
		590: begin l_1 = -15;
				 l_2 = +25; end
		3018: begin l_1 = -15;
				 l_2 = -25; end
		315: begin l_1 = +15;
				 l_2 = +26; end
		624: begin l_1 = +15;
				 l_2 = -26; end
		3923: begin l_1 = -15;
				 l_2 = +26; end
		4232: begin l_1 = -15;
				 l_2 = -26; end
		2434: begin l_1 = +15;
				 l_2 = +27; end
		3052: begin l_1 = +15;
				 l_2 = -27; end
		1495: begin l_1 = -15;
				 l_2 = +27; end
		2113: begin l_1 = -15;
				 l_2 = -27; end
		2125: begin l_1 = +15;
				 l_2 = +28; end
		3361: begin l_1 = +15;
				 l_2 = -28; end
		1186: begin l_1 = -15;
				 l_2 = +28; end
		2422: begin l_1 = -15;
				 l_2 = -28; end
		1507: begin l_1 = +15;
				 l_2 = +29; end
		3979: begin l_1 = +15;
				 l_2 = -29; end
		568: begin l_1 = -15;
				 l_2 = +29; end
		3040: begin l_1 = -15;
				 l_2 = -29; end
		2817: begin l_1 = -16;
				 l_2 = +18; end
		1730: begin l_1 = -16;
				 l_2 = -17; end
		148: begin l_1 = +16;
				 l_2 = +18; end
		4399: begin l_1 = -16;
				 l_2 = -18; end
		3904: begin l_1 = +16;
				 l_2 = +19; end
		2521: begin l_1 = +16;
				 l_2 = -19; end
		2026: begin l_1 = -16;
				 l_2 = +19; end
		643: begin l_1 = -16;
				 l_2 = -19; end
		2322: begin l_1 = +16;
				 l_2 = +20; end
		4103: begin l_1 = +16;
				 l_2 = -20; end
		444: begin l_1 = -16;
				 l_2 = +20; end
		2225: begin l_1 = -16;
				 l_2 = -20; end
		3705: begin l_1 = +16;
				 l_2 = +21; end
		2720: begin l_1 = +16;
				 l_2 = -21; end
		1827: begin l_1 = -16;
				 l_2 = +21; end
		842: begin l_1 = -16;
				 l_2 = -21; end
		1924: begin l_1 = +16;
				 l_2 = +22; end
		4501: begin l_1 = +16;
				 l_2 = -22; end
		46: begin l_1 = -16;
				 l_2 = +22; end
		2623: begin l_1 = -16;
				 l_2 = -22; end
		2909: begin l_1 = +16;
				 l_2 = +23; end
		3516: begin l_1 = +16;
				 l_2 = -23; end
		1031: begin l_1 = -16;
				 l_2 = +23; end
		1638: begin l_1 = -16;
				 l_2 = -23; end
		332: begin l_1 = +16;
				 l_2 = +24; end
		1546: begin l_1 = +16;
				 l_2 = -24; end
		3001: begin l_1 = -16;
				 l_2 = +24; end
		4215: begin l_1 = -16;
				 l_2 = -24; end
		4272: begin l_1 = +16;
				 l_2 = +25; end
		2153: begin l_1 = +16;
				 l_2 = -25; end
		2394: begin l_1 = -16;
				 l_2 = +25; end
		275: begin l_1 = -16;
				 l_2 = -25; end
		3058: begin l_1 = +16;
				 l_2 = +26; end
		3367: begin l_1 = +16;
				 l_2 = -26; end
		1180: begin l_1 = -16;
				 l_2 = +26; end
		1489: begin l_1 = -16;
				 l_2 = -26; end
		630: begin l_1 = +16;
				 l_2 = +27; end
		1248: begin l_1 = +16;
				 l_2 = -27; end
		3299: begin l_1 = -16;
				 l_2 = +27; end
		3917: begin l_1 = -16;
				 l_2 = -27; end
		321: begin l_1 = +16;
				 l_2 = +28; end
		1557: begin l_1 = +16;
				 l_2 = -28; end
		2990: begin l_1 = -16;
				 l_2 = +28; end
		4226: begin l_1 = -16;
				 l_2 = -28; end
		4250: begin l_1 = +16;
				 l_2 = +29; end
		2175: begin l_1 = +16;
				 l_2 = -29; end
		2372: begin l_1 = -16;
				 l_2 = +29; end
		297: begin l_1 = -16;
				 l_2 = -29; end
		1087: begin l_1 = -17;
				 l_2 = +19; end
		3460: begin l_1 = -17;
				 l_2 = -18; end
		296: begin l_1 = +17;
				 l_2 = +19; end
		4251: begin l_1 = -17;
				 l_2 = -19; end
		3261: begin l_1 = +17;
				 l_2 = +20; end
		495: begin l_1 = +17;
				 l_2 = -20; end
		4052: begin l_1 = -17;
				 l_2 = +20; end
		1286: begin l_1 = -17;
				 l_2 = -20; end
		97: begin l_1 = +17;
				 l_2 = +21; end
		3659: begin l_1 = +17;
				 l_2 = -21; end
		888: begin l_1 = -17;
				 l_2 = +21; end
		4450: begin l_1 = -17;
				 l_2 = -21; end
		2863: begin l_1 = +17;
				 l_2 = +22; end
		893: begin l_1 = +17;
				 l_2 = -22; end
		3654: begin l_1 = -17;
				 l_2 = +22; end
		1684: begin l_1 = -17;
				 l_2 = -22; end
		3848: begin l_1 = +17;
				 l_2 = +23; end
		4455: begin l_1 = +17;
				 l_2 = -23; end
		92: begin l_1 = -17;
				 l_2 = +23; end
		699: begin l_1 = -17;
				 l_2 = -23; end
		1271: begin l_1 = +17;
				 l_2 = +24; end
		2485: begin l_1 = +17;
				 l_2 = -24; end
		2062: begin l_1 = -17;
				 l_2 = +24; end
		3276: begin l_1 = -17;
				 l_2 = -24; end
		664: begin l_1 = +17;
				 l_2 = +25; end
		3092: begin l_1 = +17;
				 l_2 = -25; end
		1455: begin l_1 = -17;
				 l_2 = +25; end
		3883: begin l_1 = -17;
				 l_2 = -25; end
		3997: begin l_1 = +17;
				 l_2 = +26; end
		4306: begin l_1 = +17;
				 l_2 = -26; end
		241: begin l_1 = -17;
				 l_2 = +26; end
		550: begin l_1 = -17;
				 l_2 = -26; end
		1569: begin l_1 = +17;
				 l_2 = +27; end
		2187: begin l_1 = +17;
				 l_2 = -27; end
		2360: begin l_1 = -17;
				 l_2 = +27; end
		2978: begin l_1 = -17;
				 l_2 = -27; end
		1260: begin l_1 = +17;
				 l_2 = +28; end
		2496: begin l_1 = +17;
				 l_2 = -28; end
		2051: begin l_1 = -17;
				 l_2 = +28; end
		3287: begin l_1 = -17;
				 l_2 = -28; end
		642: begin l_1 = +17;
				 l_2 = +29; end
		3114: begin l_1 = +17;
				 l_2 = -29; end
		1433: begin l_1 = -17;
				 l_2 = +29; end
		3905: begin l_1 = -17;
				 l_2 = -29; end
		2174: begin l_1 = -18;
				 l_2 = +20; end
		2373: begin l_1 = -18;
				 l_2 = -19; end
		592: begin l_1 = +18;
				 l_2 = +20; end
		3955: begin l_1 = -18;
				 l_2 = -20; end
		1975: begin l_1 = +18;
				 l_2 = +21; end
		990: begin l_1 = +18;
				 l_2 = -21; end
		3557: begin l_1 = -18;
				 l_2 = +21; end
		2572: begin l_1 = -18;
				 l_2 = -21; end
		194: begin l_1 = +18;
				 l_2 = +22; end
		2771: begin l_1 = +18;
				 l_2 = -22; end
		1776: begin l_1 = -18;
				 l_2 = +22; end
		4353: begin l_1 = -18;
				 l_2 = -22; end
		1179: begin l_1 = +18;
				 l_2 = +23; end
		1786: begin l_1 = +18;
				 l_2 = -23; end
		2761: begin l_1 = -18;
				 l_2 = +23; end
		3368: begin l_1 = -18;
				 l_2 = -23; end
		3149: begin l_1 = +18;
				 l_2 = +24; end
		4363: begin l_1 = +18;
				 l_2 = -24; end
		184: begin l_1 = -18;
				 l_2 = +24; end
		1398: begin l_1 = -18;
				 l_2 = -24; end
		2542: begin l_1 = +18;
				 l_2 = +25; end
		423: begin l_1 = +18;
				 l_2 = -25; end
		4124: begin l_1 = -18;
				 l_2 = +25; end
		2005: begin l_1 = -18;
				 l_2 = -25; end
		1328: begin l_1 = +18;
				 l_2 = +26; end
		1637: begin l_1 = +18;
				 l_2 = -26; end
		2910: begin l_1 = -18;
				 l_2 = +26; end
		3219: begin l_1 = -18;
				 l_2 = -26; end
		3447: begin l_1 = +18;
				 l_2 = +27; end
		4065: begin l_1 = +18;
				 l_2 = -27; end
		482: begin l_1 = -18;
				 l_2 = +27; end
		1100: begin l_1 = -18;
				 l_2 = -27; end
		3138: begin l_1 = +18;
				 l_2 = +28; end
		4374: begin l_1 = +18;
				 l_2 = -28; end
		173: begin l_1 = -18;
				 l_2 = +28; end
		1409: begin l_1 = -18;
				 l_2 = -28; end
		2520: begin l_1 = +18;
				 l_2 = +29; end
		445: begin l_1 = +18;
				 l_2 = -29; end
		4102: begin l_1 = -18;
				 l_2 = +29; end
		2027: begin l_1 = -18;
				 l_2 = -29; end
		4348: begin l_1 = -19;
				 l_2 = +21; end
		199: begin l_1 = -19;
				 l_2 = -20; end
		1184: begin l_1 = +19;
				 l_2 = +21; end
		3363: begin l_1 = -19;
				 l_2 = -21; end
		3950: begin l_1 = +19;
				 l_2 = +22; end
		1980: begin l_1 = +19;
				 l_2 = -22; end
		2567: begin l_1 = -19;
				 l_2 = +22; end
		597: begin l_1 = -19;
				 l_2 = -22; end
		388: begin l_1 = +19;
				 l_2 = +23; end
		995: begin l_1 = +19;
				 l_2 = -23; end
		3552: begin l_1 = -19;
				 l_2 = +23; end
		4159: begin l_1 = -19;
				 l_2 = -23; end
		2358: begin l_1 = +19;
				 l_2 = +24; end
		3572: begin l_1 = +19;
				 l_2 = -24; end
		975: begin l_1 = -19;
				 l_2 = +24; end
		2189: begin l_1 = -19;
				 l_2 = -24; end
		1751: begin l_1 = +19;
				 l_2 = +25; end
		4179: begin l_1 = +19;
				 l_2 = -25; end
		368: begin l_1 = -19;
				 l_2 = +25; end
		2796: begin l_1 = -19;
				 l_2 = -25; end
		537: begin l_1 = +19;
				 l_2 = +26; end
		846: begin l_1 = +19;
				 l_2 = -26; end
		3701: begin l_1 = -19;
				 l_2 = +26; end
		4010: begin l_1 = -19;
				 l_2 = -26; end
		2656: begin l_1 = +19;
				 l_2 = +27; end
		3274: begin l_1 = +19;
				 l_2 = -27; end
		1273: begin l_1 = -19;
				 l_2 = +27; end
		1891: begin l_1 = -19;
				 l_2 = -27; end
		2347: begin l_1 = +19;
				 l_2 = +28; end
		3583: begin l_1 = +19;
				 l_2 = -28; end
		964: begin l_1 = -19;
				 l_2 = +28; end
		2200: begin l_1 = -19;
				 l_2 = -28; end
		1729: begin l_1 = +19;
				 l_2 = +29; end
		4201: begin l_1 = +19;
				 l_2 = -29; end
		346: begin l_1 = -19;
				 l_2 = +29; end
		2818: begin l_1 = -19;
				 l_2 = -29; end
		4149: begin l_1 = -20;
				 l_2 = +22; end
		398: begin l_1 = -20;
				 l_2 = -21; end
		2368: begin l_1 = +20;
				 l_2 = +22; end
		2179: begin l_1 = -20;
				 l_2 = -22; end
		3353: begin l_1 = +20;
				 l_2 = +23; end
		3960: begin l_1 = +20;
				 l_2 = -23; end
		587: begin l_1 = -20;
				 l_2 = +23; end
		1194: begin l_1 = -20;
				 l_2 = -23; end
		776: begin l_1 = +20;
				 l_2 = +24; end
		1990: begin l_1 = +20;
				 l_2 = -24; end
		2557: begin l_1 = -20;
				 l_2 = +24; end
		3771: begin l_1 = -20;
				 l_2 = -24; end
		169: begin l_1 = +20;
				 l_2 = +25; end
		2597: begin l_1 = +20;
				 l_2 = -25; end
		1950: begin l_1 = -20;
				 l_2 = +25; end
		4378: begin l_1 = -20;
				 l_2 = -25; end
		3502: begin l_1 = +20;
				 l_2 = +26; end
		3811: begin l_1 = +20;
				 l_2 = -26; end
		736: begin l_1 = -20;
				 l_2 = +26; end
		1045: begin l_1 = -20;
				 l_2 = -26; end
		1074: begin l_1 = +20;
				 l_2 = +27; end
		1692: begin l_1 = +20;
				 l_2 = -27; end
		2855: begin l_1 = -20;
				 l_2 = +27; end
		3473: begin l_1 = -20;
				 l_2 = -27; end
		765: begin l_1 = +20;
				 l_2 = +28; end
		2001: begin l_1 = +20;
				 l_2 = -28; end
		2546: begin l_1 = -20;
				 l_2 = +28; end
		3782: begin l_1 = -20;
				 l_2 = -28; end
		147: begin l_1 = +20;
				 l_2 = +29; end
		2619: begin l_1 = +20;
				 l_2 = -29; end
		1928: begin l_1 = -20;
				 l_2 = +29; end
		4400: begin l_1 = -20;
				 l_2 = -29; end
		3751: begin l_1 = -21;
				 l_2 = +23; end
		796: begin l_1 = -21;
				 l_2 = -22; end
		189: begin l_1 = +21;
				 l_2 = +23; end
		4358: begin l_1 = -21;
				 l_2 = -23; end
		2159: begin l_1 = +21;
				 l_2 = +24; end
		3373: begin l_1 = +21;
				 l_2 = -24; end
		1174: begin l_1 = -21;
				 l_2 = +24; end
		2388: begin l_1 = -21;
				 l_2 = -24; end
		1552: begin l_1 = +21;
				 l_2 = +25; end
		3980: begin l_1 = +21;
				 l_2 = -25; end
		567: begin l_1 = -21;
				 l_2 = +25; end
		2995: begin l_1 = -21;
				 l_2 = -25; end
		338: begin l_1 = +21;
				 l_2 = +26; end
		647: begin l_1 = +21;
				 l_2 = -26; end
		3900: begin l_1 = -21;
				 l_2 = +26; end
		4209: begin l_1 = -21;
				 l_2 = -26; end
		2457: begin l_1 = +21;
				 l_2 = +27; end
		3075: begin l_1 = +21;
				 l_2 = -27; end
		1472: begin l_1 = -21;
				 l_2 = +27; end
		2090: begin l_1 = -21;
				 l_2 = -27; end
		2148: begin l_1 = +21;
				 l_2 = +28; end
		3384: begin l_1 = +21;
				 l_2 = -28; end
		1163: begin l_1 = -21;
				 l_2 = +28; end
		2399: begin l_1 = -21;
				 l_2 = -28; end
		1530: begin l_1 = +21;
				 l_2 = +29; end
		4002: begin l_1 = +21;
				 l_2 = -29; end
		545: begin l_1 = -21;
				 l_2 = +29; end
		3017: begin l_1 = -21;
				 l_2 = -29; end
		2955: begin l_1 = -22;
				 l_2 = +24; end
		1592: begin l_1 = -22;
				 l_2 = -23; end
		378: begin l_1 = +22;
				 l_2 = +24; end
		4169: begin l_1 = -22;
				 l_2 = -24; end
		4318: begin l_1 = +22;
				 l_2 = +25; end
		2199: begin l_1 = +22;
				 l_2 = -25; end
		2348: begin l_1 = -22;
				 l_2 = +25; end
		229: begin l_1 = -22;
				 l_2 = -25; end
		3104: begin l_1 = +22;
				 l_2 = +26; end
		3413: begin l_1 = +22;
				 l_2 = -26; end
		1134: begin l_1 = -22;
				 l_2 = +26; end
		1443: begin l_1 = -22;
				 l_2 = -26; end
		676: begin l_1 = +22;
				 l_2 = +27; end
		1294: begin l_1 = +22;
				 l_2 = -27; end
		3253: begin l_1 = -22;
				 l_2 = +27; end
		3871: begin l_1 = -22;
				 l_2 = -27; end
		367: begin l_1 = +22;
				 l_2 = +28; end
		1603: begin l_1 = +22;
				 l_2 = -28; end
		2944: begin l_1 = -22;
				 l_2 = +28; end
		4180: begin l_1 = -22;
				 l_2 = -28; end
		4296: begin l_1 = +22;
				 l_2 = +29; end
		2221: begin l_1 = +22;
				 l_2 = -29; end
		2326: begin l_1 = -22;
				 l_2 = +29; end
		251: begin l_1 = -22;
				 l_2 = -29; end
		1363: begin l_1 = -23;
				 l_2 = +25; end
		3184: begin l_1 = -23;
				 l_2 = -24; end
		756: begin l_1 = +23;
				 l_2 = +25; end
		3791: begin l_1 = -23;
				 l_2 = -25; end
		4089: begin l_1 = +23;
				 l_2 = +26; end
		4398: begin l_1 = +23;
				 l_2 = -26; end
		149: begin l_1 = -23;
				 l_2 = +26; end
		458: begin l_1 = -23;
				 l_2 = -26; end
		1661: begin l_1 = +23;
				 l_2 = +27; end
		2279: begin l_1 = +23;
				 l_2 = -27; end
		2268: begin l_1 = -23;
				 l_2 = +27; end
		2886: begin l_1 = -23;
				 l_2 = -27; end
		1352: begin l_1 = +23;
				 l_2 = +28; end
		2588: begin l_1 = +23;
				 l_2 = -28; end
		1959: begin l_1 = -23;
				 l_2 = +28; end
		3195: begin l_1 = -23;
				 l_2 = -28; end
		734: begin l_1 = +23;
				 l_2 = +29; end
		3206: begin l_1 = +23;
				 l_2 = -29; end
		1341: begin l_1 = -23;
				 l_2 = +29; end
		3813: begin l_1 = -23;
				 l_2 = -29; end
		2726: begin l_1 = -24;
				 l_2 = +26; end
		1821: begin l_1 = -24;
				 l_2 = -25; end
		1512: begin l_1 = +24;
				 l_2 = +26; end
		3035: begin l_1 = -24;
				 l_2 = -26; end
		3631: begin l_1 = +24;
				 l_2 = +27; end
		4249: begin l_1 = +24;
				 l_2 = -27; end
		298: begin l_1 = -24;
				 l_2 = +27; end
		916: begin l_1 = -24;
				 l_2 = -27; end
		3322: begin l_1 = +24;
				 l_2 = +28; end
		11: begin l_1 = +24;
				 l_2 = -28; end
		4536: begin l_1 = -24;
				 l_2 = +28; end
		1225: begin l_1 = -24;
				 l_2 = -28; end
		2704: begin l_1 = +24;
				 l_2 = +29; end
		629: begin l_1 = +24;
				 l_2 = -29; end
		3918: begin l_1 = -24;
				 l_2 = +29; end
		1843: begin l_1 = -24;
				 l_2 = -29; end
		905: begin l_1 = -25;
				 l_2 = +27; end
		3642: begin l_1 = -25;
				 l_2 = -26; end
		3024: begin l_1 = +25;
				 l_2 = +27; end
		1523: begin l_1 = -25;
				 l_2 = -27; end
		2715: begin l_1 = +25;
				 l_2 = +28; end
		3951: begin l_1 = +25;
				 l_2 = -28; end
		596: begin l_1 = -25;
				 l_2 = +28; end
		1832: begin l_1 = -25;
				 l_2 = -28; end
		2097: begin l_1 = +25;
				 l_2 = +29; end
		22: begin l_1 = +25;
				 l_2 = -29; end
		4525: begin l_1 = -25;
				 l_2 = +29; end
		2450: begin l_1 = -25;
				 l_2 = -29; end
		1810: begin l_1 = -26;
				 l_2 = +28; end
		2737: begin l_1 = -26;
				 l_2 = -27; end
		1501: begin l_1 = +26;
				 l_2 = +28; end
		3046: begin l_1 = -26;
				 l_2 = -28; end
		883: begin l_1 = +26;
				 l_2 = +29; end
		3355: begin l_1 = +26;
				 l_2 = -29; end
		1192: begin l_1 = -26;
				 l_2 = +29; end
		3664: begin l_1 = -26;
				 l_2 = -29; end
		3620: begin l_1 = -27;
				 l_2 = +29; end
		927: begin l_1 = -27;
				 l_2 = -28; end
		3002: begin l_1 = +27;
				 l_2 = +29; end
		1545: begin l_1 = -27;
				 l_2 = -29; end
		2693: begin l_1 = +28;
				 l_2 = +29; end
		1854: begin l_1 = -28;
				 l_2 = -29; end
		default: begin l_1 = 0;
					   l_2 = 0; end
	endcase
end

endmodule

// Product (AN) Code SEC_LUT_Decoder
// SEC_LUT_Decoder16bits.v
// Received codeword W = AN + e, e is single arithmetic weight error (AWE), +2^i or -2^i.
module SEC_LUT_Decoder16bits(W, N);
input 	[28:0]	W;
output	[15:0]	N;
parameter A = 4547;

wire 	[15:0]	Q;
wire 	[12:0]	R;
assign Q = W / A;
assign R = W - (A * Q);

reg	signed	[29:0]	Delta;
always@(*) begin
	case(R)
		1: Delta = 30'sb000000000000000000000000000001;
		4546: Delta = 30'sb111111111111111111111111111111;
		2: Delta = 30'sb000000000000000000000000000010;
		4545: Delta = 30'sb111111111111111111111111111110;
		4: Delta = 30'sb000000000000000000000000000100;
		4543: Delta = 30'sb111111111111111111111111111100;
		8: Delta = 30'sb000000000000000000000000001000;
		4539: Delta = 30'sb111111111111111111111111111000;
		16: Delta = 30'sb000000000000000000000000010000;
		4531: Delta = 30'sb111111111111111111111111110000;
		32: Delta = 30'sb000000000000000000000000100000;
		4515: Delta = 30'sb111111111111111111111111100000;
		64: Delta = 30'sb000000000000000000000001000000;
		4483: Delta = 30'sb111111111111111111111111000000;
		128: Delta = 30'sb000000000000000000000010000000;
		4419: Delta = 30'sb111111111111111111111110000000;
		256: Delta = 30'sb000000000000000000000100000000;
		4291: Delta = 30'sb111111111111111111111100000000;
		512: Delta = 30'sb000000000000000000001000000000;
		4035: Delta = 30'sb111111111111111111111000000000;
		1024: Delta = 30'sb000000000000000000010000000000;
		3523: Delta = 30'sb111111111111111111110000000000;
		2048: Delta = 30'sb000000000000000000100000000000;
		2499: Delta = 30'sb111111111111111111100000000000;
		4096: Delta = 30'sb000000000000000001000000000000;
		451: Delta = 30'sb111111111111111111000000000000;
		3645: Delta = 30'sb000000000000000010000000000000;
		902: Delta = 30'sb111111111111111110000000000000;
		2743: Delta = 30'sb000000000000000100000000000000;
		1804: Delta = 30'sb111111111111111100000000000000;
		939: Delta = 30'sb000000000000001000000000000000;
		3608: Delta = 30'sb111111111111111000000000000000;
		1878: Delta = 30'sb000000000000010000000000000000;
		2669: Delta = 30'sb111111111111110000000000000000;
		3756: Delta = 30'sb000000000000100000000000000000;
		791: Delta = 30'sb111111111111100000000000000000;
		2965: Delta = 30'sb000000000001000000000000000000;
		1582: Delta = 30'sb111111111111000000000000000000;
		1383: Delta = 30'sb000000000010000000000000000000;
		3164: Delta = 30'sb111111111110000000000000000000;
		2766: Delta = 30'sb000000000100000000000000000000;
		1781: Delta = 30'sb111111111100000000000000000000;
		985: Delta = 30'sb000000001000000000000000000000;
		3562: Delta = 30'sb111111111000000000000000000000;
		1970: Delta = 30'sb000000010000000000000000000000;
		2577: Delta = 30'sb111111110000000000000000000000;
		3940: Delta = 30'sb000000100000000000000000000000;
		607: Delta = 30'sb111111100000000000000000000000;
		3333: Delta = 30'sb000001000000000000000000000000;
		1214: Delta = 30'sb111111000000000000000000000000;
		2119: Delta = 30'sb000010000000000000000000000000;
		2428: Delta = 30'sb111110000000000000000000000000;
		4238: Delta = 30'sb000100000000000000000000000000;
		309: Delta = 30'sb111100000000000000000000000000;
		3929: Delta = 30'sb001000000000000000000000000000;
		618: Delta = 30'sb111000000000000000000000000000;
		3311: Delta = 30'sb010000000000000000000000000000;
		1236: Delta = 30'sb110000000000000000000000000000;
		default: Delta =30'sb0;
	endcase
end

assign N = (W - Delta) / A;

endmodule

// Product (AN) Code DEC_LUT_Decoder
// DEC_LUT_Decoder20bits.v
// Received codeword W = AN + E, E is double AWE (E = e1 + e2), +2^i or -2^i.
module DEC_LUT_Decoder20bits_clk(clk, rst_n, W, found, N);

//=========================================================================
//   PARAMETER AND LOCALPARAM FOR FSM
//   W_BITS 要考慮 OVERFLOW 問題
//   N_BITS 也要考慮 OVERFLOW 問題
//=========================================================================
parameter A = 6311 , W_BITS = 34, A_BITS = 13 , N_BITS = 21;

localparam [1:0] idle=2'b00, pre=2'b01,load=2'b10, LUT=2'b11;

reg [1:0] ps;
//==========================================
//   INPUT AND OUTPUT DECLARATION
//==========================================
input   clk, rst_n;
input 	[W_BITS-1:0]	W;
output	reg  [N_BITS-1:0] N;
output  reg  found;

reg 	[N_BITS-1:0]	Q;
reg 	[A_BITS-1:0]	R;

reg	signed	[33:0]	Delta;
always@(*) begin
	case(R)
		1: Delta = 34'sb0000000000000000000000000000000001;
		6310: Delta = 34'sb1111111111111111111111111111111111;
		2: Delta = 34'sb0000000000000000000000000000000010;
		6309: Delta = 34'sb1111111111111111111111111111111110;
		4: Delta = 34'sb0000000000000000000000000000000100;
		6307: Delta = 34'sb1111111111111111111111111111111100;
		8: Delta = 34'sb0000000000000000000000000000001000;
		6303: Delta = 34'sb1111111111111111111111111111111000;
		16: Delta = 34'sb0000000000000000000000000000010000;
		6295: Delta = 34'sb1111111111111111111111111111110000;
		32: Delta = 34'sb0000000000000000000000000000100000;
		6279: Delta = 34'sb1111111111111111111111111111100000;
		64: Delta = 34'sb0000000000000000000000000001000000;
		6247: Delta = 34'sb1111111111111111111111111111000000;
		128: Delta = 34'sb0000000000000000000000000010000000;
		6183: Delta = 34'sb1111111111111111111111111110000000;
		256: Delta = 34'sb0000000000000000000000000100000000;
		6055: Delta = 34'sb1111111111111111111111111100000000;
		512: Delta = 34'sb0000000000000000000000001000000000;
		5799: Delta = 34'sb1111111111111111111111111000000000;
		1024: Delta = 34'sb0000000000000000000000010000000000;
		5287: Delta = 34'sb1111111111111111111111110000000000;
		2048: Delta = 34'sb0000000000000000000000100000000000;
		4263: Delta = 34'sb1111111111111111111111100000000000;
		4096: Delta = 34'sb0000000000000000000001000000000000;
		2215: Delta = 34'sb1111111111111111111111000000000000;
		1881: Delta = 34'sb0000000000000000000010000000000000;
		4430: Delta = 34'sb1111111111111111111110000000000000;
		3762: Delta = 34'sb0000000000000000000100000000000000;
		2549: Delta = 34'sb1111111111111111111100000000000000;
		1213: Delta = 34'sb0000000000000000001000000000000000;
		5098: Delta = 34'sb1111111111111111111000000000000000;
		2426: Delta = 34'sb0000000000000000010000000000000000;
		3885: Delta = 34'sb1111111111111111110000000000000000;
		4852: Delta = 34'sb0000000000000000100000000000000000;
		1459: Delta = 34'sb1111111111111111100000000000000000;
		3393: Delta = 34'sb0000000000000001000000000000000000;
		2918: Delta = 34'sb1111111111111111000000000000000000;
		475: Delta = 34'sb0000000000000010000000000000000000;
		5836: Delta = 34'sb1111111111111110000000000000000000;
		950: Delta = 34'sb0000000000000100000000000000000000;
		5361: Delta = 34'sb1111111111111100000000000000000000;
		1900: Delta = 34'sb0000000000001000000000000000000000;
		4411: Delta = 34'sb1111111111111000000000000000000000;
		3800: Delta = 34'sb0000000000010000000000000000000000;
		2511: Delta = 34'sb1111111111110000000000000000000000;
		1289: Delta = 34'sb0000000000100000000000000000000000;
		5022: Delta = 34'sb1111111111100000000000000000000000;
		2578: Delta = 34'sb0000000001000000000000000000000000;
		3733: Delta = 34'sb1111111111000000000000000000000000;
		5156: Delta = 34'sb0000000010000000000000000000000000;
		1155: Delta = 34'sb1111111110000000000000000000000000;
		4001: Delta = 34'sb0000000100000000000000000000000000;
		2310: Delta = 34'sb1111111100000000000000000000000000;
		1691: Delta = 34'sb0000001000000000000000000000000000;
		4620: Delta = 34'sb1111111000000000000000000000000000;
		3382: Delta = 34'sb0000010000000000000000000000000000;
		2929: Delta = 34'sb1111110000000000000000000000000000;
		453: Delta = 34'sb0000100000000000000000000000000000;
		5858: Delta = 34'sb1111100000000000000000000000000000;
		906: Delta = 34'sb0001000000000000000000000000000000;
		5405: Delta = 34'sb1111000000000000000000000000000000;
		1812: Delta = 34'sb0010000000000000000000000000000000;
		4499: Delta = 34'sb1110000000000000000000000000000000;
		3624: Delta = 34'sb0100000000000000000000000000000000;
		2687: Delta = 34'sb1100000000000000000000000000000000;
		3: Delta = 34'sb0000000000000000000000000000000011;
		6308: Delta = 34'sb1111111111111111111111111111111101;
		5: Delta = 34'sb0000000000000000000000000000000101;
		6306: Delta = 34'sb1111111111111111111111111111111011;
		9: Delta = 34'sb0000000000000000000000000000001001;
		6304: Delta = 34'sb1111111111111111111111111111111001;
		7: Delta = 34'sb0000000000000000000000000000000111;
		6302: Delta = 34'sb1111111111111111111111111111110111;
		17: Delta = 34'sb0000000000000000000000000000010001;
		6296: Delta = 34'sb1111111111111111111111111111110001;
		15: Delta = 34'sb0000000000000000000000000000001111;
		6294: Delta = 34'sb1111111111111111111111111111101111;
		33: Delta = 34'sb0000000000000000000000000000100001;
		6280: Delta = 34'sb1111111111111111111111111111100001;
		31: Delta = 34'sb0000000000000000000000000000011111;
		6278: Delta = 34'sb1111111111111111111111111111011111;
		65: Delta = 34'sb0000000000000000000000000001000001;
		6248: Delta = 34'sb1111111111111111111111111111000001;
		63: Delta = 34'sb0000000000000000000000000000111111;
		6246: Delta = 34'sb1111111111111111111111111110111111;
		129: Delta = 34'sb0000000000000000000000000010000001;
		6184: Delta = 34'sb1111111111111111111111111110000001;
		127: Delta = 34'sb0000000000000000000000000001111111;
		6182: Delta = 34'sb1111111111111111111111111101111111;
		257: Delta = 34'sb0000000000000000000000000100000001;
		6056: Delta = 34'sb1111111111111111111111111100000001;
		255: Delta = 34'sb0000000000000000000000000011111111;
		6054: Delta = 34'sb1111111111111111111111111011111111;
		513: Delta = 34'sb0000000000000000000000001000000001;
		5800: Delta = 34'sb1111111111111111111111111000000001;
		511: Delta = 34'sb0000000000000000000000000111111111;
		5798: Delta = 34'sb1111111111111111111111110111111111;
		1025: Delta = 34'sb0000000000000000000000010000000001;
		5288: Delta = 34'sb1111111111111111111111110000000001;
		1023: Delta = 34'sb0000000000000000000000001111111111;
		5286: Delta = 34'sb1111111111111111111111101111111111;
		2049: Delta = 34'sb0000000000000000000000100000000001;
		4264: Delta = 34'sb1111111111111111111111100000000001;
		2047: Delta = 34'sb0000000000000000000000011111111111;
		4262: Delta = 34'sb1111111111111111111111011111111111;
		4097: Delta = 34'sb0000000000000000000001000000000001;
		2216: Delta = 34'sb1111111111111111111111000000000001;
		4095: Delta = 34'sb0000000000000000000000111111111111;
		2214: Delta = 34'sb1111111111111111111110111111111111;
		1882: Delta = 34'sb0000000000000000000010000000000001;
		4431: Delta = 34'sb1111111111111111111110000000000001;
		1880: Delta = 34'sb0000000000000000000001111111111111;
		4429: Delta = 34'sb1111111111111111111101111111111111;
		3763: Delta = 34'sb0000000000000000000100000000000001;
		2550: Delta = 34'sb1111111111111111111100000000000001;
		3761: Delta = 34'sb0000000000000000000011111111111111;
		2548: Delta = 34'sb1111111111111111111011111111111111;
		1214: Delta = 34'sb0000000000000000001000000000000001;
		5099: Delta = 34'sb1111111111111111111000000000000001;
		1212: Delta = 34'sb0000000000000000000111111111111111;
		5097: Delta = 34'sb1111111111111111110111111111111111;
		2427: Delta = 34'sb0000000000000000010000000000000001;
		3886: Delta = 34'sb1111111111111111110000000000000001;
		2425: Delta = 34'sb0000000000000000001111111111111111;
		3884: Delta = 34'sb1111111111111111101111111111111111;
		4853: Delta = 34'sb0000000000000000100000000000000001;
		1460: Delta = 34'sb1111111111111111100000000000000001;
		4851: Delta = 34'sb0000000000000000011111111111111111;
		1458: Delta = 34'sb1111111111111111011111111111111111;
		3394: Delta = 34'sb0000000000000001000000000000000001;
		2919: Delta = 34'sb1111111111111111000000000000000001;
		3392: Delta = 34'sb0000000000000000111111111111111111;
		2917: Delta = 34'sb1111111111111110111111111111111111;
		476: Delta = 34'sb0000000000000010000000000000000001;
		5837: Delta = 34'sb1111111111111110000000000000000001;
		474: Delta = 34'sb0000000000000001111111111111111111;
		5835: Delta = 34'sb1111111111111101111111111111111111;
		951: Delta = 34'sb0000000000000100000000000000000001;
		5362: Delta = 34'sb1111111111111100000000000000000001;
		949: Delta = 34'sb0000000000000011111111111111111111;
		5360: Delta = 34'sb1111111111111011111111111111111111;
		1901: Delta = 34'sb0000000000001000000000000000000001;
		4412: Delta = 34'sb1111111111111000000000000000000001;
		1899: Delta = 34'sb0000000000000111111111111111111111;
		4410: Delta = 34'sb1111111111110111111111111111111111;
		3801: Delta = 34'sb0000000000010000000000000000000001;
		2512: Delta = 34'sb1111111111110000000000000000000001;
		3799: Delta = 34'sb0000000000001111111111111111111111;
		2510: Delta = 34'sb1111111111101111111111111111111111;
		1290: Delta = 34'sb0000000000100000000000000000000001;
		5023: Delta = 34'sb1111111111100000000000000000000001;
		1288: Delta = 34'sb0000000000011111111111111111111111;
		5021: Delta = 34'sb1111111111011111111111111111111111;
		2579: Delta = 34'sb0000000001000000000000000000000001;
		3734: Delta = 34'sb1111111111000000000000000000000001;
		2577: Delta = 34'sb0000000000111111111111111111111111;
		3732: Delta = 34'sb1111111110111111111111111111111111;
		5157: Delta = 34'sb0000000010000000000000000000000001;
		1156: Delta = 34'sb1111111110000000000000000000000001;
		5155: Delta = 34'sb0000000001111111111111111111111111;
		1154: Delta = 34'sb1111111101111111111111111111111111;
		4002: Delta = 34'sb0000000100000000000000000000000001;
		2311: Delta = 34'sb1111111100000000000000000000000001;
		4000: Delta = 34'sb0000000011111111111111111111111111;
		2309: Delta = 34'sb1111111011111111111111111111111111;
		1692: Delta = 34'sb0000001000000000000000000000000001;
		4621: Delta = 34'sb1111111000000000000000000000000001;
		1690: Delta = 34'sb0000000111111111111111111111111111;
		4619: Delta = 34'sb1111110111111111111111111111111111;
		3383: Delta = 34'sb0000010000000000000000000000000001;
		2930: Delta = 34'sb1111110000000000000000000000000001;
		3381: Delta = 34'sb0000001111111111111111111111111111;
		2928: Delta = 34'sb1111101111111111111111111111111111;
		454: Delta = 34'sb0000100000000000000000000000000001;
		5859: Delta = 34'sb1111100000000000000000000000000001;
		452: Delta = 34'sb0000011111111111111111111111111111;
		5857: Delta = 34'sb1111011111111111111111111111111111;
		907: Delta = 34'sb0001000000000000000000000000000001;
		5406: Delta = 34'sb1111000000000000000000000000000001;
		905: Delta = 34'sb0000111111111111111111111111111111;
		5404: Delta = 34'sb1110111111111111111111111111111111;
		1813: Delta = 34'sb0010000000000000000000000000000001;
		4500: Delta = 34'sb1110000000000000000000000000000001;
		1811: Delta = 34'sb0001111111111111111111111111111111;
		4498: Delta = 34'sb1101111111111111111111111111111111;
		3625: Delta = 34'sb0100000000000000000000000000000001;
		2688: Delta = 34'sb1100000000000000000000000000000001;
		3623: Delta = 34'sb0011111111111111111111111111111111;
		2686: Delta = 34'sb1011111111111111111111111111111111;
		6: Delta = 34'sb0000000000000000000000000000000110;
		6305: Delta = 34'sb1111111111111111111111111111111010;
		10: Delta = 34'sb0000000000000000000000000000001010;
		6301: Delta = 34'sb1111111111111111111111111111110110;
		18: Delta = 34'sb0000000000000000000000000000010010;
		6297: Delta = 34'sb1111111111111111111111111111110010;
		14: Delta = 34'sb0000000000000000000000000000001110;
		6293: Delta = 34'sb1111111111111111111111111111101110;
		34: Delta = 34'sb0000000000000000000000000000100010;
		6281: Delta = 34'sb1111111111111111111111111111100010;
		30: Delta = 34'sb0000000000000000000000000000011110;
		6277: Delta = 34'sb1111111111111111111111111111011110;
		66: Delta = 34'sb0000000000000000000000000001000010;
		6249: Delta = 34'sb1111111111111111111111111111000010;
		62: Delta = 34'sb0000000000000000000000000000111110;
		6245: Delta = 34'sb1111111111111111111111111110111110;
		130: Delta = 34'sb0000000000000000000000000010000010;
		6185: Delta = 34'sb1111111111111111111111111110000010;
		126: Delta = 34'sb0000000000000000000000000001111110;
		6181: Delta = 34'sb1111111111111111111111111101111110;
		258: Delta = 34'sb0000000000000000000000000100000010;
		6057: Delta = 34'sb1111111111111111111111111100000010;
		254: Delta = 34'sb0000000000000000000000000011111110;
		6053: Delta = 34'sb1111111111111111111111111011111110;
		514: Delta = 34'sb0000000000000000000000001000000010;
		5801: Delta = 34'sb1111111111111111111111111000000010;
		510: Delta = 34'sb0000000000000000000000000111111110;
		5797: Delta = 34'sb1111111111111111111111110111111110;
		1026: Delta = 34'sb0000000000000000000000010000000010;
		5289: Delta = 34'sb1111111111111111111111110000000010;
		1022: Delta = 34'sb0000000000000000000000001111111110;
		5285: Delta = 34'sb1111111111111111111111101111111110;
		2050: Delta = 34'sb0000000000000000000000100000000010;
		4265: Delta = 34'sb1111111111111111111111100000000010;
		2046: Delta = 34'sb0000000000000000000000011111111110;
		4261: Delta = 34'sb1111111111111111111111011111111110;
		4098: Delta = 34'sb0000000000000000000001000000000010;
		2217: Delta = 34'sb1111111111111111111111000000000010;
		4094: Delta = 34'sb0000000000000000000000111111111110;
		2213: Delta = 34'sb1111111111111111111110111111111110;
		1883: Delta = 34'sb0000000000000000000010000000000010;
		4432: Delta = 34'sb1111111111111111111110000000000010;
		1879: Delta = 34'sb0000000000000000000001111111111110;
		4428: Delta = 34'sb1111111111111111111101111111111110;
		3764: Delta = 34'sb0000000000000000000100000000000010;
		2551: Delta = 34'sb1111111111111111111100000000000010;
		3760: Delta = 34'sb0000000000000000000011111111111110;
		2547: Delta = 34'sb1111111111111111111011111111111110;
		1215: Delta = 34'sb0000000000000000001000000000000010;
		5100: Delta = 34'sb1111111111111111111000000000000010;
		1211: Delta = 34'sb0000000000000000000111111111111110;
		5096: Delta = 34'sb1111111111111111110111111111111110;
		2428: Delta = 34'sb0000000000000000010000000000000010;
		3887: Delta = 34'sb1111111111111111110000000000000010;
		2424: Delta = 34'sb0000000000000000001111111111111110;
		3883: Delta = 34'sb1111111111111111101111111111111110;
		4854: Delta = 34'sb0000000000000000100000000000000010;
		1461: Delta = 34'sb1111111111111111100000000000000010;
		4850: Delta = 34'sb0000000000000000011111111111111110;
		1457: Delta = 34'sb1111111111111111011111111111111110;
		3395: Delta = 34'sb0000000000000001000000000000000010;
		2920: Delta = 34'sb1111111111111111000000000000000010;
		3391: Delta = 34'sb0000000000000000111111111111111110;
		2916: Delta = 34'sb1111111111111110111111111111111110;
		477: Delta = 34'sb0000000000000010000000000000000010;
		5838: Delta = 34'sb1111111111111110000000000000000010;
		473: Delta = 34'sb0000000000000001111111111111111110;
		5834: Delta = 34'sb1111111111111101111111111111111110;
		952: Delta = 34'sb0000000000000100000000000000000010;
		5363: Delta = 34'sb1111111111111100000000000000000010;
		948: Delta = 34'sb0000000000000011111111111111111110;
		5359: Delta = 34'sb1111111111111011111111111111111110;
		1902: Delta = 34'sb0000000000001000000000000000000010;
		4413: Delta = 34'sb1111111111111000000000000000000010;
		1898: Delta = 34'sb0000000000000111111111111111111110;
		4409: Delta = 34'sb1111111111110111111111111111111110;
		3802: Delta = 34'sb0000000000010000000000000000000010;
		2513: Delta = 34'sb1111111111110000000000000000000010;
		3798: Delta = 34'sb0000000000001111111111111111111110;
		2509: Delta = 34'sb1111111111101111111111111111111110;
		1291: Delta = 34'sb0000000000100000000000000000000010;
		5024: Delta = 34'sb1111111111100000000000000000000010;
		1287: Delta = 34'sb0000000000011111111111111111111110;
		5020: Delta = 34'sb1111111111011111111111111111111110;
		2580: Delta = 34'sb0000000001000000000000000000000010;
		3735: Delta = 34'sb1111111111000000000000000000000010;
		2576: Delta = 34'sb0000000000111111111111111111111110;
		3731: Delta = 34'sb1111111110111111111111111111111110;
		5158: Delta = 34'sb0000000010000000000000000000000010;
		1157: Delta = 34'sb1111111110000000000000000000000010;
		5154: Delta = 34'sb0000000001111111111111111111111110;
		1153: Delta = 34'sb1111111101111111111111111111111110;
		4003: Delta = 34'sb0000000100000000000000000000000010;
		2312: Delta = 34'sb1111111100000000000000000000000010;
		3999: Delta = 34'sb0000000011111111111111111111111110;
		2308: Delta = 34'sb1111111011111111111111111111111110;
		1693: Delta = 34'sb0000001000000000000000000000000010;
		4622: Delta = 34'sb1111111000000000000000000000000010;
		1689: Delta = 34'sb0000000111111111111111111111111110;
		4618: Delta = 34'sb1111110111111111111111111111111110;
		3384: Delta = 34'sb0000010000000000000000000000000010;
		2931: Delta = 34'sb1111110000000000000000000000000010;
		3380: Delta = 34'sb0000001111111111111111111111111110;
		2927: Delta = 34'sb1111101111111111111111111111111110;
		455: Delta = 34'sb0000100000000000000000000000000010;
		5860: Delta = 34'sb1111100000000000000000000000000010;
		451: Delta = 34'sb0000011111111111111111111111111110;
		5856: Delta = 34'sb1111011111111111111111111111111110;
		908: Delta = 34'sb0001000000000000000000000000000010;
		5407: Delta = 34'sb1111000000000000000000000000000010;
		904: Delta = 34'sb0000111111111111111111111111111110;
		5403: Delta = 34'sb1110111111111111111111111111111110;
		1814: Delta = 34'sb0010000000000000000000000000000010;
		4501: Delta = 34'sb1110000000000000000000000000000010;
		1810: Delta = 34'sb0001111111111111111111111111111110;
		4497: Delta = 34'sb1101111111111111111111111111111110;
		3626: Delta = 34'sb0100000000000000000000000000000010;
		2689: Delta = 34'sb1100000000000000000000000000000010;
		3622: Delta = 34'sb0011111111111111111111111111111110;
		2685: Delta = 34'sb1011111111111111111111111111111110;
		12: Delta = 34'sb0000000000000000000000000000001100;
		6299: Delta = 34'sb1111111111111111111111111111110100;
		20: Delta = 34'sb0000000000000000000000000000010100;
		6291: Delta = 34'sb1111111111111111111111111111101100;
		36: Delta = 34'sb0000000000000000000000000000100100;
		6283: Delta = 34'sb1111111111111111111111111111100100;
		28: Delta = 34'sb0000000000000000000000000000011100;
		6275: Delta = 34'sb1111111111111111111111111111011100;
		68: Delta = 34'sb0000000000000000000000000001000100;
		6251: Delta = 34'sb1111111111111111111111111111000100;
		60: Delta = 34'sb0000000000000000000000000000111100;
		6243: Delta = 34'sb1111111111111111111111111110111100;
		132: Delta = 34'sb0000000000000000000000000010000100;
		6187: Delta = 34'sb1111111111111111111111111110000100;
		124: Delta = 34'sb0000000000000000000000000001111100;
		6179: Delta = 34'sb1111111111111111111111111101111100;
		260: Delta = 34'sb0000000000000000000000000100000100;
		6059: Delta = 34'sb1111111111111111111111111100000100;
		252: Delta = 34'sb0000000000000000000000000011111100;
		6051: Delta = 34'sb1111111111111111111111111011111100;
		516: Delta = 34'sb0000000000000000000000001000000100;
		5803: Delta = 34'sb1111111111111111111111111000000100;
		508: Delta = 34'sb0000000000000000000000000111111100;
		5795: Delta = 34'sb1111111111111111111111110111111100;
		1028: Delta = 34'sb0000000000000000000000010000000100;
		5291: Delta = 34'sb1111111111111111111111110000000100;
		1020: Delta = 34'sb0000000000000000000000001111111100;
		5283: Delta = 34'sb1111111111111111111111101111111100;
		2052: Delta = 34'sb0000000000000000000000100000000100;
		4267: Delta = 34'sb1111111111111111111111100000000100;
		2044: Delta = 34'sb0000000000000000000000011111111100;
		4259: Delta = 34'sb1111111111111111111111011111111100;
		4100: Delta = 34'sb0000000000000000000001000000000100;
		2219: Delta = 34'sb1111111111111111111111000000000100;
		4092: Delta = 34'sb0000000000000000000000111111111100;
		2211: Delta = 34'sb1111111111111111111110111111111100;
		1885: Delta = 34'sb0000000000000000000010000000000100;
		4434: Delta = 34'sb1111111111111111111110000000000100;
		1877: Delta = 34'sb0000000000000000000001111111111100;
		4426: Delta = 34'sb1111111111111111111101111111111100;
		3766: Delta = 34'sb0000000000000000000100000000000100;
		2553: Delta = 34'sb1111111111111111111100000000000100;
		3758: Delta = 34'sb0000000000000000000011111111111100;
		2545: Delta = 34'sb1111111111111111111011111111111100;
		1217: Delta = 34'sb0000000000000000001000000000000100;
		5102: Delta = 34'sb1111111111111111111000000000000100;
		1209: Delta = 34'sb0000000000000000000111111111111100;
		5094: Delta = 34'sb1111111111111111110111111111111100;
		2430: Delta = 34'sb0000000000000000010000000000000100;
		3889: Delta = 34'sb1111111111111111110000000000000100;
		2422: Delta = 34'sb0000000000000000001111111111111100;
		3881: Delta = 34'sb1111111111111111101111111111111100;
		4856: Delta = 34'sb0000000000000000100000000000000100;
		1463: Delta = 34'sb1111111111111111100000000000000100;
		4848: Delta = 34'sb0000000000000000011111111111111100;
		1455: Delta = 34'sb1111111111111111011111111111111100;
		3397: Delta = 34'sb0000000000000001000000000000000100;
		2922: Delta = 34'sb1111111111111111000000000000000100;
		3389: Delta = 34'sb0000000000000000111111111111111100;
		2914: Delta = 34'sb1111111111111110111111111111111100;
		479: Delta = 34'sb0000000000000010000000000000000100;
		5840: Delta = 34'sb1111111111111110000000000000000100;
		471: Delta = 34'sb0000000000000001111111111111111100;
		5832: Delta = 34'sb1111111111111101111111111111111100;
		954: Delta = 34'sb0000000000000100000000000000000100;
		5365: Delta = 34'sb1111111111111100000000000000000100;
		946: Delta = 34'sb0000000000000011111111111111111100;
		5357: Delta = 34'sb1111111111111011111111111111111100;
		1904: Delta = 34'sb0000000000001000000000000000000100;
		4415: Delta = 34'sb1111111111111000000000000000000100;
		1896: Delta = 34'sb0000000000000111111111111111111100;
		4407: Delta = 34'sb1111111111110111111111111111111100;
		3804: Delta = 34'sb0000000000010000000000000000000100;
		2515: Delta = 34'sb1111111111110000000000000000000100;
		3796: Delta = 34'sb0000000000001111111111111111111100;
		2507: Delta = 34'sb1111111111101111111111111111111100;
		1293: Delta = 34'sb0000000000100000000000000000000100;
		5026: Delta = 34'sb1111111111100000000000000000000100;
		1285: Delta = 34'sb0000000000011111111111111111111100;
		5018: Delta = 34'sb1111111111011111111111111111111100;
		2582: Delta = 34'sb0000000001000000000000000000000100;
		3737: Delta = 34'sb1111111111000000000000000000000100;
		2574: Delta = 34'sb0000000000111111111111111111111100;
		3729: Delta = 34'sb1111111110111111111111111111111100;
		5160: Delta = 34'sb0000000010000000000000000000000100;
		1159: Delta = 34'sb1111111110000000000000000000000100;
		5152: Delta = 34'sb0000000001111111111111111111111100;
		1151: Delta = 34'sb1111111101111111111111111111111100;
		4005: Delta = 34'sb0000000100000000000000000000000100;
		2314: Delta = 34'sb1111111100000000000000000000000100;
		3997: Delta = 34'sb0000000011111111111111111111111100;
		2306: Delta = 34'sb1111111011111111111111111111111100;
		1695: Delta = 34'sb0000001000000000000000000000000100;
		4624: Delta = 34'sb1111111000000000000000000000000100;
		1687: Delta = 34'sb0000000111111111111111111111111100;
		4616: Delta = 34'sb1111110111111111111111111111111100;
		3386: Delta = 34'sb0000010000000000000000000000000100;
		2933: Delta = 34'sb1111110000000000000000000000000100;
		3378: Delta = 34'sb0000001111111111111111111111111100;
		2925: Delta = 34'sb1111101111111111111111111111111100;
		457: Delta = 34'sb0000100000000000000000000000000100;
		5862: Delta = 34'sb1111100000000000000000000000000100;
		449: Delta = 34'sb0000011111111111111111111111111100;
		5854: Delta = 34'sb1111011111111111111111111111111100;
		910: Delta = 34'sb0001000000000000000000000000000100;
		5409: Delta = 34'sb1111000000000000000000000000000100;
		902: Delta = 34'sb0000111111111111111111111111111100;
		5401: Delta = 34'sb1110111111111111111111111111111100;
		1816: Delta = 34'sb0010000000000000000000000000000100;
		4503: Delta = 34'sb1110000000000000000000000000000100;
		1808: Delta = 34'sb0001111111111111111111111111111100;
		4495: Delta = 34'sb1101111111111111111111111111111100;
		3628: Delta = 34'sb0100000000000000000000000000000100;
		2691: Delta = 34'sb1100000000000000000000000000000100;
		3620: Delta = 34'sb0011111111111111111111111111111100;
		2683: Delta = 34'sb1011111111111111111111111111111100;
		24: Delta = 34'sb0000000000000000000000000000011000;
		6287: Delta = 34'sb1111111111111111111111111111101000;
		40: Delta = 34'sb0000000000000000000000000000101000;
		6271: Delta = 34'sb1111111111111111111111111111011000;
		72: Delta = 34'sb0000000000000000000000000001001000;
		6255: Delta = 34'sb1111111111111111111111111111001000;
		56: Delta = 34'sb0000000000000000000000000000111000;
		6239: Delta = 34'sb1111111111111111111111111110111000;
		136: Delta = 34'sb0000000000000000000000000010001000;
		6191: Delta = 34'sb1111111111111111111111111110001000;
		120: Delta = 34'sb0000000000000000000000000001111000;
		6175: Delta = 34'sb1111111111111111111111111101111000;
		264: Delta = 34'sb0000000000000000000000000100001000;
		6063: Delta = 34'sb1111111111111111111111111100001000;
		248: Delta = 34'sb0000000000000000000000000011111000;
		6047: Delta = 34'sb1111111111111111111111111011111000;
		520: Delta = 34'sb0000000000000000000000001000001000;
		5807: Delta = 34'sb1111111111111111111111111000001000;
		504: Delta = 34'sb0000000000000000000000000111111000;
		5791: Delta = 34'sb1111111111111111111111110111111000;
		1032: Delta = 34'sb0000000000000000000000010000001000;
		5295: Delta = 34'sb1111111111111111111111110000001000;
		1016: Delta = 34'sb0000000000000000000000001111111000;
		5279: Delta = 34'sb1111111111111111111111101111111000;
		2056: Delta = 34'sb0000000000000000000000100000001000;
		4271: Delta = 34'sb1111111111111111111111100000001000;
		2040: Delta = 34'sb0000000000000000000000011111111000;
		4255: Delta = 34'sb1111111111111111111111011111111000;
		4104: Delta = 34'sb0000000000000000000001000000001000;
		2223: Delta = 34'sb1111111111111111111111000000001000;
		4088: Delta = 34'sb0000000000000000000000111111111000;
		2207: Delta = 34'sb1111111111111111111110111111111000;
		1889: Delta = 34'sb0000000000000000000010000000001000;
		4438: Delta = 34'sb1111111111111111111110000000001000;
		1873: Delta = 34'sb0000000000000000000001111111111000;
		4422: Delta = 34'sb1111111111111111111101111111111000;
		3770: Delta = 34'sb0000000000000000000100000000001000;
		2557: Delta = 34'sb1111111111111111111100000000001000;
		3754: Delta = 34'sb0000000000000000000011111111111000;
		2541: Delta = 34'sb1111111111111111111011111111111000;
		1221: Delta = 34'sb0000000000000000001000000000001000;
		5106: Delta = 34'sb1111111111111111111000000000001000;
		1205: Delta = 34'sb0000000000000000000111111111111000;
		5090: Delta = 34'sb1111111111111111110111111111111000;
		2434: Delta = 34'sb0000000000000000010000000000001000;
		3893: Delta = 34'sb1111111111111111110000000000001000;
		2418: Delta = 34'sb0000000000000000001111111111111000;
		3877: Delta = 34'sb1111111111111111101111111111111000;
		4860: Delta = 34'sb0000000000000000100000000000001000;
		1467: Delta = 34'sb1111111111111111100000000000001000;
		4844: Delta = 34'sb0000000000000000011111111111111000;
		1451: Delta = 34'sb1111111111111111011111111111111000;
		3401: Delta = 34'sb0000000000000001000000000000001000;
		2926: Delta = 34'sb1111111111111111000000000000001000;
		3385: Delta = 34'sb0000000000000000111111111111111000;
		2910: Delta = 34'sb1111111111111110111111111111111000;
		483: Delta = 34'sb0000000000000010000000000000001000;
		5844: Delta = 34'sb1111111111111110000000000000001000;
		467: Delta = 34'sb0000000000000001111111111111111000;
		5828: Delta = 34'sb1111111111111101111111111111111000;
		958: Delta = 34'sb0000000000000100000000000000001000;
		5369: Delta = 34'sb1111111111111100000000000000001000;
		942: Delta = 34'sb0000000000000011111111111111111000;
		5353: Delta = 34'sb1111111111111011111111111111111000;
		1908: Delta = 34'sb0000000000001000000000000000001000;
		4419: Delta = 34'sb1111111111111000000000000000001000;
		1892: Delta = 34'sb0000000000000111111111111111111000;
		4403: Delta = 34'sb1111111111110111111111111111111000;
		3808: Delta = 34'sb0000000000010000000000000000001000;
		2519: Delta = 34'sb1111111111110000000000000000001000;
		3792: Delta = 34'sb0000000000001111111111111111111000;
		2503: Delta = 34'sb1111111111101111111111111111111000;
		1297: Delta = 34'sb0000000000100000000000000000001000;
		5030: Delta = 34'sb1111111111100000000000000000001000;
		1281: Delta = 34'sb0000000000011111111111111111111000;
		5014: Delta = 34'sb1111111111011111111111111111111000;
		2586: Delta = 34'sb0000000001000000000000000000001000;
		3741: Delta = 34'sb1111111111000000000000000000001000;
		2570: Delta = 34'sb0000000000111111111111111111111000;
		3725: Delta = 34'sb1111111110111111111111111111111000;
		5164: Delta = 34'sb0000000010000000000000000000001000;
		1163: Delta = 34'sb1111111110000000000000000000001000;
		5148: Delta = 34'sb0000000001111111111111111111111000;
		1147: Delta = 34'sb1111111101111111111111111111111000;
		4009: Delta = 34'sb0000000100000000000000000000001000;
		2318: Delta = 34'sb1111111100000000000000000000001000;
		3993: Delta = 34'sb0000000011111111111111111111111000;
		2302: Delta = 34'sb1111111011111111111111111111111000;
		1699: Delta = 34'sb0000001000000000000000000000001000;
		4628: Delta = 34'sb1111111000000000000000000000001000;
		1683: Delta = 34'sb0000000111111111111111111111111000;
		4612: Delta = 34'sb1111110111111111111111111111111000;
		3390: Delta = 34'sb0000010000000000000000000000001000;
		2937: Delta = 34'sb1111110000000000000000000000001000;
		3374: Delta = 34'sb0000001111111111111111111111111000;
		2921: Delta = 34'sb1111101111111111111111111111111000;
		461: Delta = 34'sb0000100000000000000000000000001000;
		5866: Delta = 34'sb1111100000000000000000000000001000;
		445: Delta = 34'sb0000011111111111111111111111111000;
		5850: Delta = 34'sb1111011111111111111111111111111000;
		914: Delta = 34'sb0001000000000000000000000000001000;
		5413: Delta = 34'sb1111000000000000000000000000001000;
		898: Delta = 34'sb0000111111111111111111111111111000;
		5397: Delta = 34'sb1110111111111111111111111111111000;
		1820: Delta = 34'sb0010000000000000000000000000001000;
		4507: Delta = 34'sb1110000000000000000000000000001000;
		1804: Delta = 34'sb0001111111111111111111111111111000;
		4491: Delta = 34'sb1101111111111111111111111111111000;
		3632: Delta = 34'sb0100000000000000000000000000001000;
		2695: Delta = 34'sb1100000000000000000000000000001000;
		3616: Delta = 34'sb0011111111111111111111111111111000;
		2679: Delta = 34'sb1011111111111111111111111111111000;
		48: Delta = 34'sb0000000000000000000000000000110000;
		6263: Delta = 34'sb1111111111111111111111111111010000;
		80: Delta = 34'sb0000000000000000000000000001010000;
		6231: Delta = 34'sb1111111111111111111111111110110000;
		144: Delta = 34'sb0000000000000000000000000010010000;
		6199: Delta = 34'sb1111111111111111111111111110010000;
		112: Delta = 34'sb0000000000000000000000000001110000;
		6167: Delta = 34'sb1111111111111111111111111101110000;
		272: Delta = 34'sb0000000000000000000000000100010000;
		6071: Delta = 34'sb1111111111111111111111111100010000;
		240: Delta = 34'sb0000000000000000000000000011110000;
		6039: Delta = 34'sb1111111111111111111111111011110000;
		528: Delta = 34'sb0000000000000000000000001000010000;
		5815: Delta = 34'sb1111111111111111111111111000010000;
		496: Delta = 34'sb0000000000000000000000000111110000;
		5783: Delta = 34'sb1111111111111111111111110111110000;
		1040: Delta = 34'sb0000000000000000000000010000010000;
		5303: Delta = 34'sb1111111111111111111111110000010000;
		1008: Delta = 34'sb0000000000000000000000001111110000;
		5271: Delta = 34'sb1111111111111111111111101111110000;
		2064: Delta = 34'sb0000000000000000000000100000010000;
		4279: Delta = 34'sb1111111111111111111111100000010000;
		2032: Delta = 34'sb0000000000000000000000011111110000;
		4247: Delta = 34'sb1111111111111111111111011111110000;
		4112: Delta = 34'sb0000000000000000000001000000010000;
		2231: Delta = 34'sb1111111111111111111111000000010000;
		4080: Delta = 34'sb0000000000000000000000111111110000;
		2199: Delta = 34'sb1111111111111111111110111111110000;
		1897: Delta = 34'sb0000000000000000000010000000010000;
		4446: Delta = 34'sb1111111111111111111110000000010000;
		1865: Delta = 34'sb0000000000000000000001111111110000;
		4414: Delta = 34'sb1111111111111111111101111111110000;
		3778: Delta = 34'sb0000000000000000000100000000010000;
		2565: Delta = 34'sb1111111111111111111100000000010000;
		3746: Delta = 34'sb0000000000000000000011111111110000;
		2533: Delta = 34'sb1111111111111111111011111111110000;
		1229: Delta = 34'sb0000000000000000001000000000010000;
		5114: Delta = 34'sb1111111111111111111000000000010000;
		1197: Delta = 34'sb0000000000000000000111111111110000;
		5082: Delta = 34'sb1111111111111111110111111111110000;
		2442: Delta = 34'sb0000000000000000010000000000010000;
		3901: Delta = 34'sb1111111111111111110000000000010000;
		2410: Delta = 34'sb0000000000000000001111111111110000;
		3869: Delta = 34'sb1111111111111111101111111111110000;
		4868: Delta = 34'sb0000000000000000100000000000010000;
		1475: Delta = 34'sb1111111111111111100000000000010000;
		4836: Delta = 34'sb0000000000000000011111111111110000;
		1443: Delta = 34'sb1111111111111111011111111111110000;
		3409: Delta = 34'sb0000000000000001000000000000010000;
		2934: Delta = 34'sb1111111111111111000000000000010000;
		3377: Delta = 34'sb0000000000000000111111111111110000;
		2902: Delta = 34'sb1111111111111110111111111111110000;
		491: Delta = 34'sb0000000000000010000000000000010000;
		5852: Delta = 34'sb1111111111111110000000000000010000;
		459: Delta = 34'sb0000000000000001111111111111110000;
		5820: Delta = 34'sb1111111111111101111111111111110000;
		966: Delta = 34'sb0000000000000100000000000000010000;
		5377: Delta = 34'sb1111111111111100000000000000010000;
		934: Delta = 34'sb0000000000000011111111111111110000;
		5345: Delta = 34'sb1111111111111011111111111111110000;
		1916: Delta = 34'sb0000000000001000000000000000010000;
		4427: Delta = 34'sb1111111111111000000000000000010000;
		1884: Delta = 34'sb0000000000000111111111111111110000;
		4395: Delta = 34'sb1111111111110111111111111111110000;
		3816: Delta = 34'sb0000000000010000000000000000010000;
		2527: Delta = 34'sb1111111111110000000000000000010000;
		3784: Delta = 34'sb0000000000001111111111111111110000;
		2495: Delta = 34'sb1111111111101111111111111111110000;
		1305: Delta = 34'sb0000000000100000000000000000010000;
		5038: Delta = 34'sb1111111111100000000000000000010000;
		1273: Delta = 34'sb0000000000011111111111111111110000;
		5006: Delta = 34'sb1111111111011111111111111111110000;
		2594: Delta = 34'sb0000000001000000000000000000010000;
		3749: Delta = 34'sb1111111111000000000000000000010000;
		2562: Delta = 34'sb0000000000111111111111111111110000;
		3717: Delta = 34'sb1111111110111111111111111111110000;
		5172: Delta = 34'sb0000000010000000000000000000010000;
		1171: Delta = 34'sb1111111110000000000000000000010000;
		5140: Delta = 34'sb0000000001111111111111111111110000;
		1139: Delta = 34'sb1111111101111111111111111111110000;
		4017: Delta = 34'sb0000000100000000000000000000010000;
		2326: Delta = 34'sb1111111100000000000000000000010000;
		3985: Delta = 34'sb0000000011111111111111111111110000;
		2294: Delta = 34'sb1111111011111111111111111111110000;
		1707: Delta = 34'sb0000001000000000000000000000010000;
		4636: Delta = 34'sb1111111000000000000000000000010000;
		1675: Delta = 34'sb0000000111111111111111111111110000;
		4604: Delta = 34'sb1111110111111111111111111111110000;
		3398: Delta = 34'sb0000010000000000000000000000010000;
		2945: Delta = 34'sb1111110000000000000000000000010000;
		3366: Delta = 34'sb0000001111111111111111111111110000;
		2913: Delta = 34'sb1111101111111111111111111111110000;
		469: Delta = 34'sb0000100000000000000000000000010000;
		5874: Delta = 34'sb1111100000000000000000000000010000;
		437: Delta = 34'sb0000011111111111111111111111110000;
		5842: Delta = 34'sb1111011111111111111111111111110000;
		922: Delta = 34'sb0001000000000000000000000000010000;
		5421: Delta = 34'sb1111000000000000000000000000010000;
		890: Delta = 34'sb0000111111111111111111111111110000;
		5389: Delta = 34'sb1110111111111111111111111111110000;
		1828: Delta = 34'sb0010000000000000000000000000010000;
		4515: Delta = 34'sb1110000000000000000000000000010000;
		1796: Delta = 34'sb0001111111111111111111111111110000;
		4483: Delta = 34'sb1101111111111111111111111111110000;
		3640: Delta = 34'sb0100000000000000000000000000010000;
		2703: Delta = 34'sb1100000000000000000000000000010000;
		3608: Delta = 34'sb0011111111111111111111111111110000;
		2671: Delta = 34'sb1011111111111111111111111111110000;
		96: Delta = 34'sb0000000000000000000000000001100000;
		6215: Delta = 34'sb1111111111111111111111111110100000;
		160: Delta = 34'sb0000000000000000000000000010100000;
		6151: Delta = 34'sb1111111111111111111111111101100000;
		288: Delta = 34'sb0000000000000000000000000100100000;
		6087: Delta = 34'sb1111111111111111111111111100100000;
		224: Delta = 34'sb0000000000000000000000000011100000;
		6023: Delta = 34'sb1111111111111111111111111011100000;
		544: Delta = 34'sb0000000000000000000000001000100000;
		5831: Delta = 34'sb1111111111111111111111111000100000;
		480: Delta = 34'sb0000000000000000000000000111100000;
		5767: Delta = 34'sb1111111111111111111111110111100000;
		1056: Delta = 34'sb0000000000000000000000010000100000;
		5319: Delta = 34'sb1111111111111111111111110000100000;
		992: Delta = 34'sb0000000000000000000000001111100000;
		5255: Delta = 34'sb1111111111111111111111101111100000;
		2080: Delta = 34'sb0000000000000000000000100000100000;
		4295: Delta = 34'sb1111111111111111111111100000100000;
		2016: Delta = 34'sb0000000000000000000000011111100000;
		4231: Delta = 34'sb1111111111111111111111011111100000;
		4128: Delta = 34'sb0000000000000000000001000000100000;
		2247: Delta = 34'sb1111111111111111111111000000100000;
		4064: Delta = 34'sb0000000000000000000000111111100000;
		2183: Delta = 34'sb1111111111111111111110111111100000;
		1913: Delta = 34'sb0000000000000000000010000000100000;
		4462: Delta = 34'sb1111111111111111111110000000100000;
		1849: Delta = 34'sb0000000000000000000001111111100000;
		4398: Delta = 34'sb1111111111111111111101111111100000;
		3794: Delta = 34'sb0000000000000000000100000000100000;
		2581: Delta = 34'sb1111111111111111111100000000100000;
		3730: Delta = 34'sb0000000000000000000011111111100000;
		2517: Delta = 34'sb1111111111111111111011111111100000;
		1245: Delta = 34'sb0000000000000000001000000000100000;
		5130: Delta = 34'sb1111111111111111111000000000100000;
		1181: Delta = 34'sb0000000000000000000111111111100000;
		5066: Delta = 34'sb1111111111111111110111111111100000;
		2458: Delta = 34'sb0000000000000000010000000000100000;
		3917: Delta = 34'sb1111111111111111110000000000100000;
		2394: Delta = 34'sb0000000000000000001111111111100000;
		3853: Delta = 34'sb1111111111111111101111111111100000;
		4884: Delta = 34'sb0000000000000000100000000000100000;
		1491: Delta = 34'sb1111111111111111100000000000100000;
		4820: Delta = 34'sb0000000000000000011111111111100000;
		1427: Delta = 34'sb1111111111111111011111111111100000;
		3425: Delta = 34'sb0000000000000001000000000000100000;
		2950: Delta = 34'sb1111111111111111000000000000100000;
		3361: Delta = 34'sb0000000000000000111111111111100000;
		2886: Delta = 34'sb1111111111111110111111111111100000;
		507: Delta = 34'sb0000000000000010000000000000100000;
		5868: Delta = 34'sb1111111111111110000000000000100000;
		443: Delta = 34'sb0000000000000001111111111111100000;
		5804: Delta = 34'sb1111111111111101111111111111100000;
		982: Delta = 34'sb0000000000000100000000000000100000;
		5393: Delta = 34'sb1111111111111100000000000000100000;
		918: Delta = 34'sb0000000000000011111111111111100000;
		5329: Delta = 34'sb1111111111111011111111111111100000;
		1932: Delta = 34'sb0000000000001000000000000000100000;
		4443: Delta = 34'sb1111111111111000000000000000100000;
		1868: Delta = 34'sb0000000000000111111111111111100000;
		4379: Delta = 34'sb1111111111110111111111111111100000;
		3832: Delta = 34'sb0000000000010000000000000000100000;
		2543: Delta = 34'sb1111111111110000000000000000100000;
		3768: Delta = 34'sb0000000000001111111111111111100000;
		2479: Delta = 34'sb1111111111101111111111111111100000;
		1321: Delta = 34'sb0000000000100000000000000000100000;
		5054: Delta = 34'sb1111111111100000000000000000100000;
		1257: Delta = 34'sb0000000000011111111111111111100000;
		4990: Delta = 34'sb1111111111011111111111111111100000;
		2610: Delta = 34'sb0000000001000000000000000000100000;
		3765: Delta = 34'sb1111111111000000000000000000100000;
		2546: Delta = 34'sb0000000000111111111111111111100000;
		3701: Delta = 34'sb1111111110111111111111111111100000;
		5188: Delta = 34'sb0000000010000000000000000000100000;
		1187: Delta = 34'sb1111111110000000000000000000100000;
		5124: Delta = 34'sb0000000001111111111111111111100000;
		1123: Delta = 34'sb1111111101111111111111111111100000;
		4033: Delta = 34'sb0000000100000000000000000000100000;
		2342: Delta = 34'sb1111111100000000000000000000100000;
		3969: Delta = 34'sb0000000011111111111111111111100000;
		2278: Delta = 34'sb1111111011111111111111111111100000;
		1723: Delta = 34'sb0000001000000000000000000000100000;
		4652: Delta = 34'sb1111111000000000000000000000100000;
		1659: Delta = 34'sb0000000111111111111111111111100000;
		4588: Delta = 34'sb1111110111111111111111111111100000;
		3414: Delta = 34'sb0000010000000000000000000000100000;
		2961: Delta = 34'sb1111110000000000000000000000100000;
		3350: Delta = 34'sb0000001111111111111111111111100000;
		2897: Delta = 34'sb1111101111111111111111111111100000;
		485: Delta = 34'sb0000100000000000000000000000100000;
		5890: Delta = 34'sb1111100000000000000000000000100000;
		421: Delta = 34'sb0000011111111111111111111111100000;
		5826: Delta = 34'sb1111011111111111111111111111100000;
		938: Delta = 34'sb0001000000000000000000000000100000;
		5437: Delta = 34'sb1111000000000000000000000000100000;
		874: Delta = 34'sb0000111111111111111111111111100000;
		5373: Delta = 34'sb1110111111111111111111111111100000;
		1844: Delta = 34'sb0010000000000000000000000000100000;
		4531: Delta = 34'sb1110000000000000000000000000100000;
		1780: Delta = 34'sb0001111111111111111111111111100000;
		4467: Delta = 34'sb1101111111111111111111111111100000;
		3656: Delta = 34'sb0100000000000000000000000000100000;
		2719: Delta = 34'sb1100000000000000000000000000100000;
		3592: Delta = 34'sb0011111111111111111111111111100000;
		2655: Delta = 34'sb1011111111111111111111111111100000;
		192: Delta = 34'sb0000000000000000000000000011000000;
		6119: Delta = 34'sb1111111111111111111111111101000000;
		320: Delta = 34'sb0000000000000000000000000101000000;
		5991: Delta = 34'sb1111111111111111111111111011000000;
		576: Delta = 34'sb0000000000000000000000001001000000;
		5863: Delta = 34'sb1111111111111111111111111001000000;
		448: Delta = 34'sb0000000000000000000000000111000000;
		5735: Delta = 34'sb1111111111111111111111110111000000;
		1088: Delta = 34'sb0000000000000000000000010001000000;
		5351: Delta = 34'sb1111111111111111111111110001000000;
		960: Delta = 34'sb0000000000000000000000001111000000;
		5223: Delta = 34'sb1111111111111111111111101111000000;
		2112: Delta = 34'sb0000000000000000000000100001000000;
		4327: Delta = 34'sb1111111111111111111111100001000000;
		1984: Delta = 34'sb0000000000000000000000011111000000;
		4199: Delta = 34'sb1111111111111111111111011111000000;
		4160: Delta = 34'sb0000000000000000000001000001000000;
		2279: Delta = 34'sb1111111111111111111111000001000000;
		4032: Delta = 34'sb0000000000000000000000111111000000;
		2151: Delta = 34'sb1111111111111111111110111111000000;
		1945: Delta = 34'sb0000000000000000000010000001000000;
		4494: Delta = 34'sb1111111111111111111110000001000000;
		1817: Delta = 34'sb0000000000000000000001111111000000;
		4366: Delta = 34'sb1111111111111111111101111111000000;
		3826: Delta = 34'sb0000000000000000000100000001000000;
		2613: Delta = 34'sb1111111111111111111100000001000000;
		3698: Delta = 34'sb0000000000000000000011111111000000;
		2485: Delta = 34'sb1111111111111111111011111111000000;
		1277: Delta = 34'sb0000000000000000001000000001000000;
		5162: Delta = 34'sb1111111111111111111000000001000000;
		1149: Delta = 34'sb0000000000000000000111111111000000;
		5034: Delta = 34'sb1111111111111111110111111111000000;
		2490: Delta = 34'sb0000000000000000010000000001000000;
		3949: Delta = 34'sb1111111111111111110000000001000000;
		2362: Delta = 34'sb0000000000000000001111111111000000;
		3821: Delta = 34'sb1111111111111111101111111111000000;
		4916: Delta = 34'sb0000000000000000100000000001000000;
		1523: Delta = 34'sb1111111111111111100000000001000000;
		4788: Delta = 34'sb0000000000000000011111111111000000;
		1395: Delta = 34'sb1111111111111111011111111111000000;
		3457: Delta = 34'sb0000000000000001000000000001000000;
		2982: Delta = 34'sb1111111111111111000000000001000000;
		3329: Delta = 34'sb0000000000000000111111111111000000;
		2854: Delta = 34'sb1111111111111110111111111111000000;
		539: Delta = 34'sb0000000000000010000000000001000000;
		5900: Delta = 34'sb1111111111111110000000000001000000;
		411: Delta = 34'sb0000000000000001111111111111000000;
		5772: Delta = 34'sb1111111111111101111111111111000000;
		1014: Delta = 34'sb0000000000000100000000000001000000;
		5425: Delta = 34'sb1111111111111100000000000001000000;
		886: Delta = 34'sb0000000000000011111111111111000000;
		5297: Delta = 34'sb1111111111111011111111111111000000;
		1964: Delta = 34'sb0000000000001000000000000001000000;
		4475: Delta = 34'sb1111111111111000000000000001000000;
		1836: Delta = 34'sb0000000000000111111111111111000000;
		4347: Delta = 34'sb1111111111110111111111111111000000;
		3864: Delta = 34'sb0000000000010000000000000001000000;
		2575: Delta = 34'sb1111111111110000000000000001000000;
		3736: Delta = 34'sb0000000000001111111111111111000000;
		2447: Delta = 34'sb1111111111101111111111111111000000;
		1353: Delta = 34'sb0000000000100000000000000001000000;
		5086: Delta = 34'sb1111111111100000000000000001000000;
		1225: Delta = 34'sb0000000000011111111111111111000000;
		4958: Delta = 34'sb1111111111011111111111111111000000;
		2642: Delta = 34'sb0000000001000000000000000001000000;
		3797: Delta = 34'sb1111111111000000000000000001000000;
		2514: Delta = 34'sb0000000000111111111111111111000000;
		3669: Delta = 34'sb1111111110111111111111111111000000;
		5220: Delta = 34'sb0000000010000000000000000001000000;
		1219: Delta = 34'sb1111111110000000000000000001000000;
		5092: Delta = 34'sb0000000001111111111111111111000000;
		1091: Delta = 34'sb1111111101111111111111111111000000;
		4065: Delta = 34'sb0000000100000000000000000001000000;
		2374: Delta = 34'sb1111111100000000000000000001000000;
		3937: Delta = 34'sb0000000011111111111111111111000000;
		2246: Delta = 34'sb1111111011111111111111111111000000;
		1755: Delta = 34'sb0000001000000000000000000001000000;
		4684: Delta = 34'sb1111111000000000000000000001000000;
		1627: Delta = 34'sb0000000111111111111111111111000000;
		4556: Delta = 34'sb1111110111111111111111111111000000;
		3446: Delta = 34'sb0000010000000000000000000001000000;
		2993: Delta = 34'sb1111110000000000000000000001000000;
		3318: Delta = 34'sb0000001111111111111111111111000000;
		2865: Delta = 34'sb1111101111111111111111111111000000;
		517: Delta = 34'sb0000100000000000000000000001000000;
		5922: Delta = 34'sb1111100000000000000000000001000000;
		389: Delta = 34'sb0000011111111111111111111111000000;
		5794: Delta = 34'sb1111011111111111111111111111000000;
		970: Delta = 34'sb0001000000000000000000000001000000;
		5469: Delta = 34'sb1111000000000000000000000001000000;
		842: Delta = 34'sb0000111111111111111111111111000000;
		5341: Delta = 34'sb1110111111111111111111111111000000;
		1876: Delta = 34'sb0010000000000000000000000001000000;
		4563: Delta = 34'sb1110000000000000000000000001000000;
		1748: Delta = 34'sb0001111111111111111111111111000000;
		4435: Delta = 34'sb1101111111111111111111111111000000;
		3688: Delta = 34'sb0100000000000000000000000001000000;
		2751: Delta = 34'sb1100000000000000000000000001000000;
		3560: Delta = 34'sb0011111111111111111111111111000000;
		2623: Delta = 34'sb1011111111111111111111111111000000;
		384: Delta = 34'sb0000000000000000000000000110000000;
		5927: Delta = 34'sb1111111111111111111111111010000000;
		640: Delta = 34'sb0000000000000000000000001010000000;
		5671: Delta = 34'sb1111111111111111111111110110000000;
		1152: Delta = 34'sb0000000000000000000000010010000000;
		5415: Delta = 34'sb1111111111111111111111110010000000;
		896: Delta = 34'sb0000000000000000000000001110000000;
		5159: Delta = 34'sb1111111111111111111111101110000000;
		2176: Delta = 34'sb0000000000000000000000100010000000;
		4391: Delta = 34'sb1111111111111111111111100010000000;
		1920: Delta = 34'sb0000000000000000000000011110000000;
		4135: Delta = 34'sb1111111111111111111111011110000000;
		4224: Delta = 34'sb0000000000000000000001000010000000;
		2343: Delta = 34'sb1111111111111111111111000010000000;
		3968: Delta = 34'sb0000000000000000000000111110000000;
		2087: Delta = 34'sb1111111111111111111110111110000000;
		2009: Delta = 34'sb0000000000000000000010000010000000;
		4558: Delta = 34'sb1111111111111111111110000010000000;
		1753: Delta = 34'sb0000000000000000000001111110000000;
		4302: Delta = 34'sb1111111111111111111101111110000000;
		3890: Delta = 34'sb0000000000000000000100000010000000;
		2677: Delta = 34'sb1111111111111111111100000010000000;
		3634: Delta = 34'sb0000000000000000000011111110000000;
		2421: Delta = 34'sb1111111111111111111011111110000000;
		1341: Delta = 34'sb0000000000000000001000000010000000;
		5226: Delta = 34'sb1111111111111111111000000010000000;
		1085: Delta = 34'sb0000000000000000000111111110000000;
		4970: Delta = 34'sb1111111111111111110111111110000000;
		2554: Delta = 34'sb0000000000000000010000000010000000;
		4013: Delta = 34'sb1111111111111111110000000010000000;
		2298: Delta = 34'sb0000000000000000001111111110000000;
		3757: Delta = 34'sb1111111111111111101111111110000000;
		4980: Delta = 34'sb0000000000000000100000000010000000;
		1587: Delta = 34'sb1111111111111111100000000010000000;
		4724: Delta = 34'sb0000000000000000011111111110000000;
		1331: Delta = 34'sb1111111111111111011111111110000000;
		3521: Delta = 34'sb0000000000000001000000000010000000;
		3046: Delta = 34'sb1111111111111111000000000010000000;
		3265: Delta = 34'sb0000000000000000111111111110000000;
		2790: Delta = 34'sb1111111111111110111111111110000000;
		603: Delta = 34'sb0000000000000010000000000010000000;
		5964: Delta = 34'sb1111111111111110000000000010000000;
		347: Delta = 34'sb0000000000000001111111111110000000;
		5708: Delta = 34'sb1111111111111101111111111110000000;
		1078: Delta = 34'sb0000000000000100000000000010000000;
		5489: Delta = 34'sb1111111111111100000000000010000000;
		822: Delta = 34'sb0000000000000011111111111110000000;
		5233: Delta = 34'sb1111111111111011111111111110000000;
		2028: Delta = 34'sb0000000000001000000000000010000000;
		4539: Delta = 34'sb1111111111111000000000000010000000;
		1772: Delta = 34'sb0000000000000111111111111110000000;
		4283: Delta = 34'sb1111111111110111111111111110000000;
		3928: Delta = 34'sb0000000000010000000000000010000000;
		2639: Delta = 34'sb1111111111110000000000000010000000;
		3672: Delta = 34'sb0000000000001111111111111110000000;
		2383: Delta = 34'sb1111111111101111111111111110000000;
		1417: Delta = 34'sb0000000000100000000000000010000000;
		5150: Delta = 34'sb1111111111100000000000000010000000;
		1161: Delta = 34'sb0000000000011111111111111110000000;
		4894: Delta = 34'sb1111111111011111111111111110000000;
		2706: Delta = 34'sb0000000001000000000000000010000000;
		3861: Delta = 34'sb1111111111000000000000000010000000;
		2450: Delta = 34'sb0000000000111111111111111110000000;
		3605: Delta = 34'sb1111111110111111111111111110000000;
		5284: Delta = 34'sb0000000010000000000000000010000000;
		1283: Delta = 34'sb1111111110000000000000000010000000;
		5028: Delta = 34'sb0000000001111111111111111110000000;
		1027: Delta = 34'sb1111111101111111111111111110000000;
		4129: Delta = 34'sb0000000100000000000000000010000000;
		2438: Delta = 34'sb1111111100000000000000000010000000;
		3873: Delta = 34'sb0000000011111111111111111110000000;
		2182: Delta = 34'sb1111111011111111111111111110000000;
		1819: Delta = 34'sb0000001000000000000000000010000000;
		4748: Delta = 34'sb1111111000000000000000000010000000;
		1563: Delta = 34'sb0000000111111111111111111110000000;
		4492: Delta = 34'sb1111110111111111111111111110000000;
		3510: Delta = 34'sb0000010000000000000000000010000000;
		3057: Delta = 34'sb1111110000000000000000000010000000;
		3254: Delta = 34'sb0000001111111111111111111110000000;
		2801: Delta = 34'sb1111101111111111111111111110000000;
		581: Delta = 34'sb0000100000000000000000000010000000;
		5986: Delta = 34'sb1111100000000000000000000010000000;
		325: Delta = 34'sb0000011111111111111111111110000000;
		5730: Delta = 34'sb1111011111111111111111111110000000;
		1034: Delta = 34'sb0001000000000000000000000010000000;
		5533: Delta = 34'sb1111000000000000000000000010000000;
		778: Delta = 34'sb0000111111111111111111111110000000;
		5277: Delta = 34'sb1110111111111111111111111110000000;
		1940: Delta = 34'sb0010000000000000000000000010000000;
		4627: Delta = 34'sb1110000000000000000000000010000000;
		1684: Delta = 34'sb0001111111111111111111111110000000;
		4371: Delta = 34'sb1101111111111111111111111110000000;
		3752: Delta = 34'sb0100000000000000000000000010000000;
		2815: Delta = 34'sb1100000000000000000000000010000000;
		3496: Delta = 34'sb0011111111111111111111111110000000;
		2559: Delta = 34'sb1011111111111111111111111110000000;
		768: Delta = 34'sb0000000000000000000000001100000000;
		5543: Delta = 34'sb1111111111111111111111110100000000;
		1280: Delta = 34'sb0000000000000000000000010100000000;
		5031: Delta = 34'sb1111111111111111111111101100000000;
		2304: Delta = 34'sb0000000000000000000000100100000000;
		4519: Delta = 34'sb1111111111111111111111100100000000;
		1792: Delta = 34'sb0000000000000000000000011100000000;
		4007: Delta = 34'sb1111111111111111111111011100000000;
		4352: Delta = 34'sb0000000000000000000001000100000000;
		2471: Delta = 34'sb1111111111111111111111000100000000;
		3840: Delta = 34'sb0000000000000000000000111100000000;
		1959: Delta = 34'sb1111111111111111111110111100000000;
		2137: Delta = 34'sb0000000000000000000010000100000000;
		4686: Delta = 34'sb1111111111111111111110000100000000;
		1625: Delta = 34'sb0000000000000000000001111100000000;
		4174: Delta = 34'sb1111111111111111111101111100000000;
		4018: Delta = 34'sb0000000000000000000100000100000000;
		2805: Delta = 34'sb1111111111111111111100000100000000;
		3506: Delta = 34'sb0000000000000000000011111100000000;
		2293: Delta = 34'sb1111111111111111111011111100000000;
		1469: Delta = 34'sb0000000000000000001000000100000000;
		5354: Delta = 34'sb1111111111111111111000000100000000;
		957: Delta = 34'sb0000000000000000000111111100000000;
		4842: Delta = 34'sb1111111111111111110111111100000000;
		2682: Delta = 34'sb0000000000000000010000000100000000;
		4141: Delta = 34'sb1111111111111111110000000100000000;
		2170: Delta = 34'sb0000000000000000001111111100000000;
		3629: Delta = 34'sb1111111111111111101111111100000000;
		5108: Delta = 34'sb0000000000000000100000000100000000;
		1715: Delta = 34'sb1111111111111111100000000100000000;
		4596: Delta = 34'sb0000000000000000011111111100000000;
		1203: Delta = 34'sb1111111111111111011111111100000000;
		3649: Delta = 34'sb0000000000000001000000000100000000;
		3174: Delta = 34'sb1111111111111111000000000100000000;
		3137: Delta = 34'sb0000000000000000111111111100000000;
		2662: Delta = 34'sb1111111111111110111111111100000000;
		731: Delta = 34'sb0000000000000010000000000100000000;
		6092: Delta = 34'sb1111111111111110000000000100000000;
		219: Delta = 34'sb0000000000000001111111111100000000;
		5580: Delta = 34'sb1111111111111101111111111100000000;
		1206: Delta = 34'sb0000000000000100000000000100000000;
		5617: Delta = 34'sb1111111111111100000000000100000000;
		694: Delta = 34'sb0000000000000011111111111100000000;
		5105: Delta = 34'sb1111111111111011111111111100000000;
		2156: Delta = 34'sb0000000000001000000000000100000000;
		4667: Delta = 34'sb1111111111111000000000000100000000;
		1644: Delta = 34'sb0000000000000111111111111100000000;
		4155: Delta = 34'sb1111111111110111111111111100000000;
		4056: Delta = 34'sb0000000000010000000000000100000000;
		2767: Delta = 34'sb1111111111110000000000000100000000;
		3544: Delta = 34'sb0000000000001111111111111100000000;
		2255: Delta = 34'sb1111111111101111111111111100000000;
		1545: Delta = 34'sb0000000000100000000000000100000000;
		5278: Delta = 34'sb1111111111100000000000000100000000;
		1033: Delta = 34'sb0000000000011111111111111100000000;
		4766: Delta = 34'sb1111111111011111111111111100000000;
		2834: Delta = 34'sb0000000001000000000000000100000000;
		3989: Delta = 34'sb1111111111000000000000000100000000;
		2322: Delta = 34'sb0000000000111111111111111100000000;
		3477: Delta = 34'sb1111111110111111111111111100000000;
		5412: Delta = 34'sb0000000010000000000000000100000000;
		1411: Delta = 34'sb1111111110000000000000000100000000;
		4900: Delta = 34'sb0000000001111111111111111100000000;
		899: Delta = 34'sb1111111101111111111111111100000000;
		4257: Delta = 34'sb0000000100000000000000000100000000;
		2566: Delta = 34'sb1111111100000000000000000100000000;
		3745: Delta = 34'sb0000000011111111111111111100000000;
		2054: Delta = 34'sb1111111011111111111111111100000000;
		1947: Delta = 34'sb0000001000000000000000000100000000;
		4876: Delta = 34'sb1111111000000000000000000100000000;
		1435: Delta = 34'sb0000000111111111111111111100000000;
		4364: Delta = 34'sb1111110111111111111111111100000000;
		3638: Delta = 34'sb0000010000000000000000000100000000;
		3185: Delta = 34'sb1111110000000000000000000100000000;
		3126: Delta = 34'sb0000001111111111111111111100000000;
		2673: Delta = 34'sb1111101111111111111111111100000000;
		709: Delta = 34'sb0000100000000000000000000100000000;
		6114: Delta = 34'sb1111100000000000000000000100000000;
		197: Delta = 34'sb0000011111111111111111111100000000;
		5602: Delta = 34'sb1111011111111111111111111100000000;
		1162: Delta = 34'sb0001000000000000000000000100000000;
		5661: Delta = 34'sb1111000000000000000000000100000000;
		650: Delta = 34'sb0000111111111111111111111100000000;
		5149: Delta = 34'sb1110111111111111111111111100000000;
		2068: Delta = 34'sb0010000000000000000000000100000000;
		4755: Delta = 34'sb1110000000000000000000000100000000;
		1556: Delta = 34'sb0001111111111111111111111100000000;
		4243: Delta = 34'sb1101111111111111111111111100000000;
		3880: Delta = 34'sb0100000000000000000000000100000000;
		2943: Delta = 34'sb1100000000000000000000000100000000;
		3368: Delta = 34'sb0011111111111111111111111100000000;
		2431: Delta = 34'sb1011111111111111111111111100000000;
		1536: Delta = 34'sb0000000000000000000000011000000000;
		4775: Delta = 34'sb1111111111111111111111101000000000;
		2560: Delta = 34'sb0000000000000000000000101000000000;
		3751: Delta = 34'sb1111111111111111111111011000000000;
		4608: Delta = 34'sb0000000000000000000001001000000000;
		2727: Delta = 34'sb1111111111111111111111001000000000;
		3584: Delta = 34'sb0000000000000000000000111000000000;
		1703: Delta = 34'sb1111111111111111111110111000000000;
		2393: Delta = 34'sb0000000000000000000010001000000000;
		4942: Delta = 34'sb1111111111111111111110001000000000;
		1369: Delta = 34'sb0000000000000000000001111000000000;
		3918: Delta = 34'sb1111111111111111111101111000000000;
		4274: Delta = 34'sb0000000000000000000100001000000000;
		3061: Delta = 34'sb1111111111111111111100001000000000;
		3250: Delta = 34'sb0000000000000000000011111000000000;
		2037: Delta = 34'sb1111111111111111111011111000000000;
		1725: Delta = 34'sb0000000000000000001000001000000000;
		5610: Delta = 34'sb1111111111111111111000001000000000;
		701: Delta = 34'sb0000000000000000000111111000000000;
		4586: Delta = 34'sb1111111111111111110111111000000000;
		2938: Delta = 34'sb0000000000000000010000001000000000;
		4397: Delta = 34'sb1111111111111111110000001000000000;
		1914: Delta = 34'sb0000000000000000001111111000000000;
		3373: Delta = 34'sb1111111111111111101111111000000000;
		5364: Delta = 34'sb0000000000000000100000001000000000;
		1971: Delta = 34'sb1111111111111111100000001000000000;
		4340: Delta = 34'sb0000000000000000011111111000000000;
		947: Delta = 34'sb1111111111111111011111111000000000;
		3905: Delta = 34'sb0000000000000001000000001000000000;
		3430: Delta = 34'sb1111111111111111000000001000000000;
		2881: Delta = 34'sb0000000000000000111111111000000000;
		2406: Delta = 34'sb1111111111111110111111111000000000;
		987: Delta = 34'sb0000000000000010000000001000000000;
		37: Delta = 34'sb1111111111111110000000001000000000;
		6274: Delta = 34'sb0000000000000001111111111000000000;
		5324: Delta = 34'sb1111111111111101111111111000000000;
		1462: Delta = 34'sb0000000000000100000000001000000000;
		5873: Delta = 34'sb1111111111111100000000001000000000;
		438: Delta = 34'sb0000000000000011111111111000000000;
		4849: Delta = 34'sb1111111111111011111111111000000000;
		2412: Delta = 34'sb0000000000001000000000001000000000;
		4923: Delta = 34'sb1111111111111000000000001000000000;
		1388: Delta = 34'sb0000000000000111111111111000000000;
		3899: Delta = 34'sb1111111111110111111111111000000000;
		4312: Delta = 34'sb0000000000010000000000001000000000;
		3023: Delta = 34'sb1111111111110000000000001000000000;
		3288: Delta = 34'sb0000000000001111111111111000000000;
		1999: Delta = 34'sb1111111111101111111111111000000000;
		1801: Delta = 34'sb0000000000100000000000001000000000;
		5534: Delta = 34'sb1111111111100000000000001000000000;
		777: Delta = 34'sb0000000000011111111111111000000000;
		4510: Delta = 34'sb1111111111011111111111111000000000;
		3090: Delta = 34'sb0000000001000000000000001000000000;
		4245: Delta = 34'sb1111111111000000000000001000000000;
		2066: Delta = 34'sb0000000000111111111111111000000000;
		3221: Delta = 34'sb1111111110111111111111111000000000;
		5668: Delta = 34'sb0000000010000000000000001000000000;
		1667: Delta = 34'sb1111111110000000000000001000000000;
		4644: Delta = 34'sb0000000001111111111111111000000000;
		643: Delta = 34'sb1111111101111111111111111000000000;
		4513: Delta = 34'sb0000000100000000000000001000000000;
		2822: Delta = 34'sb1111111100000000000000001000000000;
		3489: Delta = 34'sb0000000011111111111111111000000000;
		1798: Delta = 34'sb1111111011111111111111111000000000;
		2203: Delta = 34'sb0000001000000000000000001000000000;
		5132: Delta = 34'sb1111111000000000000000001000000000;
		1179: Delta = 34'sb0000000111111111111111111000000000;
		4108: Delta = 34'sb1111110111111111111111111000000000;
		3894: Delta = 34'sb0000010000000000000000001000000000;
		3441: Delta = 34'sb1111110000000000000000001000000000;
		2870: Delta = 34'sb0000001111111111111111111000000000;
		2417: Delta = 34'sb1111101111111111111111111000000000;
		965: Delta = 34'sb0000100000000000000000001000000000;
		59: Delta = 34'sb1111100000000000000000001000000000;
		6252: Delta = 34'sb0000011111111111111111111000000000;
		5346: Delta = 34'sb1111011111111111111111111000000000;
		1418: Delta = 34'sb0001000000000000000000001000000000;
		5917: Delta = 34'sb1111000000000000000000001000000000;
		394: Delta = 34'sb0000111111111111111111111000000000;
		4893: Delta = 34'sb1110111111111111111111111000000000;
		2324: Delta = 34'sb0010000000000000000000001000000000;
		5011: Delta = 34'sb1110000000000000000000001000000000;
		1300: Delta = 34'sb0001111111111111111111111000000000;
		3987: Delta = 34'sb1101111111111111111111111000000000;
		4136: Delta = 34'sb0100000000000000000000001000000000;
		3199: Delta = 34'sb1100000000000000000000001000000000;
		3112: Delta = 34'sb0011111111111111111111111000000000;
		2175: Delta = 34'sb1011111111111111111111111000000000;
		3072: Delta = 34'sb0000000000000000000000110000000000;
		3239: Delta = 34'sb1111111111111111111111010000000000;
		5120: Delta = 34'sb0000000000000000000001010000000000;
		1191: Delta = 34'sb1111111111111111111110110000000000;
		2905: Delta = 34'sb0000000000000000000010010000000000;
		5454: Delta = 34'sb1111111111111111111110010000000000;
		857: Delta = 34'sb0000000000000000000001110000000000;
		3406: Delta = 34'sb1111111111111111111101110000000000;
		4786: Delta = 34'sb0000000000000000000100010000000000;
		3573: Delta = 34'sb1111111111111111111100010000000000;
		2738: Delta = 34'sb0000000000000000000011110000000000;
		1525: Delta = 34'sb1111111111111111111011110000000000;
		2237: Delta = 34'sb0000000000000000001000010000000000;
		6122: Delta = 34'sb1111111111111111111000010000000000;
		189: Delta = 34'sb0000000000000000000111110000000000;
		4074: Delta = 34'sb1111111111111111110111110000000000;
		3450: Delta = 34'sb0000000000000000010000010000000000;
		4909: Delta = 34'sb1111111111111111110000010000000000;
		1402: Delta = 34'sb0000000000000000001111110000000000;
		2861: Delta = 34'sb1111111111111111101111110000000000;
		5876: Delta = 34'sb0000000000000000100000010000000000;
		2483: Delta = 34'sb1111111111111111100000010000000000;
		3828: Delta = 34'sb0000000000000000011111110000000000;
		435: Delta = 34'sb1111111111111111011111110000000000;
		4417: Delta = 34'sb0000000000000001000000010000000000;
		3942: Delta = 34'sb1111111111111111000000010000000000;
		2369: Delta = 34'sb0000000000000000111111110000000000;
		1894: Delta = 34'sb1111111111111110111111110000000000;
		1499: Delta = 34'sb0000000000000010000000010000000000;
		549: Delta = 34'sb1111111111111110000000010000000000;
		5762: Delta = 34'sb0000000000000001111111110000000000;
		4812: Delta = 34'sb1111111111111101111111110000000000;
		1974: Delta = 34'sb0000000000000100000000010000000000;
		74: Delta = 34'sb1111111111111100000000010000000000;
		6237: Delta = 34'sb0000000000000011111111110000000000;
		4337: Delta = 34'sb1111111111111011111111110000000000;
		2924: Delta = 34'sb0000000000001000000000010000000000;
		5435: Delta = 34'sb1111111111111000000000010000000000;
		876: Delta = 34'sb0000000000000111111111110000000000;
		3387: Delta = 34'sb1111111111110111111111110000000000;
		4824: Delta = 34'sb0000000000010000000000010000000000;
		3535: Delta = 34'sb1111111111110000000000010000000000;
		2776: Delta = 34'sb0000000000001111111111110000000000;
		1487: Delta = 34'sb1111111111101111111111110000000000;
		2313: Delta = 34'sb0000000000100000000000010000000000;
		6046: Delta = 34'sb1111111111100000000000010000000000;
		265: Delta = 34'sb0000000000011111111111110000000000;
		3998: Delta = 34'sb1111111111011111111111110000000000;
		3602: Delta = 34'sb0000000001000000000000010000000000;
		4757: Delta = 34'sb1111111111000000000000010000000000;
		1554: Delta = 34'sb0000000000111111111111110000000000;
		2709: Delta = 34'sb1111111110111111111111110000000000;
		6180: Delta = 34'sb0000000010000000000000010000000000;
		2179: Delta = 34'sb1111111110000000000000010000000000;
		4132: Delta = 34'sb0000000001111111111111110000000000;
		131: Delta = 34'sb1111111101111111111111110000000000;
		5025: Delta = 34'sb0000000100000000000000010000000000;
		3334: Delta = 34'sb1111111100000000000000010000000000;
		2977: Delta = 34'sb0000000011111111111111110000000000;
		1286: Delta = 34'sb1111111011111111111111110000000000;
		2715: Delta = 34'sb0000001000000000000000010000000000;
		5644: Delta = 34'sb1111111000000000000000010000000000;
		667: Delta = 34'sb0000000111111111111111110000000000;
		3596: Delta = 34'sb1111110111111111111111110000000000;
		4406: Delta = 34'sb0000010000000000000000010000000000;
		3953: Delta = 34'sb1111110000000000000000010000000000;
		2358: Delta = 34'sb0000001111111111111111110000000000;
		1905: Delta = 34'sb1111101111111111111111110000000000;
		1477: Delta = 34'sb0000100000000000000000010000000000;
		571: Delta = 34'sb1111100000000000000000010000000000;
		5740: Delta = 34'sb0000011111111111111111110000000000;
		4834: Delta = 34'sb1111011111111111111111110000000000;
		1930: Delta = 34'sb0001000000000000000000010000000000;
		118: Delta = 34'sb1111000000000000000000010000000000;
		6193: Delta = 34'sb0000111111111111111111110000000000;
		4381: Delta = 34'sb1110111111111111111111110000000000;
		2836: Delta = 34'sb0010000000000000000000010000000000;
		5523: Delta = 34'sb1110000000000000000000010000000000;
		788: Delta = 34'sb0001111111111111111111110000000000;
		3475: Delta = 34'sb1101111111111111111111110000000000;
		4648: Delta = 34'sb0100000000000000000000010000000000;
		3711: Delta = 34'sb1100000000000000000000010000000000;
		2600: Delta = 34'sb0011111111111111111111110000000000;
		1663: Delta = 34'sb1011111111111111111111110000000000;
		6144: Delta = 34'sb0000000000000000000001100000000000;
		167: Delta = 34'sb1111111111111111111110100000000000;
		3929: Delta = 34'sb0000000000000000000010100000000000;
		2382: Delta = 34'sb1111111111111111111101100000000000;
		5810: Delta = 34'sb0000000000000000000100100000000000;
		4597: Delta = 34'sb1111111111111111111100100000000000;
		1714: Delta = 34'sb0000000000000000000011100000000000;
		501: Delta = 34'sb1111111111111111111011100000000000;
		3261: Delta = 34'sb0000000000000000001000100000000000;
		835: Delta = 34'sb1111111111111111111000100000000000;
		5476: Delta = 34'sb0000000000000000000111100000000000;
		3050: Delta = 34'sb1111111111111111110111100000000000;
		4474: Delta = 34'sb0000000000000000010000100000000000;
		5933: Delta = 34'sb1111111111111111110000100000000000;
		378: Delta = 34'sb0000000000000000001111100000000000;
		1837: Delta = 34'sb1111111111111111101111100000000000;
		589: Delta = 34'sb0000000000000000100000100000000000;
		3507: Delta = 34'sb1111111111111111100000100000000000;
		2804: Delta = 34'sb0000000000000000011111100000000000;
		5722: Delta = 34'sb1111111111111111011111100000000000;
		5441: Delta = 34'sb0000000000000001000000100000000000;
		4966: Delta = 34'sb1111111111111111000000100000000000;
		1345: Delta = 34'sb0000000000000000111111100000000000;
		870: Delta = 34'sb1111111111111110111111100000000000;
		2523: Delta = 34'sb0000000000000010000000100000000000;
		1573: Delta = 34'sb1111111111111110000000100000000000;
		4738: Delta = 34'sb0000000000000001111111100000000000;
		3788: Delta = 34'sb1111111111111101111111100000000000;
		2998: Delta = 34'sb0000000000000100000000100000000000;
		1098: Delta = 34'sb1111111111111100000000100000000000;
		5213: Delta = 34'sb0000000000000011111111100000000000;
		3313: Delta = 34'sb1111111111111011111111100000000000;
		3948: Delta = 34'sb0000000000001000000000100000000000;
		148: Delta = 34'sb1111111111111000000000100000000000;
		6163: Delta = 34'sb0000000000000111111111100000000000;
		2363: Delta = 34'sb1111111111110111111111100000000000;
		5848: Delta = 34'sb0000000000010000000000100000000000;
		4559: Delta = 34'sb1111111111110000000000100000000000;
		1752: Delta = 34'sb0000000000001111111111100000000000;
		463: Delta = 34'sb1111111111101111111111100000000000;
		3337: Delta = 34'sb0000000000100000000000100000000000;
		759: Delta = 34'sb1111111111100000000000100000000000;
		5552: Delta = 34'sb0000000000011111111111100000000000;
		2974: Delta = 34'sb1111111111011111111111100000000000;
		4626: Delta = 34'sb0000000001000000000000100000000000;
		5781: Delta = 34'sb1111111111000000000000100000000000;
		530: Delta = 34'sb0000000000111111111111100000000000;
		1685: Delta = 34'sb1111111110111111111111100000000000;
		893: Delta = 34'sb0000000010000000000000100000000000;
		3203: Delta = 34'sb1111111110000000000000100000000000;
		3108: Delta = 34'sb0000000001111111111111100000000000;
		5418: Delta = 34'sb1111111101111111111111100000000000;
		6049: Delta = 34'sb0000000100000000000000100000000000;
		4358: Delta = 34'sb1111111100000000000000100000000000;
		1953: Delta = 34'sb0000000011111111111111100000000000;
		262: Delta = 34'sb1111111011111111111111100000000000;
		3739: Delta = 34'sb0000001000000000000000100000000000;
		357: Delta = 34'sb1111111000000000000000100000000000;
		5954: Delta = 34'sb0000000111111111111111100000000000;
		2572: Delta = 34'sb1111110111111111111111100000000000;
		5430: Delta = 34'sb0000010000000000000000100000000000;
		4977: Delta = 34'sb1111110000000000000000100000000000;
		1334: Delta = 34'sb0000001111111111111111100000000000;
		881: Delta = 34'sb1111101111111111111111100000000000;
		2501: Delta = 34'sb0000100000000000000000100000000000;
		1595: Delta = 34'sb1111100000000000000000100000000000;
		4716: Delta = 34'sb0000011111111111111111100000000000;
		3810: Delta = 34'sb1111011111111111111111100000000000;
		2954: Delta = 34'sb0001000000000000000000100000000000;
		1142: Delta = 34'sb1111000000000000000000100000000000;
		5169: Delta = 34'sb0000111111111111111111100000000000;
		3357: Delta = 34'sb1110111111111111111111100000000000;
		3860: Delta = 34'sb0010000000000000000000100000000000;
		236: Delta = 34'sb1110000000000000000000100000000000;
		6075: Delta = 34'sb0001111111111111111111100000000000;
		2451: Delta = 34'sb1101111111111111111111100000000000;
		5672: Delta = 34'sb0100000000000000000000100000000000;
		4735: Delta = 34'sb1100000000000000000000100000000000;
		1576: Delta = 34'sb0011111111111111111111100000000000;
		639: Delta = 34'sb1011111111111111111111100000000000;
		5977: Delta = 34'sb0000000000000000000011000000000000;
		334: Delta = 34'sb1111111111111111111101000000000000;
		1547: Delta = 34'sb0000000000000000000101000000000000;
		4764: Delta = 34'sb1111111111111111111011000000000000;
		5309: Delta = 34'sb0000000000000000001001000000000000;
		2883: Delta = 34'sb1111111111111111111001000000000000;
		3428: Delta = 34'sb0000000000000000000111000000000000;
		1002: Delta = 34'sb1111111111111111110111000000000000;
		211: Delta = 34'sb0000000000000000010001000000000000;
		1670: Delta = 34'sb1111111111111111110001000000000000;
		4641: Delta = 34'sb0000000000000000001111000000000000;
		6100: Delta = 34'sb1111111111111111101111000000000000;
		2637: Delta = 34'sb0000000000000000100001000000000000;
		5555: Delta = 34'sb1111111111111111100001000000000000;
		756: Delta = 34'sb0000000000000000011111000000000000;
		3674: Delta = 34'sb1111111111111111011111000000000000;
		1178: Delta = 34'sb0000000000000001000001000000000000;
		703: Delta = 34'sb1111111111111111000001000000000000;
		5608: Delta = 34'sb0000000000000000111111000000000000;
		5133: Delta = 34'sb1111111111111110111111000000000000;
		4571: Delta = 34'sb0000000000000010000001000000000000;
		3621: Delta = 34'sb1111111111111110000001000000000000;
		2690: Delta = 34'sb0000000000000001111111000000000000;
		1740: Delta = 34'sb1111111111111101111111000000000000;
		5046: Delta = 34'sb0000000000000100000001000000000000;
		3146: Delta = 34'sb1111111111111100000001000000000000;
		3165: Delta = 34'sb0000000000000011111111000000000000;
		1265: Delta = 34'sb1111111111111011111111000000000000;
		5996: Delta = 34'sb0000000000001000000001000000000000;
		2196: Delta = 34'sb1111111111111000000001000000000000;
		4115: Delta = 34'sb0000000000000111111111000000000000;
		315: Delta = 34'sb1111111111110111111111000000000000;
		1585: Delta = 34'sb0000000000010000000001000000000000;
		296: Delta = 34'sb1111111111110000000001000000000000;
		6015: Delta = 34'sb0000000000001111111111000000000000;
		4726: Delta = 34'sb1111111111101111111111000000000000;
		5385: Delta = 34'sb0000000000100000000001000000000000;
		2807: Delta = 34'sb1111111111100000000001000000000000;
		3504: Delta = 34'sb0000000000011111111111000000000000;
		926: Delta = 34'sb1111111111011111111111000000000000;
		363: Delta = 34'sb0000000001000000000001000000000000;
		1518: Delta = 34'sb1111111111000000000001000000000000;
		4793: Delta = 34'sb0000000000111111111111000000000000;
		5948: Delta = 34'sb1111111110111111111111000000000000;
		2941: Delta = 34'sb0000000010000000000001000000000000;
		5251: Delta = 34'sb1111111110000000000001000000000000;
		1060: Delta = 34'sb0000000001111111111111000000000000;
		3370: Delta = 34'sb1111111101111111111111000000000000;
		1786: Delta = 34'sb0000000100000000000001000000000000;
		95: Delta = 34'sb1111111100000000000001000000000000;
		6216: Delta = 34'sb0000000011111111111111000000000000;
		4525: Delta = 34'sb1111111011111111111111000000000000;
		5787: Delta = 34'sb0000001000000000000001000000000000;
		2405: Delta = 34'sb1111111000000000000001000000000000;
		3906: Delta = 34'sb0000000111111111111111000000000000;
		524: Delta = 34'sb1111110111111111111111000000000000;
		1167: Delta = 34'sb0000010000000000000001000000000000;
		714: Delta = 34'sb1111110000000000000001000000000000;
		5597: Delta = 34'sb0000001111111111111111000000000000;
		5144: Delta = 34'sb1111101111111111111111000000000000;
		4549: Delta = 34'sb0000100000000000000001000000000000;
		3643: Delta = 34'sb1111100000000000000001000000000000;
		2668: Delta = 34'sb0000011111111111111111000000000000;
		1762: Delta = 34'sb1111011111111111111111000000000000;
		5002: Delta = 34'sb0001000000000000000001000000000000;
		3190: Delta = 34'sb1111000000000000000001000000000000;
		3121: Delta = 34'sb0000111111111111111111000000000000;
		1309: Delta = 34'sb1110111111111111111111000000000000;
		5908: Delta = 34'sb0010000000000000000001000000000000;
		2284: Delta = 34'sb1110000000000000000001000000000000;
		4027: Delta = 34'sb0001111111111111111111000000000000;
		403: Delta = 34'sb1101111111111111111111000000000000;
		1409: Delta = 34'sb0100000000000000000001000000000000;
		472: Delta = 34'sb1100000000000000000001000000000000;
		5839: Delta = 34'sb0011111111111111111111000000000000;
		4902: Delta = 34'sb1011111111111111111111000000000000;
		5643: Delta = 34'sb0000000000000000000110000000000000;
		668: Delta = 34'sb1111111111111111111010000000000000;
		3094: Delta = 34'sb0000000000000000001010000000000000;
		3217: Delta = 34'sb1111111111111111110110000000000000;
		4307: Delta = 34'sb0000000000000000010010000000000000;
		5766: Delta = 34'sb1111111111111111110010000000000000;
		545: Delta = 34'sb0000000000000000001110000000000000;
		2004: Delta = 34'sb1111111111111111101110000000000000;
		422: Delta = 34'sb0000000000000000100010000000000000;
		3340: Delta = 34'sb1111111111111111100010000000000000;
		2971: Delta = 34'sb0000000000000000011110000000000000;
		5889: Delta = 34'sb1111111111111111011110000000000000;
		5274: Delta = 34'sb0000000000000001000010000000000000;
		4799: Delta = 34'sb1111111111111111000010000000000000;
		1512: Delta = 34'sb0000000000000000111110000000000000;
		1037: Delta = 34'sb1111111111111110111110000000000000;
		2356: Delta = 34'sb0000000000000010000010000000000000;
		1406: Delta = 34'sb1111111111111110000010000000000000;
		4905: Delta = 34'sb0000000000000001111110000000000000;
		3955: Delta = 34'sb1111111111111101111110000000000000;
		2831: Delta = 34'sb0000000000000100000010000000000000;
		931: Delta = 34'sb1111111111111100000010000000000000;
		5380: Delta = 34'sb0000000000000011111110000000000000;
		3480: Delta = 34'sb1111111111111011111110000000000000;
		3781: Delta = 34'sb0000000000001000000010000000000000;
		6292: Delta = 34'sb1111111111111000000010000000000000;
		19: Delta = 34'sb0000000000000111111110000000000000;
		2530: Delta = 34'sb1111111111110111111110000000000000;
		5681: Delta = 34'sb0000000000010000000010000000000000;
		4392: Delta = 34'sb1111111111110000000010000000000000;
		1919: Delta = 34'sb0000000000001111111110000000000000;
		630: Delta = 34'sb1111111111101111111110000000000000;
		3170: Delta = 34'sb0000000000100000000010000000000000;
		592: Delta = 34'sb1111111111100000000010000000000000;
		5719: Delta = 34'sb0000000000011111111110000000000000;
		3141: Delta = 34'sb1111111111011111111110000000000000;
		4459: Delta = 34'sb0000000001000000000010000000000000;
		5614: Delta = 34'sb1111111111000000000010000000000000;
		697: Delta = 34'sb0000000000111111111110000000000000;
		1852: Delta = 34'sb1111111110111111111110000000000000;
		726: Delta = 34'sb0000000010000000000010000000000000;
		3036: Delta = 34'sb1111111110000000000010000000000000;
		3275: Delta = 34'sb0000000001111111111110000000000000;
		5585: Delta = 34'sb1111111101111111111110000000000000;
		5882: Delta = 34'sb0000000100000000000010000000000000;
		4191: Delta = 34'sb1111111100000000000010000000000000;
		2120: Delta = 34'sb0000000011111111111110000000000000;
		429: Delta = 34'sb1111111011111111111110000000000000;
		3572: Delta = 34'sb0000001000000000000010000000000000;
		190: Delta = 34'sb1111111000000000000010000000000000;
		6121: Delta = 34'sb0000000111111111111110000000000000;
		2739: Delta = 34'sb1111110111111111111110000000000000;
		5263: Delta = 34'sb0000010000000000000010000000000000;
		4810: Delta = 34'sb1111110000000000000010000000000000;
		1501: Delta = 34'sb0000001111111111111110000000000000;
		1048: Delta = 34'sb1111101111111111111110000000000000;
		2334: Delta = 34'sb0000100000000000000010000000000000;
		1428: Delta = 34'sb1111100000000000000010000000000000;
		4883: Delta = 34'sb0000011111111111111110000000000000;
		3977: Delta = 34'sb1111011111111111111110000000000000;
		2787: Delta = 34'sb0001000000000000000010000000000000;
		975: Delta = 34'sb1111000000000000000010000000000000;
		5336: Delta = 34'sb0000111111111111111110000000000000;
		3524: Delta = 34'sb1110111111111111111110000000000000;
		3693: Delta = 34'sb0010000000000000000010000000000000;
		69: Delta = 34'sb1110000000000000000010000000000000;
		6242: Delta = 34'sb0001111111111111111110000000000000;
		2618: Delta = 34'sb1101111111111111111110000000000000;
		5505: Delta = 34'sb0100000000000000000010000000000000;
		4568: Delta = 34'sb1100000000000000000010000000000000;
		1743: Delta = 34'sb0011111111111111111110000000000000;
		806: Delta = 34'sb1011111111111111111110000000000000;
		4975: Delta = 34'sb0000000000000000001100000000000000;
		1336: Delta = 34'sb1111111111111111110100000000000000;
		6188: Delta = 34'sb0000000000000000010100000000000000;
		123: Delta = 34'sb1111111111111111101100000000000000;
		2303: Delta = 34'sb0000000000000000100100000000000000;
		5221: Delta = 34'sb1111111111111111100100000000000000;
		1090: Delta = 34'sb0000000000000000011100000000000000;
		4008: Delta = 34'sb1111111111111111011100000000000000;
		844: Delta = 34'sb0000000000000001000100000000000000;
		369: Delta = 34'sb1111111111111111000100000000000000;
		5942: Delta = 34'sb0000000000000000111100000000000000;
		5467: Delta = 34'sb1111111111111110111100000000000000;
		4237: Delta = 34'sb0000000000000010000100000000000000;
		3287: Delta = 34'sb1111111111111110000100000000000000;
		3024: Delta = 34'sb0000000000000001111100000000000000;
		2074: Delta = 34'sb1111111111111101111100000000000000;
		4712: Delta = 34'sb0000000000000100000100000000000000;
		2812: Delta = 34'sb1111111111111100000100000000000000;
		3499: Delta = 34'sb0000000000000011111100000000000000;
		1599: Delta = 34'sb1111111111111011111100000000000000;
		5662: Delta = 34'sb0000000000001000000100000000000000;
		1862: Delta = 34'sb1111111111111000000100000000000000;
		4449: Delta = 34'sb0000000000000111111100000000000000;
		649: Delta = 34'sb1111111111110111111100000000000000;
		1251: Delta = 34'sb0000000000010000000100000000000000;
		6273: Delta = 34'sb1111111111110000000100000000000000;
		38: Delta = 34'sb0000000000001111111100000000000000;
		5060: Delta = 34'sb1111111111101111111100000000000000;
		5051: Delta = 34'sb0000000000100000000100000000000000;
		2473: Delta = 34'sb1111111111100000000100000000000000;
		3838: Delta = 34'sb0000000000011111111100000000000000;
		1260: Delta = 34'sb1111111111011111111100000000000000;
		29: Delta = 34'sb0000000001000000000100000000000000;
		1184: Delta = 34'sb1111111111000000000100000000000000;
		5127: Delta = 34'sb0000000000111111111100000000000000;
		6282: Delta = 34'sb1111111110111111111100000000000000;
		2607: Delta = 34'sb0000000010000000000100000000000000;
		4917: Delta = 34'sb1111111110000000000100000000000000;
		1394: Delta = 34'sb0000000001111111111100000000000000;
		3704: Delta = 34'sb1111111101111111111100000000000000;
		1452: Delta = 34'sb0000000100000000000100000000000000;
		6072: Delta = 34'sb1111111100000000000100000000000000;
		239: Delta = 34'sb0000000011111111111100000000000000;
		4859: Delta = 34'sb1111111011111111111100000000000000;
		5453: Delta = 34'sb0000001000000000000100000000000000;
		2071: Delta = 34'sb1111111000000000000100000000000000;
		4240: Delta = 34'sb0000000111111111111100000000000000;
		858: Delta = 34'sb1111110111111111111100000000000000;
		833: Delta = 34'sb0000010000000000000100000000000000;
		380: Delta = 34'sb1111110000000000000100000000000000;
		5931: Delta = 34'sb0000001111111111111100000000000000;
		5478: Delta = 34'sb1111101111111111111100000000000000;
		4215: Delta = 34'sb0000100000000000000100000000000000;
		3309: Delta = 34'sb1111100000000000000100000000000000;
		3002: Delta = 34'sb0000011111111111111100000000000000;
		2096: Delta = 34'sb1111011111111111111100000000000000;
		4668: Delta = 34'sb0001000000000000000100000000000000;
		2856: Delta = 34'sb1111000000000000000100000000000000;
		3455: Delta = 34'sb0000111111111111111100000000000000;
		1643: Delta = 34'sb1110111111111111111100000000000000;
		5574: Delta = 34'sb0010000000000000000100000000000000;
		1950: Delta = 34'sb1110000000000000000100000000000000;
		4361: Delta = 34'sb0001111111111111111100000000000000;
		737: Delta = 34'sb1101111111111111111100000000000000;
		1075: Delta = 34'sb0100000000000000000100000000000000;
		138: Delta = 34'sb1100000000000000000100000000000000;
		6173: Delta = 34'sb0011111111111111111100000000000000;
		5236: Delta = 34'sb1011111111111111111100000000000000;
		3639: Delta = 34'sb0000000000000000011000000000000000;
		2672: Delta = 34'sb1111111111111111101000000000000000;
		6065: Delta = 34'sb0000000000000000101000000000000000;
		246: Delta = 34'sb1111111111111111011000000000000000;
		4606: Delta = 34'sb0000000000000001001000000000000000;
		4131: Delta = 34'sb1111111111111111001000000000000000;
		2180: Delta = 34'sb0000000000000000111000000000000000;
		1705: Delta = 34'sb1111111111111110111000000000000000;
		1688: Delta = 34'sb0000000000000010001000000000000000;
		738: Delta = 34'sb1111111111111110001000000000000000;
		5573: Delta = 34'sb0000000000000001111000000000000000;
		4623: Delta = 34'sb1111111111111101111000000000000000;
		2163: Delta = 34'sb0000000000000100001000000000000000;
		263: Delta = 34'sb1111111111111100001000000000000000;
		6048: Delta = 34'sb0000000000000011111000000000000000;
		4148: Delta = 34'sb1111111111111011111000000000000000;
		3113: Delta = 34'sb0000000000001000001000000000000000;
		5624: Delta = 34'sb1111111111111000001000000000000000;
		687: Delta = 34'sb0000000000000111111000000000000000;
		3198: Delta = 34'sb1111111111110111111000000000000000;
		5013: Delta = 34'sb0000000000010000001000000000000000;
		3724: Delta = 34'sb1111111111110000001000000000000000;
		2587: Delta = 34'sb0000000000001111111000000000000000;
		1298: Delta = 34'sb1111111111101111111000000000000000;
		2502: Delta = 34'sb0000000000100000001000000000000000;
		6235: Delta = 34'sb1111111111100000001000000000000000;
		76: Delta = 34'sb0000000000011111111000000000000000;
		3809: Delta = 34'sb1111111111011111111000000000000000;
		3791: Delta = 34'sb0000000001000000001000000000000000;
		4946: Delta = 34'sb1111111111000000001000000000000000;
		1365: Delta = 34'sb0000000000111111111000000000000000;
		2520: Delta = 34'sb1111111110111111111000000000000000;
		58: Delta = 34'sb0000000010000000001000000000000000;
		2368: Delta = 34'sb1111111110000000001000000000000000;
		3943: Delta = 34'sb0000000001111111111000000000000000;
		6253: Delta = 34'sb1111111101111111111000000000000000;
		5214: Delta = 34'sb0000000100000000001000000000000000;
		3523: Delta = 34'sb1111111100000000001000000000000000;
		2788: Delta = 34'sb0000000011111111111000000000000000;
		1097: Delta = 34'sb1111111011111111111000000000000000;
		2904: Delta = 34'sb0000001000000000001000000000000000;
		5833: Delta = 34'sb1111111000000000001000000000000000;
		478: Delta = 34'sb0000000111111111111000000000000000;
		3407: Delta = 34'sb1111110111111111111000000000000000;
		4595: Delta = 34'sb0000010000000000001000000000000000;
		4142: Delta = 34'sb1111110000000000001000000000000000;
		2169: Delta = 34'sb0000001111111111111000000000000000;
		1716: Delta = 34'sb1111101111111111111000000000000000;
		1666: Delta = 34'sb0000100000000000001000000000000000;
		760: Delta = 34'sb1111100000000000001000000000000000;
		5551: Delta = 34'sb0000011111111111111000000000000000;
		4645: Delta = 34'sb1111011111111111111000000000000000;
		2119: Delta = 34'sb0001000000000000001000000000000000;
		307: Delta = 34'sb1111000000000000001000000000000000;
		6004: Delta = 34'sb0000111111111111111000000000000000;
		4192: Delta = 34'sb1110111111111111111000000000000000;
		3025: Delta = 34'sb0010000000000000001000000000000000;
		5712: Delta = 34'sb1110000000000000001000000000000000;
		599: Delta = 34'sb0001111111111111111000000000000000;
		3286: Delta = 34'sb1101111111111111111000000000000000;
		4837: Delta = 34'sb0100000000000000001000000000000000;
		3900: Delta = 34'sb1100000000000000001000000000000000;
		2411: Delta = 34'sb0011111111111111111000000000000000;
		1474: Delta = 34'sb1011111111111111111000000000000000;
		967: Delta = 34'sb0000000000000000110000000000000000;
		5344: Delta = 34'sb1111111111111111010000000000000000;
		5819: Delta = 34'sb0000000000000001010000000000000000;
		492: Delta = 34'sb1111111111111110110000000000000000;
		2901: Delta = 34'sb0000000000000010010000000000000000;
		1951: Delta = 34'sb1111111111111110010000000000000000;
		4360: Delta = 34'sb0000000000000001110000000000000000;
		3410: Delta = 34'sb1111111111111101110000000000000000;
		3376: Delta = 34'sb0000000000000100010000000000000000;
		1476: Delta = 34'sb1111111111111100010000000000000000;
		4835: Delta = 34'sb0000000000000011110000000000000000;
		2935: Delta = 34'sb1111111111111011110000000000000000;
		4326: Delta = 34'sb0000000000001000010000000000000000;
		526: Delta = 34'sb1111111111111000010000000000000000;
		5785: Delta = 34'sb0000000000000111110000000000000000;
		1985: Delta = 34'sb1111111111110111110000000000000000;
		6226: Delta = 34'sb0000000000010000010000000000000000;
		4937: Delta = 34'sb1111111111110000010000000000000000;
		1374: Delta = 34'sb0000000000001111110000000000000000;
		85: Delta = 34'sb1111111111101111110000000000000000;
		3715: Delta = 34'sb0000000000100000010000000000000000;
		1137: Delta = 34'sb1111111111100000010000000000000000;
		5174: Delta = 34'sb0000000000011111110000000000000000;
		2596: Delta = 34'sb1111111111011111110000000000000000;
		5004: Delta = 34'sb0000000001000000010000000000000000;
		6159: Delta = 34'sb1111111111000000010000000000000000;
		152: Delta = 34'sb0000000000111111110000000000000000;
		1307: Delta = 34'sb1111111110111111110000000000000000;
		1271: Delta = 34'sb0000000010000000010000000000000000;
		3581: Delta = 34'sb1111111110000000010000000000000000;
		2730: Delta = 34'sb0000000001111111110000000000000000;
		5040: Delta = 34'sb1111111101111111110000000000000000;
		116: Delta = 34'sb0000000100000000010000000000000000;
		4736: Delta = 34'sb1111111100000000010000000000000000;
		1575: Delta = 34'sb0000000011111111110000000000000000;
		6195: Delta = 34'sb1111111011111111110000000000000000;
		4117: Delta = 34'sb0000001000000000010000000000000000;
		735: Delta = 34'sb1111111000000000010000000000000000;
		5576: Delta = 34'sb0000000111111111110000000000000000;
		2194: Delta = 34'sb1111110111111111110000000000000000;
		5808: Delta = 34'sb0000010000000000010000000000000000;
		5355: Delta = 34'sb1111110000000000010000000000000000;
		956: Delta = 34'sb0000001111111111110000000000000000;
		503: Delta = 34'sb1111101111111111110000000000000000;
		2879: Delta = 34'sb0000100000000000010000000000000000;
		1973: Delta = 34'sb1111100000000000010000000000000000;
		4338: Delta = 34'sb0000011111111111110000000000000000;
		3432: Delta = 34'sb1111011111111111110000000000000000;
		3332: Delta = 34'sb0001000000000000010000000000000000;
		1520: Delta = 34'sb1111000000000000010000000000000000;
		4791: Delta = 34'sb0000111111111111110000000000000000;
		2979: Delta = 34'sb1110111111111111110000000000000000;
		4238: Delta = 34'sb0010000000000000010000000000000000;
		614: Delta = 34'sb1110000000000000010000000000000000;
		5697: Delta = 34'sb0001111111111111110000000000000000;
		2073: Delta = 34'sb1101111111111111110000000000000000;
		6050: Delta = 34'sb0100000000000000010000000000000000;
		5113: Delta = 34'sb1100000000000000010000000000000000;
		1198: Delta = 34'sb0011111111111111110000000000000000;
		261: Delta = 34'sb1011111111111111110000000000000000;
		1934: Delta = 34'sb0000000000000001100000000000000000;
		4377: Delta = 34'sb1111111111111110100000000000000000;
		5327: Delta = 34'sb0000000000000010100000000000000000;
		984: Delta = 34'sb1111111111111101100000000000000000;
		5802: Delta = 34'sb0000000000000100100000000000000000;
		3902: Delta = 34'sb1111111111111100100000000000000000;
		2409: Delta = 34'sb0000000000000011100000000000000000;
		509: Delta = 34'sb1111111111111011100000000000000000;
		441: Delta = 34'sb0000000000001000100000000000000000;
		2952: Delta = 34'sb1111111111111000100000000000000000;
		3359: Delta = 34'sb0000000000000111100000000000000000;
		5870: Delta = 34'sb1111111111110111100000000000000000;
		2341: Delta = 34'sb0000000000010000100000000000000000;
		1052: Delta = 34'sb1111111111110000100000000000000000;
		5259: Delta = 34'sb0000000000001111100000000000000000;
		3970: Delta = 34'sb1111111111101111100000000000000000;
		6141: Delta = 34'sb0000000000100000100000000000000000;
		3563: Delta = 34'sb1111111111100000100000000000000000;
		2748: Delta = 34'sb0000000000011111100000000000000000;
		170: Delta = 34'sb1111111111011111100000000000000000;
		1119: Delta = 34'sb0000000001000000100000000000000000;
		2274: Delta = 34'sb1111111111000000100000000000000000;
		4037: Delta = 34'sb0000000000111111100000000000000000;
		5192: Delta = 34'sb1111111110111111100000000000000000;
		3697: Delta = 34'sb0000000010000000100000000000000000;
		6007: Delta = 34'sb1111111110000000100000000000000000;
		304: Delta = 34'sb0000000001111111100000000000000000;
		2614: Delta = 34'sb1111111101111111100000000000000000;
		2542: Delta = 34'sb0000000100000000100000000000000000;
		851: Delta = 34'sb1111111100000000100000000000000000;
		5460: Delta = 34'sb0000000011111111100000000000000000;
		3769: Delta = 34'sb1111111011111111100000000000000000;
		232: Delta = 34'sb0000001000000000100000000000000000;
		3161: Delta = 34'sb1111111000000000100000000000000000;
		3150: Delta = 34'sb0000000111111111100000000000000000;
		6079: Delta = 34'sb1111110111111111100000000000000000;
		1923: Delta = 34'sb0000010000000000100000000000000000;
		1470: Delta = 34'sb1111110000000000100000000000000000;
		4841: Delta = 34'sb0000001111111111100000000000000000;
		4388: Delta = 34'sb1111101111111111100000000000000000;
		5305: Delta = 34'sb0000100000000000100000000000000000;
		4399: Delta = 34'sb1111100000000000100000000000000000;
		1912: Delta = 34'sb0000011111111111100000000000000000;
		1006: Delta = 34'sb1111011111111111100000000000000000;
		5758: Delta = 34'sb0001000000000000100000000000000000;
		3946: Delta = 34'sb1111000000000000100000000000000000;
		2365: Delta = 34'sb0000111111111111100000000000000000;
		553: Delta = 34'sb1110111111111111100000000000000000;
		353: Delta = 34'sb0010000000000000100000000000000000;
		3040: Delta = 34'sb1110000000000000100000000000000000;
		3271: Delta = 34'sb0001111111111111100000000000000000;
		5958: Delta = 34'sb1101111111111111100000000000000000;
		2165: Delta = 34'sb0100000000000000100000000000000000;
		1228: Delta = 34'sb1100000000000000100000000000000000;
		5083: Delta = 34'sb0011111111111111100000000000000000;
		4146: Delta = 34'sb1011111111111111100000000000000000;
		3868: Delta = 34'sb0000000000000011000000000000000000;
		2443: Delta = 34'sb1111111111111101000000000000000000;
		4343: Delta = 34'sb0000000000000101000000000000000000;
		1968: Delta = 34'sb1111111111111011000000000000000000;
		5293: Delta = 34'sb0000000000001001000000000000000000;
		1493: Delta = 34'sb1111111111111001000000000000000000;
		4818: Delta = 34'sb0000000000000111000000000000000000;
		1018: Delta = 34'sb1111111111110111000000000000000000;
		882: Delta = 34'sb0000000000010001000000000000000000;
		5904: Delta = 34'sb1111111111110001000000000000000000;
		407: Delta = 34'sb0000000000001111000000000000000000;
		5429: Delta = 34'sb1111111111101111000000000000000000;
		4682: Delta = 34'sb0000000000100001000000000000000000;
		2104: Delta = 34'sb1111111111100001000000000000000000;
		4207: Delta = 34'sb0000000000011111000000000000000000;
		1629: Delta = 34'sb1111111111011111000000000000000000;
		5971: Delta = 34'sb0000000001000001000000000000000000;
		815: Delta = 34'sb1111111111000001000000000000000000;
		5496: Delta = 34'sb0000000000111111000000000000000000;
		340: Delta = 34'sb1111111110111111000000000000000000;
		2238: Delta = 34'sb0000000010000001000000000000000000;
		4548: Delta = 34'sb1111111110000001000000000000000000;
		1763: Delta = 34'sb0000000001111111000000000000000000;
		4073: Delta = 34'sb1111111101111111000000000000000000;
		1083: Delta = 34'sb0000000100000001000000000000000000;
		5703: Delta = 34'sb1111111100000001000000000000000000;
		608: Delta = 34'sb0000000011111111000000000000000000;
		5228: Delta = 34'sb1111111011111111000000000000000000;
		5084: Delta = 34'sb0000001000000001000000000000000000;
		1702: Delta = 34'sb1111111000000001000000000000000000;
		4609: Delta = 34'sb0000000111111111000000000000000000;
		1227: Delta = 34'sb1111110111111111000000000000000000;
		464: Delta = 34'sb0000010000000001000000000000000000;
		11: Delta = 34'sb1111110000000001000000000000000000;
		6300: Delta = 34'sb0000001111111111000000000000000000;
		5847: Delta = 34'sb1111101111111111000000000000000000;
		3846: Delta = 34'sb0000100000000001000000000000000000;
		2940: Delta = 34'sb1111100000000001000000000000000000;
		3371: Delta = 34'sb0000011111111111000000000000000000;
		2465: Delta = 34'sb1111011111111111000000000000000000;
		4299: Delta = 34'sb0001000000000001000000000000000000;
		2487: Delta = 34'sb1111000000000001000000000000000000;
		3824: Delta = 34'sb0000111111111111000000000000000000;
		2012: Delta = 34'sb1110111111111111000000000000000000;
		5205: Delta = 34'sb0010000000000001000000000000000000;
		1581: Delta = 34'sb1110000000000001000000000000000000;
		4730: Delta = 34'sb0001111111111111000000000000000000;
		1106: Delta = 34'sb1101111111111111000000000000000000;
		706: Delta = 34'sb0100000000000001000000000000000000;
		6080: Delta = 34'sb1100000000000001000000000000000000;
		231: Delta = 34'sb0011111111111111000000000000000000;
		5605: Delta = 34'sb1011111111111111000000000000000000;
		1425: Delta = 34'sb0000000000000110000000000000000000;
		4886: Delta = 34'sb1111111111111010000000000000000000;
		2375: Delta = 34'sb0000000000001010000000000000000000;
		3936: Delta = 34'sb1111111111110110000000000000000000;
		4275: Delta = 34'sb0000000000010010000000000000000000;
		2986: Delta = 34'sb1111111111110010000000000000000000;
		3325: Delta = 34'sb0000000000001110000000000000000000;
		2036: Delta = 34'sb1111111111101110000000000000000000;
		1764: Delta = 34'sb0000000000100010000000000000000000;
		5497: Delta = 34'sb1111111111100010000000000000000000;
		814: Delta = 34'sb0000000000011110000000000000000000;
		4547: Delta = 34'sb1111111111011110000000000000000000;
		3053: Delta = 34'sb0000000001000010000000000000000000;
		4208: Delta = 34'sb1111111111000010000000000000000000;
		2103: Delta = 34'sb0000000000111110000000000000000000;
		3258: Delta = 34'sb1111111110111110000000000000000000;
		5631: Delta = 34'sb0000000010000010000000000000000000;
		1630: Delta = 34'sb1111111110000010000000000000000000;
		4681: Delta = 34'sb0000000001111110000000000000000000;
		680: Delta = 34'sb1111111101111110000000000000000000;
		4476: Delta = 34'sb0000000100000010000000000000000000;
		2785: Delta = 34'sb1111111100000010000000000000000000;
		3526: Delta = 34'sb0000000011111110000000000000000000;
		1835: Delta = 34'sb1111111011111110000000000000000000;
		2166: Delta = 34'sb0000001000000010000000000000000000;
		5095: Delta = 34'sb1111111000000010000000000000000000;
		1216: Delta = 34'sb0000000111111110000000000000000000;
		4145: Delta = 34'sb1111110111111110000000000000000000;
		3857: Delta = 34'sb0000010000000010000000000000000000;
		3404: Delta = 34'sb1111110000000010000000000000000000;
		2907: Delta = 34'sb0000001111111110000000000000000000;
		2454: Delta = 34'sb1111101111111110000000000000000000;
		928: Delta = 34'sb0000100000000010000000000000000000;
		22: Delta = 34'sb1111100000000010000000000000000000;
		6289: Delta = 34'sb0000011111111110000000000000000000;
		5383: Delta = 34'sb1111011111111110000000000000000000;
		1381: Delta = 34'sb0001000000000010000000000000000000;
		5880: Delta = 34'sb1111000000000010000000000000000000;
		431: Delta = 34'sb0000111111111110000000000000000000;
		4930: Delta = 34'sb1110111111111110000000000000000000;
		2287: Delta = 34'sb0010000000000010000000000000000000;
		4974: Delta = 34'sb1110000000000010000000000000000000;
		1337: Delta = 34'sb0001111111111110000000000000000000;
		4024: Delta = 34'sb1101111111111110000000000000000000;
		4099: Delta = 34'sb0100000000000010000000000000000000;
		3162: Delta = 34'sb1100000000000010000000000000000000;
		3149: Delta = 34'sb0011111111111110000000000000000000;
		2212: Delta = 34'sb1011111111111110000000000000000000;
		2850: Delta = 34'sb0000000000001100000000000000000000;
		3461: Delta = 34'sb1111111111110100000000000000000000;
		4750: Delta = 34'sb0000000000010100000000000000000000;
		1561: Delta = 34'sb1111111111101100000000000000000000;
		2239: Delta = 34'sb0000000000100100000000000000000000;
		5972: Delta = 34'sb1111111111100100000000000000000000;
		339: Delta = 34'sb0000000000011100000000000000000000;
		4072: Delta = 34'sb1111111111011100000000000000000000;
		3528: Delta = 34'sb0000000001000100000000000000000000;
		4683: Delta = 34'sb1111111111000100000000000000000000;
		1628: Delta = 34'sb0000000000111100000000000000000000;
		2783: Delta = 34'sb1111111110111100000000000000000000;
		6106: Delta = 34'sb0000000010000100000000000000000000;
		2105: Delta = 34'sb1111111110000100000000000000000000;
		4206: Delta = 34'sb0000000001111100000000000000000000;
		205: Delta = 34'sb1111111101111100000000000000000000;
		4951: Delta = 34'sb0000000100000100000000000000000000;
		3260: Delta = 34'sb1111111100000100000000000000000000;
		3051: Delta = 34'sb0000000011111100000000000000000000;
		1360: Delta = 34'sb1111111011111100000000000000000000;
		2641: Delta = 34'sb0000001000000100000000000000000000;
		5570: Delta = 34'sb1111111000000100000000000000000000;
		741: Delta = 34'sb0000000111111100000000000000000000;
		3670: Delta = 34'sb1111110111111100000000000000000000;
		4332: Delta = 34'sb0000010000000100000000000000000000;
		3879: Delta = 34'sb1111110000000100000000000000000000;
		2432: Delta = 34'sb0000001111111100000000000000000000;
		1979: Delta = 34'sb1111101111111100000000000000000000;
		1403: Delta = 34'sb0000100000000100000000000000000000;
		497: Delta = 34'sb1111100000000100000000000000000000;
		5814: Delta = 34'sb0000011111111100000000000000000000;
		4908: Delta = 34'sb1111011111111100000000000000000000;
		1856: Delta = 34'sb0001000000000100000000000000000000;
		44: Delta = 34'sb1111000000000100000000000000000000;
		6267: Delta = 34'sb0000111111111100000000000000000000;
		4455: Delta = 34'sb1110111111111100000000000000000000;
		2762: Delta = 34'sb0010000000000100000000000000000000;
		5449: Delta = 34'sb1110000000000100000000000000000000;
		862: Delta = 34'sb0001111111111100000000000000000000;
		3549: Delta = 34'sb1101111111111100000000000000000000;
		4574: Delta = 34'sb0100000000000100000000000000000000;
		3637: Delta = 34'sb1100000000000100000000000000000000;
		2674: Delta = 34'sb0011111111111100000000000000000000;
		1737: Delta = 34'sb1011111111111100000000000000000000;
		5700: Delta = 34'sb0000000000011000000000000000000000;
		611: Delta = 34'sb1111111111101000000000000000000000;
		3189: Delta = 34'sb0000000000101000000000000000000000;
		3122: Delta = 34'sb1111111111011000000000000000000000;
		4478: Delta = 34'sb0000000001001000000000000000000000;
		5633: Delta = 34'sb1111111111001000000000000000000000;
		678: Delta = 34'sb0000000000111000000000000000000000;
		1833: Delta = 34'sb1111111110111000000000000000000000;
		745: Delta = 34'sb0000000010001000000000000000000000;
		3055: Delta = 34'sb1111111110001000000000000000000000;
		3256: Delta = 34'sb0000000001111000000000000000000000;
		5566: Delta = 34'sb1111111101111000000000000000000000;
		5901: Delta = 34'sb0000000100001000000000000000000000;
		4210: Delta = 34'sb1111111100001000000000000000000000;
		2101: Delta = 34'sb0000000011111000000000000000000000;
		410: Delta = 34'sb1111111011111000000000000000000000;
		3591: Delta = 34'sb0000001000001000000000000000000000;
		209: Delta = 34'sb1111111000001000000000000000000000;
		6102: Delta = 34'sb0000000111111000000000000000000000;
		2720: Delta = 34'sb1111110111111000000000000000000000;
		5282: Delta = 34'sb0000010000001000000000000000000000;
		4829: Delta = 34'sb1111110000001000000000000000000000;
		1482: Delta = 34'sb0000001111111000000000000000000000;
		1029: Delta = 34'sb1111101111111000000000000000000000;
		2353: Delta = 34'sb0000100000001000000000000000000000;
		1447: Delta = 34'sb1111100000001000000000000000000000;
		4864: Delta = 34'sb0000011111111000000000000000000000;
		3958: Delta = 34'sb1111011111111000000000000000000000;
		2806: Delta = 34'sb0001000000001000000000000000000000;
		994: Delta = 34'sb1111000000001000000000000000000000;
		5317: Delta = 34'sb0000111111111000000000000000000000;
		3505: Delta = 34'sb1110111111111000000000000000000000;
		3712: Delta = 34'sb0010000000001000000000000000000000;
		88: Delta = 34'sb1110000000001000000000000000000000;
		6223: Delta = 34'sb0001111111111000000000000000000000;
		2599: Delta = 34'sb1101111111111000000000000000000000;
		5524: Delta = 34'sb0100000000001000000000000000000000;
		4587: Delta = 34'sb1100000000001000000000000000000000;
		1724: Delta = 34'sb0011111111111000000000000000000000;
		787: Delta = 34'sb1011111111111000000000000000000000;
		5089: Delta = 34'sb0000000000110000000000000000000000;
		1222: Delta = 34'sb1111111111010000000000000000000000;
		67: Delta = 34'sb0000000001010000000000000000000000;
		6244: Delta = 34'sb1111111110110000000000000000000000;
		2645: Delta = 34'sb0000000010010000000000000000000000;
		4955: Delta = 34'sb1111111110010000000000000000000000;
		1356: Delta = 34'sb0000000001110000000000000000000000;
		3666: Delta = 34'sb1111111101110000000000000000000000;
		1490: Delta = 34'sb0000000100010000000000000000000000;
		6110: Delta = 34'sb1111111100010000000000000000000000;
		201: Delta = 34'sb0000000011110000000000000000000000;
		4821: Delta = 34'sb1111111011110000000000000000000000;
		5491: Delta = 34'sb0000001000010000000000000000000000;
		2109: Delta = 34'sb1111111000010000000000000000000000;
		4202: Delta = 34'sb0000000111110000000000000000000000;
		820: Delta = 34'sb1111110111110000000000000000000000;
		871: Delta = 34'sb0000010000010000000000000000000000;
		418: Delta = 34'sb1111110000010000000000000000000000;
		5893: Delta = 34'sb0000001111110000000000000000000000;
		5440: Delta = 34'sb1111101111110000000000000000000000;
		4253: Delta = 34'sb0000100000010000000000000000000000;
		3347: Delta = 34'sb1111100000010000000000000000000000;
		2964: Delta = 34'sb0000011111110000000000000000000000;
		2058: Delta = 34'sb1111011111110000000000000000000000;
		4706: Delta = 34'sb0001000000010000000000000000000000;
		2894: Delta = 34'sb1111000000010000000000000000000000;
		3417: Delta = 34'sb0000111111110000000000000000000000;
		1605: Delta = 34'sb1110111111110000000000000000000000;
		5612: Delta = 34'sb0010000000010000000000000000000000;
		1988: Delta = 34'sb1110000000010000000000000000000000;
		4323: Delta = 34'sb0001111111110000000000000000000000;
		699: Delta = 34'sb1101111111110000000000000000000000;
		1113: Delta = 34'sb0100000000010000000000000000000000;
		176: Delta = 34'sb1100000000010000000000000000000000;
		6135: Delta = 34'sb0011111111110000000000000000000000;
		5198: Delta = 34'sb1011111111110000000000000000000000;
		3867: Delta = 34'sb0000000001100000000000000000000000;
		2444: Delta = 34'sb1111111110100000000000000000000000;
		134: Delta = 34'sb0000000010100000000000000000000000;
		6177: Delta = 34'sb1111111101100000000000000000000000;
		5290: Delta = 34'sb0000000100100000000000000000000000;
		3599: Delta = 34'sb1111111100100000000000000000000000;
		2712: Delta = 34'sb0000000011100000000000000000000000;
		1021: Delta = 34'sb1111111011100000000000000000000000;
		2980: Delta = 34'sb0000001000100000000000000000000000;
		5909: Delta = 34'sb1111111000100000000000000000000000;
		402: Delta = 34'sb0000000111100000000000000000000000;
		3331: Delta = 34'sb1111110111100000000000000000000000;
		4671: Delta = 34'sb0000010000100000000000000000000000;
		4218: Delta = 34'sb1111110000100000000000000000000000;
		2093: Delta = 34'sb0000001111100000000000000000000000;
		1640: Delta = 34'sb1111101111100000000000000000000000;
		1742: Delta = 34'sb0000100000100000000000000000000000;
		836: Delta = 34'sb1111100000100000000000000000000000;
		5475: Delta = 34'sb0000011111100000000000000000000000;
		4569: Delta = 34'sb1111011111100000000000000000000000;
		2195: Delta = 34'sb0001000000100000000000000000000000;
		383: Delta = 34'sb1111000000100000000000000000000000;
		5928: Delta = 34'sb0000111111100000000000000000000000;
		4116: Delta = 34'sb1110111111100000000000000000000000;
		3101: Delta = 34'sb0010000000100000000000000000000000;
		5788: Delta = 34'sb1110000000100000000000000000000000;
		523: Delta = 34'sb0001111111100000000000000000000000;
		3210: Delta = 34'sb1101111111100000000000000000000000;
		4913: Delta = 34'sb0100000000100000000000000000000000;
		3976: Delta = 34'sb1100000000100000000000000000000000;
		2335: Delta = 34'sb0011111111100000000000000000000000;
		1398: Delta = 34'sb1011111111100000000000000000000000;
		1423: Delta = 34'sb0000000011000000000000000000000000;
		4888: Delta = 34'sb1111111101000000000000000000000000;
		268: Delta = 34'sb0000000101000000000000000000000000;
		6043: Delta = 34'sb1111111011000000000000000000000000;
		4269: Delta = 34'sb0000001001000000000000000000000000;
		887: Delta = 34'sb1111111001000000000000000000000000;
		5424: Delta = 34'sb0000000111000000000000000000000000;
		2042: Delta = 34'sb1111110111000000000000000000000000;
		5960: Delta = 34'sb0000010001000000000000000000000000;
		5507: Delta = 34'sb1111110001000000000000000000000000;
		804: Delta = 34'sb0000001111000000000000000000000000;
		351: Delta = 34'sb1111101111000000000000000000000000;
		3031: Delta = 34'sb0000100001000000000000000000000000;
		2125: Delta = 34'sb1111100001000000000000000000000000;
		4186: Delta = 34'sb0000011111000000000000000000000000;
		3280: Delta = 34'sb1111011111000000000000000000000000;
		3484: Delta = 34'sb0001000001000000000000000000000000;
		1672: Delta = 34'sb1111000001000000000000000000000000;
		4639: Delta = 34'sb0000111111000000000000000000000000;
		2827: Delta = 34'sb1110111111000000000000000000000000;
		4390: Delta = 34'sb0010000001000000000000000000000000;
		766: Delta = 34'sb1110000001000000000000000000000000;
		5545: Delta = 34'sb0001111111000000000000000000000000;
		1921: Delta = 34'sb1101111111000000000000000000000000;
		6202: Delta = 34'sb0100000001000000000000000000000000;
		5265: Delta = 34'sb1100000001000000000000000000000000;
		1046: Delta = 34'sb0011111111000000000000000000000000;
		109: Delta = 34'sb1011111111000000000000000000000000;
		2846: Delta = 34'sb0000000110000000000000000000000000;
		3465: Delta = 34'sb1111111010000000000000000000000000;
		536: Delta = 34'sb0000001010000000000000000000000000;
		5775: Delta = 34'sb1111110110000000000000000000000000;
		2227: Delta = 34'sb0000010010000000000000000000000000;
		1774: Delta = 34'sb1111110010000000000000000000000000;
		4537: Delta = 34'sb0000001110000000000000000000000000;
		4084: Delta = 34'sb1111101110000000000000000000000000;
		5609: Delta = 34'sb0000100010000000000000000000000000;
		4703: Delta = 34'sb1111100010000000000000000000000000;
		1608: Delta = 34'sb0000011110000000000000000000000000;
		702: Delta = 34'sb1111011110000000000000000000000000;
		6062: Delta = 34'sb0001000010000000000000000000000000;
		4250: Delta = 34'sb1111000010000000000000000000000000;
		2061: Delta = 34'sb0000111110000000000000000000000000;
		249: Delta = 34'sb1110111110000000000000000000000000;
		657: Delta = 34'sb0010000010000000000000000000000000;
		3344: Delta = 34'sb1110000010000000000000000000000000;
		2967: Delta = 34'sb0001111110000000000000000000000000;
		5654: Delta = 34'sb1101111110000000000000000000000000;
		2469: Delta = 34'sb0100000010000000000000000000000000;
		1532: Delta = 34'sb1100000010000000000000000000000000;
		4779: Delta = 34'sb0011111110000000000000000000000000;
		3842: Delta = 34'sb1011111110000000000000000000000000;
		5692: Delta = 34'sb0000001100000000000000000000000000;
		619: Delta = 34'sb1111110100000000000000000000000000;
		1072: Delta = 34'sb0000010100000000000000000000000000;
		5239: Delta = 34'sb1111101100000000000000000000000000;
		4454: Delta = 34'sb0000100100000000000000000000000000;
		3548: Delta = 34'sb1111100100000000000000000000000000;
		2763: Delta = 34'sb0000011100000000000000000000000000;
		1857: Delta = 34'sb1111011100000000000000000000000000;
		4907: Delta = 34'sb0001000100000000000000000000000000;
		3095: Delta = 34'sb1111000100000000000000000000000000;
		3216: Delta = 34'sb0000111100000000000000000000000000;
		1404: Delta = 34'sb1110111100000000000000000000000000;
		5813: Delta = 34'sb0010000100000000000000000000000000;
		2189: Delta = 34'sb1110000100000000000000000000000000;
		4122: Delta = 34'sb0001111100000000000000000000000000;
		498: Delta = 34'sb1101111100000000000000000000000000;
		1314: Delta = 34'sb0100000100000000000000000000000000;
		377: Delta = 34'sb1100000100000000000000000000000000;
		5934: Delta = 34'sb0011111100000000000000000000000000;
		4997: Delta = 34'sb1011111100000000000000000000000000;
		5073: Delta = 34'sb0000011000000000000000000000000000;
		1238: Delta = 34'sb1111101000000000000000000000000000;
		2144: Delta = 34'sb0000101000000000000000000000000000;
		4167: Delta = 34'sb1111011000000000000000000000000000;
		2597: Delta = 34'sb0001001000000000000000000000000000;
		785: Delta = 34'sb1111001000000000000000000000000000;
		5526: Delta = 34'sb0000111000000000000000000000000000;
		3714: Delta = 34'sb1110111000000000000000000000000000;
		3503: Delta = 34'sb0010001000000000000000000000000000;
		6190: Delta = 34'sb1110001000000000000000000000000000;
		121: Delta = 34'sb0001111000000000000000000000000000;
		2808: Delta = 34'sb1101111000000000000000000000000000;
		5315: Delta = 34'sb0100001000000000000000000000000000;
		4378: Delta = 34'sb1100001000000000000000000000000000;
		1933: Delta = 34'sb0011111000000000000000000000000000;
		996: Delta = 34'sb1011111000000000000000000000000000;
		3835: Delta = 34'sb0000110000000000000000000000000000;
		2476: Delta = 34'sb1111010000000000000000000000000000;
		4288: Delta = 34'sb0001010000000000000000000000000000;
		2023: Delta = 34'sb1110110000000000000000000000000000;
		5194: Delta = 34'sb0010010000000000000000000000000000;
		1570: Delta = 34'sb1110010000000000000000000000000000;
		4741: Delta = 34'sb0001110000000000000000000000000000;
		1117: Delta = 34'sb1101110000000000000000000000000000;
		695: Delta = 34'sb0100010000000000000000000000000000;
		6069: Delta = 34'sb1100010000000000000000000000000000;
		242: Delta = 34'sb0011110000000000000000000000000000;
		5616: Delta = 34'sb1011110000000000000000000000000000;
		1359: Delta = 34'sb0001100000000000000000000000000000;
		4952: Delta = 34'sb1110100000000000000000000000000000;
		2265: Delta = 34'sb0010100000000000000000000000000000;
		4046: Delta = 34'sb1101100000000000000000000000000000;
		4077: Delta = 34'sb0100100000000000000000000000000000;
		3140: Delta = 34'sb1100100000000000000000000000000000;
		3171: Delta = 34'sb0011100000000000000000000000000000;
		2234: Delta = 34'sb1011100000000000000000000000000000;
		2718: Delta = 34'sb0011000000000000000000000000000000;
		3593: Delta = 34'sb1101000000000000000000000000000000;
		4530: Delta = 34'sb0101000000000000000000000000000000;
		1781: Delta = 34'sb1011000000000000000000000000000000;
		5436: Delta = 34'sb0110000000000000000000000000000000;
		875: Delta = 34'sb1010000000000000000000000000000000;
		default: Delta =34'sb0;
	endcase
end

wire signed [W_BITS-1:0] W_signed;
assign W_signed = (W - Delta);

always@(posedge clk or negedge rst_n) begin
   if(!rst_n) begin
     	ps <= idle;
    end
   else begin
        case(ps)
            idle: begin
                found <= 0;
                R <= 0;
        	Q <= 0;
                ps <= pre;
                end
	    pre: begin
		 Q <= W / A;
		 ps <= load;
		end
            load: begin
                 R <= W - (A * Q);
		 ps <= LUT;
		end
	    LUT: begin
		  if(Delta != 0)begin
		      N <= W_signed / A ;	
		      found <= 1;
                      ps <= idle;
		  end
		  else begin
		      N <= Q;
		      found <= 1;
                      ps <= idle;
		  end
		end
	endcase
    end
end

endmodule


// Product (AN) Code DEC r-LUT
// DEC_rLUT4bits.v
// Used to do DEC, but corrected errors by locations, not AWE
// Received remainder r, output two error locations.
module DEC_rLUT4bits(r, l_1, l_2);
input 	[9:0]	r;
output	reg	signed	[4:0]	l_1;
output	reg	signed	[4:0]	l_2;
always@(*) begin
	case(r)
		1: begin l_1 = -1;
				 l_2 = +2; end
		654: begin l_1 = +1;
				 l_2 = -2; end
		2: begin l_1 = +1;
				 l_2 = +1; end
		653: begin l_1 = -1;
				 l_2 = -1; end
		4: begin l_1 = +2;
				 l_2 = +2; end
		651: begin l_1 = -2;
				 l_2 = -2; end
		8: begin l_1 = +3;
				 l_2 = +3; end
		647: begin l_1 = -3;
				 l_2 = -3; end
		16: begin l_1 = +4;
				 l_2 = +4; end
		639: begin l_1 = -4;
				 l_2 = -4; end
		32: begin l_1 = +5;
				 l_2 = +5; end
		623: begin l_1 = -5;
				 l_2 = -5; end
		64: begin l_1 = +6;
				 l_2 = +6; end
		591: begin l_1 = -6;
				 l_2 = -6; end
		128: begin l_1 = +7;
				 l_2 = +7; end
		527: begin l_1 = -7;
				 l_2 = -7; end
		256: begin l_1 = +8;
				 l_2 = +8; end
		399: begin l_1 = -8;
				 l_2 = -8; end
		512: begin l_1 = +9;
				 l_2 = +9; end
		143: begin l_1 = -9;
				 l_2 = -9; end
		369: begin l_1 = +10;
				 l_2 = +10; end
		286: begin l_1 = -10;
				 l_2 = -10; end
		83: begin l_1 = +11;
				 l_2 = +11; end
		572: begin l_1 = -11;
				 l_2 = -11; end
		166: begin l_1 = +12;
				 l_2 = +12; end
		489: begin l_1 = -12;
				 l_2 = -12; end
		332: begin l_1 = +13;
				 l_2 = +13; end
		323: begin l_1 = -13;
				 l_2 = -13; end
		3: begin l_1 = -1;
				 l_2 = +3; end
		652: begin l_1 = -1;
				 l_2 = -2; end
		5: begin l_1 = +1;
				 l_2 = +3; end
		650: begin l_1 = -1;
				 l_2 = -3; end
		9: begin l_1 = +1;
				 l_2 = +4; end
		648: begin l_1 = +1;
				 l_2 = -4; end
		7: begin l_1 = -1;
				 l_2 = +4; end
		646: begin l_1 = -1;
				 l_2 = -4; end
		17: begin l_1 = +1;
				 l_2 = +5; end
		640: begin l_1 = +1;
				 l_2 = -5; end
		15: begin l_1 = -1;
				 l_2 = +5; end
		638: begin l_1 = -1;
				 l_2 = -5; end
		33: begin l_1 = +1;
				 l_2 = +6; end
		624: begin l_1 = +1;
				 l_2 = -6; end
		31: begin l_1 = -1;
				 l_2 = +6; end
		622: begin l_1 = -1;
				 l_2 = -6; end
		65: begin l_1 = +1;
				 l_2 = +7; end
		592: begin l_1 = +1;
				 l_2 = -7; end
		63: begin l_1 = -1;
				 l_2 = +7; end
		590: begin l_1 = -1;
				 l_2 = -7; end
		129: begin l_1 = +1;
				 l_2 = +8; end
		528: begin l_1 = +1;
				 l_2 = -8; end
		127: begin l_1 = -1;
				 l_2 = +8; end
		526: begin l_1 = -1;
				 l_2 = -8; end
		257: begin l_1 = +1;
				 l_2 = +9; end
		400: begin l_1 = +1;
				 l_2 = -9; end
		255: begin l_1 = -1;
				 l_2 = +9; end
		398: begin l_1 = -1;
				 l_2 = -9; end
		513: begin l_1 = +1;
				 l_2 = +10; end
		144: begin l_1 = +1;
				 l_2 = -10; end
		511: begin l_1 = -1;
				 l_2 = +10; end
		142: begin l_1 = -1;
				 l_2 = -10; end
		370: begin l_1 = +1;
				 l_2 = +11; end
		287: begin l_1 = +1;
				 l_2 = -11; end
		368: begin l_1 = -1;
				 l_2 = +11; end
		285: begin l_1 = -1;
				 l_2 = -11; end
		84: begin l_1 = +1;
				 l_2 = +12; end
		573: begin l_1 = +1;
				 l_2 = -12; end
		82: begin l_1 = -1;
				 l_2 = +12; end
		571: begin l_1 = -1;
				 l_2 = -12; end
		167: begin l_1 = +1;
				 l_2 = +13; end
		490: begin l_1 = +1;
				 l_2 = -13; end
		165: begin l_1 = -1;
				 l_2 = +13; end
		488: begin l_1 = -1;
				 l_2 = -13; end
		333: begin l_1 = +1;
				 l_2 = +14; end
		324: begin l_1 = +1;
				 l_2 = -14; end
		331: begin l_1 = -1;
				 l_2 = +14; end
		322: begin l_1 = -1;
				 l_2 = -14; end
		6: begin l_1 = -2;
				 l_2 = +4; end
		649: begin l_1 = -2;
				 l_2 = -3; end
		10: begin l_1 = +2;
				 l_2 = +4; end
		645: begin l_1 = -2;
				 l_2 = -4; end
		18: begin l_1 = +2;
				 l_2 = +5; end
		641: begin l_1 = +2;
				 l_2 = -5; end
		14: begin l_1 = -2;
				 l_2 = +5; end
		637: begin l_1 = -2;
				 l_2 = -5; end
		34: begin l_1 = +2;
				 l_2 = +6; end
		625: begin l_1 = +2;
				 l_2 = -6; end
		30: begin l_1 = -2;
				 l_2 = +6; end
		621: begin l_1 = -2;
				 l_2 = -6; end
		66: begin l_1 = +2;
				 l_2 = +7; end
		593: begin l_1 = +2;
				 l_2 = -7; end
		62: begin l_1 = -2;
				 l_2 = +7; end
		589: begin l_1 = -2;
				 l_2 = -7; end
		130: begin l_1 = +2;
				 l_2 = +8; end
		529: begin l_1 = +2;
				 l_2 = -8; end
		126: begin l_1 = -2;
				 l_2 = +8; end
		525: begin l_1 = -2;
				 l_2 = -8; end
		258: begin l_1 = +2;
				 l_2 = +9; end
		401: begin l_1 = +2;
				 l_2 = -9; end
		254: begin l_1 = -2;
				 l_2 = +9; end
		397: begin l_1 = -2;
				 l_2 = -9; end
		514: begin l_1 = +2;
				 l_2 = +10; end
		145: begin l_1 = +2;
				 l_2 = -10; end
		510: begin l_1 = -2;
				 l_2 = +10; end
		141: begin l_1 = -2;
				 l_2 = -10; end
		371: begin l_1 = +2;
				 l_2 = +11; end
		288: begin l_1 = +2;
				 l_2 = -11; end
		367: begin l_1 = -2;
				 l_2 = +11; end
		284: begin l_1 = -2;
				 l_2 = -11; end
		85: begin l_1 = +2;
				 l_2 = +12; end
		574: begin l_1 = +2;
				 l_2 = -12; end
		81: begin l_1 = -2;
				 l_2 = +12; end
		570: begin l_1 = -2;
				 l_2 = -12; end
		168: begin l_1 = +2;
				 l_2 = +13; end
		491: begin l_1 = +2;
				 l_2 = -13; end
		164: begin l_1 = -2;
				 l_2 = +13; end
		487: begin l_1 = -2;
				 l_2 = -13; end
		334: begin l_1 = +2;
				 l_2 = +14; end
		325: begin l_1 = +2;
				 l_2 = -14; end
		330: begin l_1 = -2;
				 l_2 = +14; end
		321: begin l_1 = -2;
				 l_2 = -14; end
		12: begin l_1 = -3;
				 l_2 = +5; end
		643: begin l_1 = -3;
				 l_2 = -4; end
		20: begin l_1 = +3;
				 l_2 = +5; end
		635: begin l_1 = -3;
				 l_2 = -5; end
		36: begin l_1 = +3;
				 l_2 = +6; end
		627: begin l_1 = +3;
				 l_2 = -6; end
		28: begin l_1 = -3;
				 l_2 = +6; end
		619: begin l_1 = -3;
				 l_2 = -6; end
		68: begin l_1 = +3;
				 l_2 = +7; end
		595: begin l_1 = +3;
				 l_2 = -7; end
		60: begin l_1 = -3;
				 l_2 = +7; end
		587: begin l_1 = -3;
				 l_2 = -7; end
		132: begin l_1 = +3;
				 l_2 = +8; end
		531: begin l_1 = +3;
				 l_2 = -8; end
		124: begin l_1 = -3;
				 l_2 = +8; end
		523: begin l_1 = -3;
				 l_2 = -8; end
		260: begin l_1 = +3;
				 l_2 = +9; end
		403: begin l_1 = +3;
				 l_2 = -9; end
		252: begin l_1 = -3;
				 l_2 = +9; end
		395: begin l_1 = -3;
				 l_2 = -9; end
		516: begin l_1 = +3;
				 l_2 = +10; end
		147: begin l_1 = +3;
				 l_2 = -10; end
		508: begin l_1 = -3;
				 l_2 = +10; end
		139: begin l_1 = -3;
				 l_2 = -10; end
		373: begin l_1 = +3;
				 l_2 = +11; end
		290: begin l_1 = +3;
				 l_2 = -11; end
		365: begin l_1 = -3;
				 l_2 = +11; end
		282: begin l_1 = -3;
				 l_2 = -11; end
		87: begin l_1 = +3;
				 l_2 = +12; end
		576: begin l_1 = +3;
				 l_2 = -12; end
		79: begin l_1 = -3;
				 l_2 = +12; end
		568: begin l_1 = -3;
				 l_2 = -12; end
		170: begin l_1 = +3;
				 l_2 = +13; end
		493: begin l_1 = +3;
				 l_2 = -13; end
		162: begin l_1 = -3;
				 l_2 = +13; end
		485: begin l_1 = -3;
				 l_2 = -13; end
		336: begin l_1 = +3;
				 l_2 = +14; end
		327: begin l_1 = +3;
				 l_2 = -14; end
		328: begin l_1 = -3;
				 l_2 = +14; end
		319: begin l_1 = -3;
				 l_2 = -14; end
		24: begin l_1 = -4;
				 l_2 = +6; end
		631: begin l_1 = -4;
				 l_2 = -5; end
		40: begin l_1 = +4;
				 l_2 = +6; end
		615: begin l_1 = -4;
				 l_2 = -6; end
		72: begin l_1 = +4;
				 l_2 = +7; end
		599: begin l_1 = +4;
				 l_2 = -7; end
		56: begin l_1 = -4;
				 l_2 = +7; end
		583: begin l_1 = -4;
				 l_2 = -7; end
		136: begin l_1 = +4;
				 l_2 = +8; end
		535: begin l_1 = +4;
				 l_2 = -8; end
		120: begin l_1 = -4;
				 l_2 = +8; end
		519: begin l_1 = -4;
				 l_2 = -8; end
		264: begin l_1 = +4;
				 l_2 = +9; end
		407: begin l_1 = +4;
				 l_2 = -9; end
		248: begin l_1 = -4;
				 l_2 = +9; end
		391: begin l_1 = -4;
				 l_2 = -9; end
		520: begin l_1 = +4;
				 l_2 = +10; end
		151: begin l_1 = +4;
				 l_2 = -10; end
		504: begin l_1 = -4;
				 l_2 = +10; end
		135: begin l_1 = -4;
				 l_2 = -10; end
		377: begin l_1 = +4;
				 l_2 = +11; end
		294: begin l_1 = +4;
				 l_2 = -11; end
		361: begin l_1 = -4;
				 l_2 = +11; end
		278: begin l_1 = -4;
				 l_2 = -11; end
		91: begin l_1 = +4;
				 l_2 = +12; end
		580: begin l_1 = +4;
				 l_2 = -12; end
		75: begin l_1 = -4;
				 l_2 = +12; end
		564: begin l_1 = -4;
				 l_2 = -12; end
		174: begin l_1 = +4;
				 l_2 = +13; end
		497: begin l_1 = +4;
				 l_2 = -13; end
		158: begin l_1 = -4;
				 l_2 = +13; end
		481: begin l_1 = -4;
				 l_2 = -13; end
		340: begin l_1 = +4;
				 l_2 = +14; end
		331: begin l_1 = -1;
				 l_2 = +14; end
		324: begin l_1 = +1;
				 l_2 = -14; end
		315: begin l_1 = -4;
				 l_2 = -14; end
		48: begin l_1 = -5;
				 l_2 = +7; end
		607: begin l_1 = -5;
				 l_2 = -6; end
		80: begin l_1 = +5;
				 l_2 = +7; end
		575: begin l_1 = -5;
				 l_2 = -7; end
		144: begin l_1 = +1;
				 l_2 = -10; end
		543: begin l_1 = +5;
				 l_2 = -8; end
		112: begin l_1 = -5;
				 l_2 = +8; end
		511: begin l_1 = -1;
				 l_2 = +10; end
		272: begin l_1 = +5;
				 l_2 = +9; end
		415: begin l_1 = +5;
				 l_2 = -9; end
		240: begin l_1 = -5;
				 l_2 = +9; end
		383: begin l_1 = -5;
				 l_2 = -9; end
		528: begin l_1 = +1;
				 l_2 = -8; end
		159: begin l_1 = +5;
				 l_2 = -10; end
		496: begin l_1 = -5;
				 l_2 = +10; end
		127: begin l_1 = -1;
				 l_2 = +8; end
		385: begin l_1 = +5;
				 l_2 = +11; end
		302: begin l_1 = +5;
				 l_2 = -11; end
		353: begin l_1 = -5;
				 l_2 = +11; end
		270: begin l_1 = -5;
				 l_2 = -11; end
		99: begin l_1 = +5;
				 l_2 = +12; end
		588: begin l_1 = +5;
				 l_2 = -12; end
		67: begin l_1 = -5;
				 l_2 = +12; end
		556: begin l_1 = -5;
				 l_2 = -12; end
		182: begin l_1 = +5;
				 l_2 = +13; end
		505: begin l_1 = +5;
				 l_2 = -13; end
		150: begin l_1 = -5;
				 l_2 = +13; end
		473: begin l_1 = -5;
				 l_2 = -13; end
		348: begin l_1 = +5;
				 l_2 = +14; end
		339: begin l_1 = +5;
				 l_2 = -14; end
		316: begin l_1 = -5;
				 l_2 = +14; end
		307: begin l_1 = -5;
				 l_2 = -14; end
		96: begin l_1 = -6;
				 l_2 = +8; end
		559: begin l_1 = -6;
				 l_2 = -7; end
		160: begin l_1 = +6;
				 l_2 = +8; end
		495: begin l_1 = -6;
				 l_2 = -8; end
		288: begin l_1 = +2;
				 l_2 = -11; end
		431: begin l_1 = +6;
				 l_2 = -9; end
		224: begin l_1 = -6;
				 l_2 = +9; end
		367: begin l_1 = -2;
				 l_2 = +11; end
		544: begin l_1 = +6;
				 l_2 = +10; end
		175: begin l_1 = +6;
				 l_2 = -10; end
		480: begin l_1 = -6;
				 l_2 = +10; end
		111: begin l_1 = -6;
				 l_2 = -10; end
		401: begin l_1 = +2;
				 l_2 = -9; end
		318: begin l_1 = +6;
				 l_2 = -11; end
		337: begin l_1 = -6;
				 l_2 = +11; end
		254: begin l_1 = -2;
				 l_2 = +9; end
		115: begin l_1 = +6;
				 l_2 = +12; end
		604: begin l_1 = +6;
				 l_2 = -12; end
		51: begin l_1 = -6;
				 l_2 = +12; end
		540: begin l_1 = -6;
				 l_2 = -12; end
		198: begin l_1 = +6;
				 l_2 = +13; end
		521: begin l_1 = +6;
				 l_2 = -13; end
		134: begin l_1 = -6;
				 l_2 = +13; end
		457: begin l_1 = -6;
				 l_2 = -13; end
		364: begin l_1 = +6;
				 l_2 = +14; end
		355: begin l_1 = +6;
				 l_2 = -14; end
		300: begin l_1 = -6;
				 l_2 = +14; end
		291: begin l_1 = -6;
				 l_2 = -14; end
		192: begin l_1 = -7;
				 l_2 = +9; end
		463: begin l_1 = -7;
				 l_2 = -8; end
		320: begin l_1 = +7;
				 l_2 = +9; end
		335: begin l_1 = -7;
				 l_2 = -9; end
		576: begin l_1 = +3;
				 l_2 = -12; end
		207: begin l_1 = +7;
				 l_2 = -10; end
		448: begin l_1 = -7;
				 l_2 = +10; end
		79: begin l_1 = -3;
				 l_2 = +12; end
		433: begin l_1 = +7;
				 l_2 = +11; end
		350: begin l_1 = +7;
				 l_2 = -11; end
		305: begin l_1 = -7;
				 l_2 = +11; end
		222: begin l_1 = -7;
				 l_2 = -11; end
		147: begin l_1 = +3;
				 l_2 = -10; end
		636: begin l_1 = +7;
				 l_2 = -12; end
		19: begin l_1 = -7;
				 l_2 = +12; end
		508: begin l_1 = -3;
				 l_2 = +10; end
		230: begin l_1 = +7;
				 l_2 = +13; end
		553: begin l_1 = +7;
				 l_2 = -13; end
		102: begin l_1 = -7;
				 l_2 = +13; end
		425: begin l_1 = -7;
				 l_2 = -13; end
		396: begin l_1 = +7;
				 l_2 = +14; end
		387: begin l_1 = +7;
				 l_2 = -14; end
		268: begin l_1 = -7;
				 l_2 = +14; end
		259: begin l_1 = -7;
				 l_2 = -14; end
		384: begin l_1 = -8;
				 l_2 = +10; end
		271: begin l_1 = -8;
				 l_2 = -9; end
		640: begin l_1 = +1;
				 l_2 = -5; end
		15: begin l_1 = -1;
				 l_2 = +5; end
		497: begin l_1 = +4;
				 l_2 = -13; end
		414: begin l_1 = +8;
				 l_2 = -11; end
		241: begin l_1 = -8;
				 l_2 = +11; end
		158: begin l_1 = -4;
				 l_2 = +13; end
		211: begin l_1 = +8;
				 l_2 = +12; end
		45: begin l_1 = +8;
				 l_2 = -12; end
		610: begin l_1 = -8;
				 l_2 = +12; end
		444: begin l_1 = -8;
				 l_2 = -12; end
		294: begin l_1 = +4;
				 l_2 = -11; end
		617: begin l_1 = +8;
				 l_2 = -13; end
		38: begin l_1 = -8;
				 l_2 = +13; end
		361: begin l_1 = -4;
				 l_2 = +11; end
		460: begin l_1 = +8;
				 l_2 = +14; end
		451: begin l_1 = +8;
				 l_2 = -14; end
		204: begin l_1 = -8;
				 l_2 = +14; end
		195: begin l_1 = -8;
				 l_2 = -14; end
		113: begin l_1 = -9;
				 l_2 = +11; end
		542: begin l_1 = -9;
				 l_2 = -10; end
		625: begin l_1 = +2;
				 l_2 = -6; end
		30: begin l_1 = -2;
				 l_2 = +6; end
		339: begin l_1 = +5;
				 l_2 = -14; end
		173: begin l_1 = +9;
				 l_2 = -12; end
		482: begin l_1 = -9;
				 l_2 = +12; end
		316: begin l_1 = -5;
				 l_2 = +14; end
		422: begin l_1 = +9;
				 l_2 = +13; end
		90: begin l_1 = +9;
				 l_2 = -13; end
		565: begin l_1 = -9;
				 l_2 = +13; end
		233: begin l_1 = -9;
				 l_2 = -13; end
		588: begin l_1 = +5;
				 l_2 = -12; end
		579: begin l_1 = +9;
				 l_2 = -14; end
		76: begin l_1 = -9;
				 l_2 = +14; end
		67: begin l_1 = -5;
				 l_2 = +12; end
		226: begin l_1 = -10;
				 l_2 = +12; end
		429: begin l_1 = -10;
				 l_2 = -11; end
		595: begin l_1 = +3;
				 l_2 = -7; end
		60: begin l_1 = -3;
				 l_2 = +7; end
		23: begin l_1 = +10;
				 l_2 = +13; end
		346: begin l_1 = +10;
				 l_2 = -13; end
		309: begin l_1 = -10;
				 l_2 = +13; end
		632: begin l_1 = -10;
				 l_2 = -13; end
		189: begin l_1 = +10;
				 l_2 = +14; end
		180: begin l_1 = +10;
				 l_2 = -14; end
		475: begin l_1 = -10;
				 l_2 = +14; end
		466: begin l_1 = -10;
				 l_2 = -14; end
		452: begin l_1 = -11;
				 l_2 = +13; end
		203: begin l_1 = -11;
				 l_2 = -12; end
		535: begin l_1 = +4;
				 l_2 = -8; end
		120: begin l_1 = -4;
				 l_2 = +8; end
		46: begin l_1 = +11;
				 l_2 = +14; end
		37: begin l_1 = +11;
				 l_2 = -14; end
		618: begin l_1 = -11;
				 l_2 = +14; end
		609: begin l_1 = -11;
				 l_2 = -14; end
		249: begin l_1 = -12;
				 l_2 = +14; end
		406: begin l_1 = -12;
				 l_2 = -13; end
		415: begin l_1 = +5;
				 l_2 = -9; end
		240: begin l_1 = -5;
				 l_2 = +9; end
		498: begin l_1 = +13;
				 l_2 = +14; end
		157: begin l_1 = -13;
				 l_2 = -14; end
		default: begin l_1 = 0;
					   l_2 = 0; end
	endcase
end

endmodule

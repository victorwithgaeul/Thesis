// Product (AN) Code SEC r-LUT
// SEC_rLUT52bits.v
// Received remainder r, output single error location.
module SEC_rLUT52bits(r, l);
input 	[15:0]	r;
output	reg	signed	[7:0]	l;
always@(*) begin
	case(r)
		1: l = +1;
		50860: l = -1;
		2: l = +2;
		50859: l = -2;
		4: l = +3;
		50857: l = -3;
		8: l = +4;
		50853: l = -4;
		16: l = +5;
		50845: l = -5;
		32: l = +6;
		50829: l = -6;
		64: l = +7;
		50797: l = -7;
		128: l = +8;
		50733: l = -8;
		256: l = +9;
		50605: l = -9;
		512: l = +10;
		50349: l = -10;
		1024: l = +11;
		49837: l = -11;
		2048: l = +12;
		48813: l = -12;
		4096: l = +13;
		46765: l = -13;
		8192: l = +14;
		42669: l = -14;
		16384: l = +15;
		34477: l = -15;
		32768: l = +16;
		18093: l = -16;
		14675: l = +17;
		36186: l = -17;
		29350: l = +18;
		21511: l = -18;
		7839: l = +19;
		43022: l = -19;
		15678: l = +20;
		35183: l = -20;
		31356: l = +21;
		19505: l = -21;
		11851: l = +22;
		39010: l = -22;
		23702: l = +23;
		27159: l = -23;
		47404: l = +24;
		3457: l = -24;
		43947: l = +25;
		6914: l = -25;
		37033: l = +26;
		13828: l = -26;
		23205: l = +27;
		27656: l = -27;
		46410: l = +28;
		4451: l = -28;
		41959: l = +29;
		8902: l = -29;
		33057: l = +30;
		17804: l = -30;
		15253: l = +31;
		35608: l = -31;
		30506: l = +32;
		20355: l = -32;
		10151: l = +33;
		40710: l = -33;
		20302: l = +34;
		30559: l = -34;
		40604: l = +35;
		10257: l = -35;
		30347: l = +36;
		20514: l = -36;
		9833: l = +37;
		41028: l = -37;
		19666: l = +38;
		31195: l = -38;
		39332: l = +39;
		11529: l = -39;
		27803: l = +40;
		23058: l = -40;
		4745: l = +41;
		46116: l = -41;
		9490: l = +42;
		41371: l = -42;
		18980: l = +43;
		31881: l = -43;
		37960: l = +44;
		12901: l = -44;
		25059: l = +45;
		25802: l = -45;
		50118: l = +46;
		743: l = -46;
		49375: l = +47;
		1486: l = -47;
		47889: l = +48;
		2972: l = -48;
		44917: l = +49;
		5944: l = -49;
		38973: l = +50;
		11888: l = -50;
		27085: l = +51;
		23776: l = -51;
		3309: l = +52;
		47552: l = -52;
		6618: l = +53;
		44243: l = -53;
		13236: l = +54;
		37625: l = -54;
		26472: l = +55;
		24389: l = -55;
		2083: l = +56;
		48778: l = -56;
		4166: l = +57;
		46695: l = -57;
		8332: l = +58;
		42529: l = -58;
		16664: l = +59;
		34197: l = -59;
		33328: l = +60;
		17533: l = -60;
		15795: l = +61;
		35066: l = -61;
		31590: l = +62;
		19271: l = -62;
		12319: l = +63;
		38542: l = -63;
		24638: l = +64;
		26223: l = -64;
		49276: l = +65;
		1585: l = -65;
		47691: l = +66;
		3170: l = -66;
		44521: l = +67;
		6340: l = -67;
		38181: l = +68;
		12680: l = -68;
		default: l = 0;
	endcase
end

endmodule

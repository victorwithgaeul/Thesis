// Product (AN) Code DEC r-LUT
// DEC_rLUT28bits.v
// Used to do DEC, but corrected errors by locations, not AWE
// Received remainder r, output two error locations.
module DEC_rLUT28bits(r, l_1, l_2);
input 	[14:0]	r;
output	reg	signed	[6:0]	l_1;
output	reg	signed	[6:0]	l_2;
always@(*) begin
	case(r)
		1: begin l_1 = -1;
				 l_2 = +2; end
		17618: begin l_1 = +1;
				 l_2 = -2; end
		2: begin l_1 = +1;
				 l_2 = +1; end
		17617: begin l_1 = -1;
				 l_2 = -1; end
		4: begin l_1 = +2;
				 l_2 = +2; end
		17615: begin l_1 = -2;
				 l_2 = -2; end
		8: begin l_1 = +3;
				 l_2 = +3; end
		17611: begin l_1 = -3;
				 l_2 = -3; end
		16: begin l_1 = +4;
				 l_2 = +4; end
		17603: begin l_1 = -4;
				 l_2 = -4; end
		32: begin l_1 = +5;
				 l_2 = +5; end
		17587: begin l_1 = -5;
				 l_2 = -5; end
		64: begin l_1 = +6;
				 l_2 = +6; end
		17555: begin l_1 = -6;
				 l_2 = -6; end
		128: begin l_1 = +7;
				 l_2 = +7; end
		17491: begin l_1 = -7;
				 l_2 = -7; end
		256: begin l_1 = +8;
				 l_2 = +8; end
		17363: begin l_1 = -8;
				 l_2 = -8; end
		512: begin l_1 = +9;
				 l_2 = +9; end
		17107: begin l_1 = -9;
				 l_2 = -9; end
		1024: begin l_1 = +10;
				 l_2 = +10; end
		16595: begin l_1 = -10;
				 l_2 = -10; end
		2048: begin l_1 = +11;
				 l_2 = +11; end
		15571: begin l_1 = -11;
				 l_2 = -11; end
		4096: begin l_1 = +12;
				 l_2 = +12; end
		13523: begin l_1 = -12;
				 l_2 = -12; end
		8192: begin l_1 = +13;
				 l_2 = +13; end
		9427: begin l_1 = -13;
				 l_2 = -13; end
		16384: begin l_1 = +14;
				 l_2 = +14; end
		1235: begin l_1 = -14;
				 l_2 = -14; end
		15149: begin l_1 = +15;
				 l_2 = +15; end
		2470: begin l_1 = -15;
				 l_2 = -15; end
		12679: begin l_1 = +16;
				 l_2 = +16; end
		4940: begin l_1 = -16;
				 l_2 = -16; end
		7739: begin l_1 = +17;
				 l_2 = +17; end
		9880: begin l_1 = -17;
				 l_2 = -17; end
		15478: begin l_1 = +18;
				 l_2 = +18; end
		2141: begin l_1 = -18;
				 l_2 = -18; end
		13337: begin l_1 = +19;
				 l_2 = +19; end
		4282: begin l_1 = -19;
				 l_2 = -19; end
		9055: begin l_1 = +20;
				 l_2 = +20; end
		8564: begin l_1 = -20;
				 l_2 = -20; end
		491: begin l_1 = +21;
				 l_2 = +21; end
		17128: begin l_1 = -21;
				 l_2 = -21; end
		982: begin l_1 = +22;
				 l_2 = +22; end
		16637: begin l_1 = -22;
				 l_2 = -22; end
		1964: begin l_1 = +23;
				 l_2 = +23; end
		15655: begin l_1 = -23;
				 l_2 = -23; end
		3928: begin l_1 = +24;
				 l_2 = +24; end
		13691: begin l_1 = -24;
				 l_2 = -24; end
		7856: begin l_1 = +25;
				 l_2 = +25; end
		9763: begin l_1 = -25;
				 l_2 = -25; end
		15712: begin l_1 = +26;
				 l_2 = +26; end
		1907: begin l_1 = -26;
				 l_2 = -26; end
		13805: begin l_1 = +27;
				 l_2 = +27; end
		3814: begin l_1 = -27;
				 l_2 = -27; end
		9991: begin l_1 = +28;
				 l_2 = +28; end
		7628: begin l_1 = -28;
				 l_2 = -28; end
		2363: begin l_1 = +29;
				 l_2 = +29; end
		15256: begin l_1 = -29;
				 l_2 = -29; end
		4726: begin l_1 = +30;
				 l_2 = +30; end
		12893: begin l_1 = -30;
				 l_2 = -30; end
		9452: begin l_1 = +31;
				 l_2 = +31; end
		8167: begin l_1 = -31;
				 l_2 = -31; end
		1285: begin l_1 = +32;
				 l_2 = +32; end
		16334: begin l_1 = -32;
				 l_2 = -32; end
		2570: begin l_1 = +33;
				 l_2 = +33; end
		15049: begin l_1 = -33;
				 l_2 = -33; end
		5140: begin l_1 = +34;
				 l_2 = +34; end
		12479: begin l_1 = -34;
				 l_2 = -34; end
		10280: begin l_1 = +35;
				 l_2 = +35; end
		7339: begin l_1 = -35;
				 l_2 = -35; end
		2941: begin l_1 = +36;
				 l_2 = +36; end
		14678: begin l_1 = -36;
				 l_2 = -36; end
		5882: begin l_1 = +37;
				 l_2 = +37; end
		11737: begin l_1 = -37;
				 l_2 = -37; end
		11764: begin l_1 = +38;
				 l_2 = +38; end
		5855: begin l_1 = -38;
				 l_2 = -38; end
		5909: begin l_1 = +39;
				 l_2 = +39; end
		11710: begin l_1 = -39;
				 l_2 = -39; end
		11818: begin l_1 = +40;
				 l_2 = +40; end
		5801: begin l_1 = -40;
				 l_2 = -40; end
		6017: begin l_1 = +41;
				 l_2 = +41; end
		11602: begin l_1 = -41;
				 l_2 = -41; end
		12034: begin l_1 = +42;
				 l_2 = +42; end
		5585: begin l_1 = -42;
				 l_2 = -42; end
		3: begin l_1 = -1;
				 l_2 = +3; end
		17616: begin l_1 = -1;
				 l_2 = -2; end
		5: begin l_1 = +1;
				 l_2 = +3; end
		17614: begin l_1 = -1;
				 l_2 = -3; end
		9: begin l_1 = +1;
				 l_2 = +4; end
		17612: begin l_1 = +1;
				 l_2 = -4; end
		7: begin l_1 = -1;
				 l_2 = +4; end
		17610: begin l_1 = -1;
				 l_2 = -4; end
		17: begin l_1 = +1;
				 l_2 = +5; end
		17604: begin l_1 = +1;
				 l_2 = -5; end
		15: begin l_1 = -1;
				 l_2 = +5; end
		17602: begin l_1 = -1;
				 l_2 = -5; end
		33: begin l_1 = +1;
				 l_2 = +6; end
		17588: begin l_1 = +1;
				 l_2 = -6; end
		31: begin l_1 = -1;
				 l_2 = +6; end
		17586: begin l_1 = -1;
				 l_2 = -6; end
		65: begin l_1 = +1;
				 l_2 = +7; end
		17556: begin l_1 = +1;
				 l_2 = -7; end
		63: begin l_1 = -1;
				 l_2 = +7; end
		17554: begin l_1 = -1;
				 l_2 = -7; end
		129: begin l_1 = +1;
				 l_2 = +8; end
		17492: begin l_1 = +1;
				 l_2 = -8; end
		127: begin l_1 = -1;
				 l_2 = +8; end
		17490: begin l_1 = -1;
				 l_2 = -8; end
		257: begin l_1 = +1;
				 l_2 = +9; end
		17364: begin l_1 = +1;
				 l_2 = -9; end
		255: begin l_1 = -1;
				 l_2 = +9; end
		17362: begin l_1 = -1;
				 l_2 = -9; end
		513: begin l_1 = +1;
				 l_2 = +10; end
		17108: begin l_1 = +1;
				 l_2 = -10; end
		511: begin l_1 = -1;
				 l_2 = +10; end
		17106: begin l_1 = -1;
				 l_2 = -10; end
		1025: begin l_1 = +1;
				 l_2 = +11; end
		16596: begin l_1 = +1;
				 l_2 = -11; end
		1023: begin l_1 = -1;
				 l_2 = +11; end
		16594: begin l_1 = -1;
				 l_2 = -11; end
		2049: begin l_1 = +1;
				 l_2 = +12; end
		15572: begin l_1 = +1;
				 l_2 = -12; end
		2047: begin l_1 = -1;
				 l_2 = +12; end
		15570: begin l_1 = -1;
				 l_2 = -12; end
		4097: begin l_1 = +1;
				 l_2 = +13; end
		13524: begin l_1 = +1;
				 l_2 = -13; end
		4095: begin l_1 = -1;
				 l_2 = +13; end
		13522: begin l_1 = -1;
				 l_2 = -13; end
		8193: begin l_1 = +1;
				 l_2 = +14; end
		9428: begin l_1 = +1;
				 l_2 = -14; end
		8191: begin l_1 = -1;
				 l_2 = +14; end
		9426: begin l_1 = -1;
				 l_2 = -14; end
		16385: begin l_1 = +1;
				 l_2 = +15; end
		1236: begin l_1 = +1;
				 l_2 = -15; end
		16383: begin l_1 = -1;
				 l_2 = +15; end
		1234: begin l_1 = -1;
				 l_2 = -15; end
		15150: begin l_1 = +1;
				 l_2 = +16; end
		2471: begin l_1 = +1;
				 l_2 = -16; end
		15148: begin l_1 = -1;
				 l_2 = +16; end
		2469: begin l_1 = -1;
				 l_2 = -16; end
		12680: begin l_1 = +1;
				 l_2 = +17; end
		4941: begin l_1 = +1;
				 l_2 = -17; end
		12678: begin l_1 = -1;
				 l_2 = +17; end
		4939: begin l_1 = -1;
				 l_2 = -17; end
		7740: begin l_1 = +1;
				 l_2 = +18; end
		9881: begin l_1 = +1;
				 l_2 = -18; end
		7738: begin l_1 = -1;
				 l_2 = +18; end
		9879: begin l_1 = -1;
				 l_2 = -18; end
		15479: begin l_1 = +1;
				 l_2 = +19; end
		2142: begin l_1 = +1;
				 l_2 = -19; end
		15477: begin l_1 = -1;
				 l_2 = +19; end
		2140: begin l_1 = -1;
				 l_2 = -19; end
		13338: begin l_1 = +1;
				 l_2 = +20; end
		4283: begin l_1 = +1;
				 l_2 = -20; end
		13336: begin l_1 = -1;
				 l_2 = +20; end
		4281: begin l_1 = -1;
				 l_2 = -20; end
		9056: begin l_1 = +1;
				 l_2 = +21; end
		8565: begin l_1 = +1;
				 l_2 = -21; end
		9054: begin l_1 = -1;
				 l_2 = +21; end
		8563: begin l_1 = -1;
				 l_2 = -21; end
		492: begin l_1 = +1;
				 l_2 = +22; end
		17129: begin l_1 = +1;
				 l_2 = -22; end
		490: begin l_1 = -1;
				 l_2 = +22; end
		17127: begin l_1 = -1;
				 l_2 = -22; end
		983: begin l_1 = +1;
				 l_2 = +23; end
		16638: begin l_1 = +1;
				 l_2 = -23; end
		981: begin l_1 = -1;
				 l_2 = +23; end
		16636: begin l_1 = -1;
				 l_2 = -23; end
		1965: begin l_1 = +1;
				 l_2 = +24; end
		15656: begin l_1 = +1;
				 l_2 = -24; end
		1963: begin l_1 = -1;
				 l_2 = +24; end
		15654: begin l_1 = -1;
				 l_2 = -24; end
		3929: begin l_1 = +1;
				 l_2 = +25; end
		13692: begin l_1 = +1;
				 l_2 = -25; end
		3927: begin l_1 = -1;
				 l_2 = +25; end
		13690: begin l_1 = -1;
				 l_2 = -25; end
		7857: begin l_1 = +1;
				 l_2 = +26; end
		9764: begin l_1 = +1;
				 l_2 = -26; end
		7855: begin l_1 = -1;
				 l_2 = +26; end
		9762: begin l_1 = -1;
				 l_2 = -26; end
		15713: begin l_1 = +1;
				 l_2 = +27; end
		1908: begin l_1 = +1;
				 l_2 = -27; end
		15711: begin l_1 = -1;
				 l_2 = +27; end
		1906: begin l_1 = -1;
				 l_2 = -27; end
		13806: begin l_1 = +1;
				 l_2 = +28; end
		3815: begin l_1 = +1;
				 l_2 = -28; end
		13804: begin l_1 = -1;
				 l_2 = +28; end
		3813: begin l_1 = -1;
				 l_2 = -28; end
		9992: begin l_1 = +1;
				 l_2 = +29; end
		7629: begin l_1 = +1;
				 l_2 = -29; end
		9990: begin l_1 = -1;
				 l_2 = +29; end
		7627: begin l_1 = -1;
				 l_2 = -29; end
		2364: begin l_1 = +1;
				 l_2 = +30; end
		15257: begin l_1 = +1;
				 l_2 = -30; end
		2362: begin l_1 = -1;
				 l_2 = +30; end
		15255: begin l_1 = -1;
				 l_2 = -30; end
		4727: begin l_1 = +1;
				 l_2 = +31; end
		12894: begin l_1 = +1;
				 l_2 = -31; end
		4725: begin l_1 = -1;
				 l_2 = +31; end
		12892: begin l_1 = -1;
				 l_2 = -31; end
		9453: begin l_1 = +1;
				 l_2 = +32; end
		8168: begin l_1 = +1;
				 l_2 = -32; end
		9451: begin l_1 = -1;
				 l_2 = +32; end
		8166: begin l_1 = -1;
				 l_2 = -32; end
		1286: begin l_1 = +1;
				 l_2 = +33; end
		16335: begin l_1 = +1;
				 l_2 = -33; end
		1284: begin l_1 = -1;
				 l_2 = +33; end
		16333: begin l_1 = -1;
				 l_2 = -33; end
		2571: begin l_1 = +1;
				 l_2 = +34; end
		15050: begin l_1 = +1;
				 l_2 = -34; end
		2569: begin l_1 = -1;
				 l_2 = +34; end
		15048: begin l_1 = -1;
				 l_2 = -34; end
		5141: begin l_1 = +1;
				 l_2 = +35; end
		12480: begin l_1 = +1;
				 l_2 = -35; end
		5139: begin l_1 = -1;
				 l_2 = +35; end
		12478: begin l_1 = -1;
				 l_2 = -35; end
		10281: begin l_1 = +1;
				 l_2 = +36; end
		7340: begin l_1 = +1;
				 l_2 = -36; end
		10279: begin l_1 = -1;
				 l_2 = +36; end
		7338: begin l_1 = -1;
				 l_2 = -36; end
		2942: begin l_1 = +1;
				 l_2 = +37; end
		14679: begin l_1 = +1;
				 l_2 = -37; end
		2940: begin l_1 = -1;
				 l_2 = +37; end
		14677: begin l_1 = -1;
				 l_2 = -37; end
		5883: begin l_1 = +1;
				 l_2 = +38; end
		11738: begin l_1 = +1;
				 l_2 = -38; end
		5881: begin l_1 = -1;
				 l_2 = +38; end
		11736: begin l_1 = -1;
				 l_2 = -38; end
		11765: begin l_1 = +1;
				 l_2 = +39; end
		5856: begin l_1 = +1;
				 l_2 = -39; end
		11763: begin l_1 = -1;
				 l_2 = +39; end
		5854: begin l_1 = -1;
				 l_2 = -39; end
		5910: begin l_1 = +1;
				 l_2 = +40; end
		11711: begin l_1 = +1;
				 l_2 = -40; end
		5908: begin l_1 = -1;
				 l_2 = +40; end
		11709: begin l_1 = -1;
				 l_2 = -40; end
		11819: begin l_1 = +1;
				 l_2 = +41; end
		5802: begin l_1 = +1;
				 l_2 = -41; end
		11817: begin l_1 = -1;
				 l_2 = +41; end
		5800: begin l_1 = -1;
				 l_2 = -41; end
		6018: begin l_1 = +1;
				 l_2 = +42; end
		11603: begin l_1 = +1;
				 l_2 = -42; end
		6016: begin l_1 = -1;
				 l_2 = +42; end
		11601: begin l_1 = -1;
				 l_2 = -42; end
		12035: begin l_1 = +1;
				 l_2 = +43; end
		5586: begin l_1 = +1;
				 l_2 = -43; end
		12033: begin l_1 = -1;
				 l_2 = +43; end
		5584: begin l_1 = -1;
				 l_2 = -43; end
		6: begin l_1 = -2;
				 l_2 = +4; end
		17613: begin l_1 = -2;
				 l_2 = -3; end
		10: begin l_1 = +2;
				 l_2 = +4; end
		17609: begin l_1 = -2;
				 l_2 = -4; end
		18: begin l_1 = +2;
				 l_2 = +5; end
		17605: begin l_1 = +2;
				 l_2 = -5; end
		14: begin l_1 = -2;
				 l_2 = +5; end
		17601: begin l_1 = -2;
				 l_2 = -5; end
		34: begin l_1 = +2;
				 l_2 = +6; end
		17589: begin l_1 = +2;
				 l_2 = -6; end
		30: begin l_1 = -2;
				 l_2 = +6; end
		17585: begin l_1 = -2;
				 l_2 = -6; end
		66: begin l_1 = +2;
				 l_2 = +7; end
		17557: begin l_1 = +2;
				 l_2 = -7; end
		62: begin l_1 = -2;
				 l_2 = +7; end
		17553: begin l_1 = -2;
				 l_2 = -7; end
		130: begin l_1 = +2;
				 l_2 = +8; end
		17493: begin l_1 = +2;
				 l_2 = -8; end
		126: begin l_1 = -2;
				 l_2 = +8; end
		17489: begin l_1 = -2;
				 l_2 = -8; end
		258: begin l_1 = +2;
				 l_2 = +9; end
		17365: begin l_1 = +2;
				 l_2 = -9; end
		254: begin l_1 = -2;
				 l_2 = +9; end
		17361: begin l_1 = -2;
				 l_2 = -9; end
		514: begin l_1 = +2;
				 l_2 = +10; end
		17109: begin l_1 = +2;
				 l_2 = -10; end
		510: begin l_1 = -2;
				 l_2 = +10; end
		17105: begin l_1 = -2;
				 l_2 = -10; end
		1026: begin l_1 = +2;
				 l_2 = +11; end
		16597: begin l_1 = +2;
				 l_2 = -11; end
		1022: begin l_1 = -2;
				 l_2 = +11; end
		16593: begin l_1 = -2;
				 l_2 = -11; end
		2050: begin l_1 = +2;
				 l_2 = +12; end
		15573: begin l_1 = +2;
				 l_2 = -12; end
		2046: begin l_1 = -2;
				 l_2 = +12; end
		15569: begin l_1 = -2;
				 l_2 = -12; end
		4098: begin l_1 = +2;
				 l_2 = +13; end
		13525: begin l_1 = +2;
				 l_2 = -13; end
		4094: begin l_1 = -2;
				 l_2 = +13; end
		13521: begin l_1 = -2;
				 l_2 = -13; end
		8194: begin l_1 = +2;
				 l_2 = +14; end
		9429: begin l_1 = +2;
				 l_2 = -14; end
		8190: begin l_1 = -2;
				 l_2 = +14; end
		9425: begin l_1 = -2;
				 l_2 = -14; end
		16386: begin l_1 = +2;
				 l_2 = +15; end
		1237: begin l_1 = +2;
				 l_2 = -15; end
		16382: begin l_1 = -2;
				 l_2 = +15; end
		1233: begin l_1 = -2;
				 l_2 = -15; end
		15151: begin l_1 = +2;
				 l_2 = +16; end
		2472: begin l_1 = +2;
				 l_2 = -16; end
		15147: begin l_1 = -2;
				 l_2 = +16; end
		2468: begin l_1 = -2;
				 l_2 = -16; end
		12681: begin l_1 = +2;
				 l_2 = +17; end
		4942: begin l_1 = +2;
				 l_2 = -17; end
		12677: begin l_1 = -2;
				 l_2 = +17; end
		4938: begin l_1 = -2;
				 l_2 = -17; end
		7741: begin l_1 = +2;
				 l_2 = +18; end
		9882: begin l_1 = +2;
				 l_2 = -18; end
		7737: begin l_1 = -2;
				 l_2 = +18; end
		9878: begin l_1 = -2;
				 l_2 = -18; end
		15480: begin l_1 = +2;
				 l_2 = +19; end
		2143: begin l_1 = +2;
				 l_2 = -19; end
		15476: begin l_1 = -2;
				 l_2 = +19; end
		2139: begin l_1 = -2;
				 l_2 = -19; end
		13339: begin l_1 = +2;
				 l_2 = +20; end
		4284: begin l_1 = +2;
				 l_2 = -20; end
		13335: begin l_1 = -2;
				 l_2 = +20; end
		4280: begin l_1 = -2;
				 l_2 = -20; end
		9057: begin l_1 = +2;
				 l_2 = +21; end
		8566: begin l_1 = +2;
				 l_2 = -21; end
		9053: begin l_1 = -2;
				 l_2 = +21; end
		8562: begin l_1 = -2;
				 l_2 = -21; end
		493: begin l_1 = +2;
				 l_2 = +22; end
		17130: begin l_1 = +2;
				 l_2 = -22; end
		489: begin l_1 = -2;
				 l_2 = +22; end
		17126: begin l_1 = -2;
				 l_2 = -22; end
		984: begin l_1 = +2;
				 l_2 = +23; end
		16639: begin l_1 = +2;
				 l_2 = -23; end
		980: begin l_1 = -2;
				 l_2 = +23; end
		16635: begin l_1 = -2;
				 l_2 = -23; end
		1966: begin l_1 = +2;
				 l_2 = +24; end
		15657: begin l_1 = +2;
				 l_2 = -24; end
		1962: begin l_1 = -2;
				 l_2 = +24; end
		15653: begin l_1 = -2;
				 l_2 = -24; end
		3930: begin l_1 = +2;
				 l_2 = +25; end
		13693: begin l_1 = +2;
				 l_2 = -25; end
		3926: begin l_1 = -2;
				 l_2 = +25; end
		13689: begin l_1 = -2;
				 l_2 = -25; end
		7858: begin l_1 = +2;
				 l_2 = +26; end
		9765: begin l_1 = +2;
				 l_2 = -26; end
		7854: begin l_1 = -2;
				 l_2 = +26; end
		9761: begin l_1 = -2;
				 l_2 = -26; end
		15714: begin l_1 = +2;
				 l_2 = +27; end
		1909: begin l_1 = +2;
				 l_2 = -27; end
		15710: begin l_1 = -2;
				 l_2 = +27; end
		1905: begin l_1 = -2;
				 l_2 = -27; end
		13807: begin l_1 = +2;
				 l_2 = +28; end
		3816: begin l_1 = +2;
				 l_2 = -28; end
		13803: begin l_1 = -2;
				 l_2 = +28; end
		3812: begin l_1 = -2;
				 l_2 = -28; end
		9993: begin l_1 = +2;
				 l_2 = +29; end
		7630: begin l_1 = +2;
				 l_2 = -29; end
		9989: begin l_1 = -2;
				 l_2 = +29; end
		7626: begin l_1 = -2;
				 l_2 = -29; end
		2365: begin l_1 = +2;
				 l_2 = +30; end
		15258: begin l_1 = +2;
				 l_2 = -30; end
		2361: begin l_1 = -2;
				 l_2 = +30; end
		15254: begin l_1 = -2;
				 l_2 = -30; end
		4728: begin l_1 = +2;
				 l_2 = +31; end
		12895: begin l_1 = +2;
				 l_2 = -31; end
		4724: begin l_1 = -2;
				 l_2 = +31; end
		12891: begin l_1 = -2;
				 l_2 = -31; end
		9454: begin l_1 = +2;
				 l_2 = +32; end
		8169: begin l_1 = +2;
				 l_2 = -32; end
		9450: begin l_1 = -2;
				 l_2 = +32; end
		8165: begin l_1 = -2;
				 l_2 = -32; end
		1287: begin l_1 = +2;
				 l_2 = +33; end
		16336: begin l_1 = +2;
				 l_2 = -33; end
		1283: begin l_1 = -2;
				 l_2 = +33; end
		16332: begin l_1 = -2;
				 l_2 = -33; end
		2572: begin l_1 = +2;
				 l_2 = +34; end
		15051: begin l_1 = +2;
				 l_2 = -34; end
		2568: begin l_1 = -2;
				 l_2 = +34; end
		15047: begin l_1 = -2;
				 l_2 = -34; end
		5142: begin l_1 = +2;
				 l_2 = +35; end
		12481: begin l_1 = +2;
				 l_2 = -35; end
		5138: begin l_1 = -2;
				 l_2 = +35; end
		12477: begin l_1 = -2;
				 l_2 = -35; end
		10282: begin l_1 = +2;
				 l_2 = +36; end
		7341: begin l_1 = +2;
				 l_2 = -36; end
		10278: begin l_1 = -2;
				 l_2 = +36; end
		7337: begin l_1 = -2;
				 l_2 = -36; end
		2943: begin l_1 = +2;
				 l_2 = +37; end
		14680: begin l_1 = +2;
				 l_2 = -37; end
		2939: begin l_1 = -2;
				 l_2 = +37; end
		14676: begin l_1 = -2;
				 l_2 = -37; end
		5884: begin l_1 = +2;
				 l_2 = +38; end
		11739: begin l_1 = +2;
				 l_2 = -38; end
		5880: begin l_1 = -2;
				 l_2 = +38; end
		11735: begin l_1 = -2;
				 l_2 = -38; end
		11766: begin l_1 = +2;
				 l_2 = +39; end
		5857: begin l_1 = +2;
				 l_2 = -39; end
		11762: begin l_1 = -2;
				 l_2 = +39; end
		5853: begin l_1 = -2;
				 l_2 = -39; end
		5911: begin l_1 = +2;
				 l_2 = +40; end
		11712: begin l_1 = +2;
				 l_2 = -40; end
		5907: begin l_1 = -2;
				 l_2 = +40; end
		11708: begin l_1 = -2;
				 l_2 = -40; end
		11820: begin l_1 = +2;
				 l_2 = +41; end
		5803: begin l_1 = +2;
				 l_2 = -41; end
		11816: begin l_1 = -2;
				 l_2 = +41; end
		5799: begin l_1 = -2;
				 l_2 = -41; end
		6019: begin l_1 = +2;
				 l_2 = +42; end
		11604: begin l_1 = +2;
				 l_2 = -42; end
		6015: begin l_1 = -2;
				 l_2 = +42; end
		11600: begin l_1 = -2;
				 l_2 = -42; end
		12036: begin l_1 = +2;
				 l_2 = +43; end
		5587: begin l_1 = +2;
				 l_2 = -43; end
		12032: begin l_1 = -2;
				 l_2 = +43; end
		5583: begin l_1 = -2;
				 l_2 = -43; end
		12: begin l_1 = -3;
				 l_2 = +5; end
		17607: begin l_1 = -3;
				 l_2 = -4; end
		20: begin l_1 = +3;
				 l_2 = +5; end
		17599: begin l_1 = -3;
				 l_2 = -5; end
		36: begin l_1 = +3;
				 l_2 = +6; end
		17591: begin l_1 = +3;
				 l_2 = -6; end
		28: begin l_1 = -3;
				 l_2 = +6; end
		17583: begin l_1 = -3;
				 l_2 = -6; end
		68: begin l_1 = +3;
				 l_2 = +7; end
		17559: begin l_1 = +3;
				 l_2 = -7; end
		60: begin l_1 = -3;
				 l_2 = +7; end
		17551: begin l_1 = -3;
				 l_2 = -7; end
		132: begin l_1 = +3;
				 l_2 = +8; end
		17495: begin l_1 = +3;
				 l_2 = -8; end
		124: begin l_1 = -3;
				 l_2 = +8; end
		17487: begin l_1 = -3;
				 l_2 = -8; end
		260: begin l_1 = +3;
				 l_2 = +9; end
		17367: begin l_1 = +3;
				 l_2 = -9; end
		252: begin l_1 = -3;
				 l_2 = +9; end
		17359: begin l_1 = -3;
				 l_2 = -9; end
		516: begin l_1 = +3;
				 l_2 = +10; end
		17111: begin l_1 = +3;
				 l_2 = -10; end
		508: begin l_1 = -3;
				 l_2 = +10; end
		17103: begin l_1 = -3;
				 l_2 = -10; end
		1028: begin l_1 = +3;
				 l_2 = +11; end
		16599: begin l_1 = +3;
				 l_2 = -11; end
		1020: begin l_1 = -3;
				 l_2 = +11; end
		16591: begin l_1 = -3;
				 l_2 = -11; end
		2052: begin l_1 = +3;
				 l_2 = +12; end
		15575: begin l_1 = +3;
				 l_2 = -12; end
		2044: begin l_1 = -3;
				 l_2 = +12; end
		15567: begin l_1 = -3;
				 l_2 = -12; end
		4100: begin l_1 = +3;
				 l_2 = +13; end
		13527: begin l_1 = +3;
				 l_2 = -13; end
		4092: begin l_1 = -3;
				 l_2 = +13; end
		13519: begin l_1 = -3;
				 l_2 = -13; end
		8196: begin l_1 = +3;
				 l_2 = +14; end
		9431: begin l_1 = +3;
				 l_2 = -14; end
		8188: begin l_1 = -3;
				 l_2 = +14; end
		9423: begin l_1 = -3;
				 l_2 = -14; end
		16388: begin l_1 = +3;
				 l_2 = +15; end
		1239: begin l_1 = +3;
				 l_2 = -15; end
		16380: begin l_1 = -3;
				 l_2 = +15; end
		1231: begin l_1 = -3;
				 l_2 = -15; end
		15153: begin l_1 = +3;
				 l_2 = +16; end
		2474: begin l_1 = +3;
				 l_2 = -16; end
		15145: begin l_1 = -3;
				 l_2 = +16; end
		2466: begin l_1 = -3;
				 l_2 = -16; end
		12683: begin l_1 = +3;
				 l_2 = +17; end
		4944: begin l_1 = +3;
				 l_2 = -17; end
		12675: begin l_1 = -3;
				 l_2 = +17; end
		4936: begin l_1 = -3;
				 l_2 = -17; end
		7743: begin l_1 = +3;
				 l_2 = +18; end
		9884: begin l_1 = +3;
				 l_2 = -18; end
		7735: begin l_1 = -3;
				 l_2 = +18; end
		9876: begin l_1 = -3;
				 l_2 = -18; end
		15482: begin l_1 = +3;
				 l_2 = +19; end
		2145: begin l_1 = +3;
				 l_2 = -19; end
		15474: begin l_1 = -3;
				 l_2 = +19; end
		2137: begin l_1 = -3;
				 l_2 = -19; end
		13341: begin l_1 = +3;
				 l_2 = +20; end
		4286: begin l_1 = +3;
				 l_2 = -20; end
		13333: begin l_1 = -3;
				 l_2 = +20; end
		4278: begin l_1 = -3;
				 l_2 = -20; end
		9059: begin l_1 = +3;
				 l_2 = +21; end
		8568: begin l_1 = +3;
				 l_2 = -21; end
		9051: begin l_1 = -3;
				 l_2 = +21; end
		8560: begin l_1 = -3;
				 l_2 = -21; end
		495: begin l_1 = +3;
				 l_2 = +22; end
		17132: begin l_1 = +3;
				 l_2 = -22; end
		487: begin l_1 = -3;
				 l_2 = +22; end
		17124: begin l_1 = -3;
				 l_2 = -22; end
		986: begin l_1 = +3;
				 l_2 = +23; end
		16641: begin l_1 = +3;
				 l_2 = -23; end
		978: begin l_1 = -3;
				 l_2 = +23; end
		16633: begin l_1 = -3;
				 l_2 = -23; end
		1968: begin l_1 = +3;
				 l_2 = +24; end
		15659: begin l_1 = +3;
				 l_2 = -24; end
		1960: begin l_1 = -3;
				 l_2 = +24; end
		15651: begin l_1 = -3;
				 l_2 = -24; end
		3932: begin l_1 = +3;
				 l_2 = +25; end
		13695: begin l_1 = +3;
				 l_2 = -25; end
		3924: begin l_1 = -3;
				 l_2 = +25; end
		13687: begin l_1 = -3;
				 l_2 = -25; end
		7860: begin l_1 = +3;
				 l_2 = +26; end
		9767: begin l_1 = +3;
				 l_2 = -26; end
		7852: begin l_1 = -3;
				 l_2 = +26; end
		9759: begin l_1 = -3;
				 l_2 = -26; end
		15716: begin l_1 = +3;
				 l_2 = +27; end
		1911: begin l_1 = +3;
				 l_2 = -27; end
		15708: begin l_1 = -3;
				 l_2 = +27; end
		1903: begin l_1 = -3;
				 l_2 = -27; end
		13809: begin l_1 = +3;
				 l_2 = +28; end
		3818: begin l_1 = +3;
				 l_2 = -28; end
		13801: begin l_1 = -3;
				 l_2 = +28; end
		3810: begin l_1 = -3;
				 l_2 = -28; end
		9995: begin l_1 = +3;
				 l_2 = +29; end
		7632: begin l_1 = +3;
				 l_2 = -29; end
		9987: begin l_1 = -3;
				 l_2 = +29; end
		7624: begin l_1 = -3;
				 l_2 = -29; end
		2367: begin l_1 = +3;
				 l_2 = +30; end
		15260: begin l_1 = +3;
				 l_2 = -30; end
		2359: begin l_1 = -3;
				 l_2 = +30; end
		15252: begin l_1 = -3;
				 l_2 = -30; end
		4730: begin l_1 = +3;
				 l_2 = +31; end
		12897: begin l_1 = +3;
				 l_2 = -31; end
		4722: begin l_1 = -3;
				 l_2 = +31; end
		12889: begin l_1 = -3;
				 l_2 = -31; end
		9456: begin l_1 = +3;
				 l_2 = +32; end
		8171: begin l_1 = +3;
				 l_2 = -32; end
		9448: begin l_1 = -3;
				 l_2 = +32; end
		8163: begin l_1 = -3;
				 l_2 = -32; end
		1289: begin l_1 = +3;
				 l_2 = +33; end
		16338: begin l_1 = +3;
				 l_2 = -33; end
		1281: begin l_1 = -3;
				 l_2 = +33; end
		16330: begin l_1 = -3;
				 l_2 = -33; end
		2574: begin l_1 = +3;
				 l_2 = +34; end
		15053: begin l_1 = +3;
				 l_2 = -34; end
		2566: begin l_1 = -3;
				 l_2 = +34; end
		15045: begin l_1 = -3;
				 l_2 = -34; end
		5144: begin l_1 = +3;
				 l_2 = +35; end
		12483: begin l_1 = +3;
				 l_2 = -35; end
		5136: begin l_1 = -3;
				 l_2 = +35; end
		12475: begin l_1 = -3;
				 l_2 = -35; end
		10284: begin l_1 = +3;
				 l_2 = +36; end
		7343: begin l_1 = +3;
				 l_2 = -36; end
		10276: begin l_1 = -3;
				 l_2 = +36; end
		7335: begin l_1 = -3;
				 l_2 = -36; end
		2945: begin l_1 = +3;
				 l_2 = +37; end
		14682: begin l_1 = +3;
				 l_2 = -37; end
		2937: begin l_1 = -3;
				 l_2 = +37; end
		14674: begin l_1 = -3;
				 l_2 = -37; end
		5886: begin l_1 = +3;
				 l_2 = +38; end
		11741: begin l_1 = +3;
				 l_2 = -38; end
		5878: begin l_1 = -3;
				 l_2 = +38; end
		11733: begin l_1 = -3;
				 l_2 = -38; end
		11768: begin l_1 = +3;
				 l_2 = +39; end
		5859: begin l_1 = +3;
				 l_2 = -39; end
		11760: begin l_1 = -3;
				 l_2 = +39; end
		5851: begin l_1 = -3;
				 l_2 = -39; end
		5913: begin l_1 = +3;
				 l_2 = +40; end
		11714: begin l_1 = +3;
				 l_2 = -40; end
		5905: begin l_1 = -3;
				 l_2 = +40; end
		11706: begin l_1 = -3;
				 l_2 = -40; end
		11822: begin l_1 = +3;
				 l_2 = +41; end
		5805: begin l_1 = +3;
				 l_2 = -41; end
		11814: begin l_1 = -3;
				 l_2 = +41; end
		5797: begin l_1 = -3;
				 l_2 = -41; end
		6021: begin l_1 = +3;
				 l_2 = +42; end
		11606: begin l_1 = +3;
				 l_2 = -42; end
		6013: begin l_1 = -3;
				 l_2 = +42; end
		11598: begin l_1 = -3;
				 l_2 = -42; end
		12038: begin l_1 = +3;
				 l_2 = +43; end
		5589: begin l_1 = +3;
				 l_2 = -43; end
		12030: begin l_1 = -3;
				 l_2 = +43; end
		5581: begin l_1 = -3;
				 l_2 = -43; end
		24: begin l_1 = -4;
				 l_2 = +6; end
		17595: begin l_1 = -4;
				 l_2 = -5; end
		40: begin l_1 = +4;
				 l_2 = +6; end
		17579: begin l_1 = -4;
				 l_2 = -6; end
		72: begin l_1 = +4;
				 l_2 = +7; end
		17563: begin l_1 = +4;
				 l_2 = -7; end
		56: begin l_1 = -4;
				 l_2 = +7; end
		17547: begin l_1 = -4;
				 l_2 = -7; end
		136: begin l_1 = +4;
				 l_2 = +8; end
		17499: begin l_1 = +4;
				 l_2 = -8; end
		120: begin l_1 = -4;
				 l_2 = +8; end
		17483: begin l_1 = -4;
				 l_2 = -8; end
		264: begin l_1 = +4;
				 l_2 = +9; end
		17371: begin l_1 = +4;
				 l_2 = -9; end
		248: begin l_1 = -4;
				 l_2 = +9; end
		17355: begin l_1 = -4;
				 l_2 = -9; end
		520: begin l_1 = +4;
				 l_2 = +10; end
		17115: begin l_1 = +4;
				 l_2 = -10; end
		504: begin l_1 = -4;
				 l_2 = +10; end
		17099: begin l_1 = -4;
				 l_2 = -10; end
		1032: begin l_1 = +4;
				 l_2 = +11; end
		16603: begin l_1 = +4;
				 l_2 = -11; end
		1016: begin l_1 = -4;
				 l_2 = +11; end
		16587: begin l_1 = -4;
				 l_2 = -11; end
		2056: begin l_1 = +4;
				 l_2 = +12; end
		15579: begin l_1 = +4;
				 l_2 = -12; end
		2040: begin l_1 = -4;
				 l_2 = +12; end
		15563: begin l_1 = -4;
				 l_2 = -12; end
		4104: begin l_1 = +4;
				 l_2 = +13; end
		13531: begin l_1 = +4;
				 l_2 = -13; end
		4088: begin l_1 = -4;
				 l_2 = +13; end
		13515: begin l_1 = -4;
				 l_2 = -13; end
		8200: begin l_1 = +4;
				 l_2 = +14; end
		9435: begin l_1 = +4;
				 l_2 = -14; end
		8184: begin l_1 = -4;
				 l_2 = +14; end
		9419: begin l_1 = -4;
				 l_2 = -14; end
		16392: begin l_1 = +4;
				 l_2 = +15; end
		1243: begin l_1 = +4;
				 l_2 = -15; end
		16376: begin l_1 = -4;
				 l_2 = +15; end
		1227: begin l_1 = -4;
				 l_2 = -15; end
		15157: begin l_1 = +4;
				 l_2 = +16; end
		2478: begin l_1 = +4;
				 l_2 = -16; end
		15141: begin l_1 = -4;
				 l_2 = +16; end
		2462: begin l_1 = -4;
				 l_2 = -16; end
		12687: begin l_1 = +4;
				 l_2 = +17; end
		4948: begin l_1 = +4;
				 l_2 = -17; end
		12671: begin l_1 = -4;
				 l_2 = +17; end
		4932: begin l_1 = -4;
				 l_2 = -17; end
		7747: begin l_1 = +4;
				 l_2 = +18; end
		9888: begin l_1 = +4;
				 l_2 = -18; end
		7731: begin l_1 = -4;
				 l_2 = +18; end
		9872: begin l_1 = -4;
				 l_2 = -18; end
		15486: begin l_1 = +4;
				 l_2 = +19; end
		2149: begin l_1 = +4;
				 l_2 = -19; end
		15470: begin l_1 = -4;
				 l_2 = +19; end
		2133: begin l_1 = -4;
				 l_2 = -19; end
		13345: begin l_1 = +4;
				 l_2 = +20; end
		4290: begin l_1 = +4;
				 l_2 = -20; end
		13329: begin l_1 = -4;
				 l_2 = +20; end
		4274: begin l_1 = -4;
				 l_2 = -20; end
		9063: begin l_1 = +4;
				 l_2 = +21; end
		8572: begin l_1 = +4;
				 l_2 = -21; end
		9047: begin l_1 = -4;
				 l_2 = +21; end
		8556: begin l_1 = -4;
				 l_2 = -21; end
		499: begin l_1 = +4;
				 l_2 = +22; end
		17136: begin l_1 = +4;
				 l_2 = -22; end
		483: begin l_1 = -4;
				 l_2 = +22; end
		17120: begin l_1 = -4;
				 l_2 = -22; end
		990: begin l_1 = +4;
				 l_2 = +23; end
		16645: begin l_1 = +4;
				 l_2 = -23; end
		974: begin l_1 = -4;
				 l_2 = +23; end
		16629: begin l_1 = -4;
				 l_2 = -23; end
		1972: begin l_1 = +4;
				 l_2 = +24; end
		15663: begin l_1 = +4;
				 l_2 = -24; end
		1956: begin l_1 = -4;
				 l_2 = +24; end
		15647: begin l_1 = -4;
				 l_2 = -24; end
		3936: begin l_1 = +4;
				 l_2 = +25; end
		13699: begin l_1 = +4;
				 l_2 = -25; end
		3920: begin l_1 = -4;
				 l_2 = +25; end
		13683: begin l_1 = -4;
				 l_2 = -25; end
		7864: begin l_1 = +4;
				 l_2 = +26; end
		9771: begin l_1 = +4;
				 l_2 = -26; end
		7848: begin l_1 = -4;
				 l_2 = +26; end
		9755: begin l_1 = -4;
				 l_2 = -26; end
		15720: begin l_1 = +4;
				 l_2 = +27; end
		1915: begin l_1 = +4;
				 l_2 = -27; end
		15704: begin l_1 = -4;
				 l_2 = +27; end
		1899: begin l_1 = -4;
				 l_2 = -27; end
		13813: begin l_1 = +4;
				 l_2 = +28; end
		3822: begin l_1 = +4;
				 l_2 = -28; end
		13797: begin l_1 = -4;
				 l_2 = +28; end
		3806: begin l_1 = -4;
				 l_2 = -28; end
		9999: begin l_1 = +4;
				 l_2 = +29; end
		7636: begin l_1 = +4;
				 l_2 = -29; end
		9983: begin l_1 = -4;
				 l_2 = +29; end
		7620: begin l_1 = -4;
				 l_2 = -29; end
		2371: begin l_1 = +4;
				 l_2 = +30; end
		15264: begin l_1 = +4;
				 l_2 = -30; end
		2355: begin l_1 = -4;
				 l_2 = +30; end
		15248: begin l_1 = -4;
				 l_2 = -30; end
		4734: begin l_1 = +4;
				 l_2 = +31; end
		12901: begin l_1 = +4;
				 l_2 = -31; end
		4718: begin l_1 = -4;
				 l_2 = +31; end
		12885: begin l_1 = -4;
				 l_2 = -31; end
		9460: begin l_1 = +4;
				 l_2 = +32; end
		8175: begin l_1 = +4;
				 l_2 = -32; end
		9444: begin l_1 = -4;
				 l_2 = +32; end
		8159: begin l_1 = -4;
				 l_2 = -32; end
		1293: begin l_1 = +4;
				 l_2 = +33; end
		16342: begin l_1 = +4;
				 l_2 = -33; end
		1277: begin l_1 = -4;
				 l_2 = +33; end
		16326: begin l_1 = -4;
				 l_2 = -33; end
		2578: begin l_1 = +4;
				 l_2 = +34; end
		15057: begin l_1 = +4;
				 l_2 = -34; end
		2562: begin l_1 = -4;
				 l_2 = +34; end
		15041: begin l_1 = -4;
				 l_2 = -34; end
		5148: begin l_1 = +4;
				 l_2 = +35; end
		12487: begin l_1 = +4;
				 l_2 = -35; end
		5132: begin l_1 = -4;
				 l_2 = +35; end
		12471: begin l_1 = -4;
				 l_2 = -35; end
		10288: begin l_1 = +4;
				 l_2 = +36; end
		7347: begin l_1 = +4;
				 l_2 = -36; end
		10272: begin l_1 = -4;
				 l_2 = +36; end
		7331: begin l_1 = -4;
				 l_2 = -36; end
		2949: begin l_1 = +4;
				 l_2 = +37; end
		14686: begin l_1 = +4;
				 l_2 = -37; end
		2933: begin l_1 = -4;
				 l_2 = +37; end
		14670: begin l_1 = -4;
				 l_2 = -37; end
		5890: begin l_1 = +4;
				 l_2 = +38; end
		11745: begin l_1 = +4;
				 l_2 = -38; end
		5874: begin l_1 = -4;
				 l_2 = +38; end
		11729: begin l_1 = -4;
				 l_2 = -38; end
		11772: begin l_1 = +4;
				 l_2 = +39; end
		5863: begin l_1 = +4;
				 l_2 = -39; end
		11756: begin l_1 = -4;
				 l_2 = +39; end
		5847: begin l_1 = -4;
				 l_2 = -39; end
		5917: begin l_1 = +4;
				 l_2 = +40; end
		11718: begin l_1 = +4;
				 l_2 = -40; end
		5901: begin l_1 = -4;
				 l_2 = +40; end
		11702: begin l_1 = -4;
				 l_2 = -40; end
		11826: begin l_1 = +4;
				 l_2 = +41; end
		5809: begin l_1 = +4;
				 l_2 = -41; end
		11810: begin l_1 = -4;
				 l_2 = +41; end
		5793: begin l_1 = -4;
				 l_2 = -41; end
		6025: begin l_1 = +4;
				 l_2 = +42; end
		11610: begin l_1 = +4;
				 l_2 = -42; end
		6009: begin l_1 = -4;
				 l_2 = +42; end
		11594: begin l_1 = -4;
				 l_2 = -42; end
		12042: begin l_1 = +4;
				 l_2 = +43; end
		5593: begin l_1 = +4;
				 l_2 = -43; end
		12026: begin l_1 = -4;
				 l_2 = +43; end
		5577: begin l_1 = -4;
				 l_2 = -43; end
		48: begin l_1 = -5;
				 l_2 = +7; end
		17571: begin l_1 = -5;
				 l_2 = -6; end
		80: begin l_1 = +5;
				 l_2 = +7; end
		17539: begin l_1 = -5;
				 l_2 = -7; end
		144: begin l_1 = +5;
				 l_2 = +8; end
		17507: begin l_1 = +5;
				 l_2 = -8; end
		112: begin l_1 = -5;
				 l_2 = +8; end
		17475: begin l_1 = -5;
				 l_2 = -8; end
		272: begin l_1 = +5;
				 l_2 = +9; end
		17379: begin l_1 = +5;
				 l_2 = -9; end
		240: begin l_1 = -5;
				 l_2 = +9; end
		17347: begin l_1 = -5;
				 l_2 = -9; end
		528: begin l_1 = +5;
				 l_2 = +10; end
		17123: begin l_1 = +5;
				 l_2 = -10; end
		496: begin l_1 = -5;
				 l_2 = +10; end
		17091: begin l_1 = -5;
				 l_2 = -10; end
		1040: begin l_1 = +5;
				 l_2 = +11; end
		16611: begin l_1 = +5;
				 l_2 = -11; end
		1008: begin l_1 = -5;
				 l_2 = +11; end
		16579: begin l_1 = -5;
				 l_2 = -11; end
		2064: begin l_1 = +5;
				 l_2 = +12; end
		15587: begin l_1 = +5;
				 l_2 = -12; end
		2032: begin l_1 = -5;
				 l_2 = +12; end
		15555: begin l_1 = -5;
				 l_2 = -12; end
		4112: begin l_1 = +5;
				 l_2 = +13; end
		13539: begin l_1 = +5;
				 l_2 = -13; end
		4080: begin l_1 = -5;
				 l_2 = +13; end
		13507: begin l_1 = -5;
				 l_2 = -13; end
		8208: begin l_1 = +5;
				 l_2 = +14; end
		9443: begin l_1 = +5;
				 l_2 = -14; end
		8176: begin l_1 = -5;
				 l_2 = +14; end
		9411: begin l_1 = -5;
				 l_2 = -14; end
		16400: begin l_1 = +5;
				 l_2 = +15; end
		1251: begin l_1 = +5;
				 l_2 = -15; end
		16368: begin l_1 = -5;
				 l_2 = +15; end
		1219: begin l_1 = -5;
				 l_2 = -15; end
		15165: begin l_1 = +5;
				 l_2 = +16; end
		2486: begin l_1 = +5;
				 l_2 = -16; end
		15133: begin l_1 = -5;
				 l_2 = +16; end
		2454: begin l_1 = -5;
				 l_2 = -16; end
		12695: begin l_1 = +5;
				 l_2 = +17; end
		4956: begin l_1 = +5;
				 l_2 = -17; end
		12663: begin l_1 = -5;
				 l_2 = +17; end
		4924: begin l_1 = -5;
				 l_2 = -17; end
		7755: begin l_1 = +5;
				 l_2 = +18; end
		9896: begin l_1 = +5;
				 l_2 = -18; end
		7723: begin l_1 = -5;
				 l_2 = +18; end
		9864: begin l_1 = -5;
				 l_2 = -18; end
		15494: begin l_1 = +5;
				 l_2 = +19; end
		2157: begin l_1 = +5;
				 l_2 = -19; end
		15462: begin l_1 = -5;
				 l_2 = +19; end
		2125: begin l_1 = -5;
				 l_2 = -19; end
		13353: begin l_1 = +5;
				 l_2 = +20; end
		4298: begin l_1 = +5;
				 l_2 = -20; end
		13321: begin l_1 = -5;
				 l_2 = +20; end
		4266: begin l_1 = -5;
				 l_2 = -20; end
		9071: begin l_1 = +5;
				 l_2 = +21; end
		8580: begin l_1 = +5;
				 l_2 = -21; end
		9039: begin l_1 = -5;
				 l_2 = +21; end
		8548: begin l_1 = -5;
				 l_2 = -21; end
		507: begin l_1 = +5;
				 l_2 = +22; end
		17144: begin l_1 = +5;
				 l_2 = -22; end
		475: begin l_1 = -5;
				 l_2 = +22; end
		17112: begin l_1 = -5;
				 l_2 = -22; end
		998: begin l_1 = +5;
				 l_2 = +23; end
		16653: begin l_1 = +5;
				 l_2 = -23; end
		966: begin l_1 = -5;
				 l_2 = +23; end
		16621: begin l_1 = -5;
				 l_2 = -23; end
		1980: begin l_1 = +5;
				 l_2 = +24; end
		15671: begin l_1 = +5;
				 l_2 = -24; end
		1948: begin l_1 = -5;
				 l_2 = +24; end
		15639: begin l_1 = -5;
				 l_2 = -24; end
		3944: begin l_1 = +5;
				 l_2 = +25; end
		13707: begin l_1 = +5;
				 l_2 = -25; end
		3912: begin l_1 = -5;
				 l_2 = +25; end
		13675: begin l_1 = -5;
				 l_2 = -25; end
		7872: begin l_1 = +5;
				 l_2 = +26; end
		9779: begin l_1 = +5;
				 l_2 = -26; end
		7840: begin l_1 = -5;
				 l_2 = +26; end
		9747: begin l_1 = -5;
				 l_2 = -26; end
		15728: begin l_1 = +5;
				 l_2 = +27; end
		1923: begin l_1 = +5;
				 l_2 = -27; end
		15696: begin l_1 = -5;
				 l_2 = +27; end
		1891: begin l_1 = -5;
				 l_2 = -27; end
		13821: begin l_1 = +5;
				 l_2 = +28; end
		3830: begin l_1 = +5;
				 l_2 = -28; end
		13789: begin l_1 = -5;
				 l_2 = +28; end
		3798: begin l_1 = -5;
				 l_2 = -28; end
		10007: begin l_1 = +5;
				 l_2 = +29; end
		7644: begin l_1 = +5;
				 l_2 = -29; end
		9975: begin l_1 = -5;
				 l_2 = +29; end
		7612: begin l_1 = -5;
				 l_2 = -29; end
		2379: begin l_1 = +5;
				 l_2 = +30; end
		15272: begin l_1 = +5;
				 l_2 = -30; end
		2347: begin l_1 = -5;
				 l_2 = +30; end
		15240: begin l_1 = -5;
				 l_2 = -30; end
		4742: begin l_1 = +5;
				 l_2 = +31; end
		12909: begin l_1 = +5;
				 l_2 = -31; end
		4710: begin l_1 = -5;
				 l_2 = +31; end
		12877: begin l_1 = -5;
				 l_2 = -31; end
		9468: begin l_1 = +5;
				 l_2 = +32; end
		8183: begin l_1 = +5;
				 l_2 = -32; end
		9436: begin l_1 = -5;
				 l_2 = +32; end
		8151: begin l_1 = -5;
				 l_2 = -32; end
		1301: begin l_1 = +5;
				 l_2 = +33; end
		16350: begin l_1 = +5;
				 l_2 = -33; end
		1269: begin l_1 = -5;
				 l_2 = +33; end
		16318: begin l_1 = -5;
				 l_2 = -33; end
		2586: begin l_1 = +5;
				 l_2 = +34; end
		15065: begin l_1 = +5;
				 l_2 = -34; end
		2554: begin l_1 = -5;
				 l_2 = +34; end
		15033: begin l_1 = -5;
				 l_2 = -34; end
		5156: begin l_1 = +5;
				 l_2 = +35; end
		12495: begin l_1 = +5;
				 l_2 = -35; end
		5124: begin l_1 = -5;
				 l_2 = +35; end
		12463: begin l_1 = -5;
				 l_2 = -35; end
		10296: begin l_1 = +5;
				 l_2 = +36; end
		7355: begin l_1 = +5;
				 l_2 = -36; end
		10264: begin l_1 = -5;
				 l_2 = +36; end
		7323: begin l_1 = -5;
				 l_2 = -36; end
		2957: begin l_1 = +5;
				 l_2 = +37; end
		14694: begin l_1 = +5;
				 l_2 = -37; end
		2925: begin l_1 = -5;
				 l_2 = +37; end
		14662: begin l_1 = -5;
				 l_2 = -37; end
		5898: begin l_1 = +5;
				 l_2 = +38; end
		11753: begin l_1 = +5;
				 l_2 = -38; end
		5866: begin l_1 = -5;
				 l_2 = +38; end
		11721: begin l_1 = -5;
				 l_2 = -38; end
		11780: begin l_1 = +5;
				 l_2 = +39; end
		5871: begin l_1 = +5;
				 l_2 = -39; end
		11748: begin l_1 = -5;
				 l_2 = +39; end
		5839: begin l_1 = -5;
				 l_2 = -39; end
		5925: begin l_1 = +5;
				 l_2 = +40; end
		11726: begin l_1 = +5;
				 l_2 = -40; end
		5893: begin l_1 = -5;
				 l_2 = +40; end
		11694: begin l_1 = -5;
				 l_2 = -40; end
		11834: begin l_1 = +5;
				 l_2 = +41; end
		5817: begin l_1 = +5;
				 l_2 = -41; end
		11802: begin l_1 = -5;
				 l_2 = +41; end
		5785: begin l_1 = -5;
				 l_2 = -41; end
		6033: begin l_1 = +5;
				 l_2 = +42; end
		11618: begin l_1 = +5;
				 l_2 = -42; end
		6001: begin l_1 = -5;
				 l_2 = +42; end
		11586: begin l_1 = -5;
				 l_2 = -42; end
		12050: begin l_1 = +5;
				 l_2 = +43; end
		5601: begin l_1 = +5;
				 l_2 = -43; end
		12018: begin l_1 = -5;
				 l_2 = +43; end
		5569: begin l_1 = -5;
				 l_2 = -43; end
		96: begin l_1 = -6;
				 l_2 = +8; end
		17523: begin l_1 = -6;
				 l_2 = -7; end
		160: begin l_1 = +6;
				 l_2 = +8; end
		17459: begin l_1 = -6;
				 l_2 = -8; end
		288: begin l_1 = +6;
				 l_2 = +9; end
		17395: begin l_1 = +6;
				 l_2 = -9; end
		224: begin l_1 = -6;
				 l_2 = +9; end
		17331: begin l_1 = -6;
				 l_2 = -9; end
		544: begin l_1 = +6;
				 l_2 = +10; end
		17139: begin l_1 = +6;
				 l_2 = -10; end
		480: begin l_1 = -6;
				 l_2 = +10; end
		17075: begin l_1 = -6;
				 l_2 = -10; end
		1056: begin l_1 = +6;
				 l_2 = +11; end
		16627: begin l_1 = +6;
				 l_2 = -11; end
		992: begin l_1 = -6;
				 l_2 = +11; end
		16563: begin l_1 = -6;
				 l_2 = -11; end
		2080: begin l_1 = +6;
				 l_2 = +12; end
		15603: begin l_1 = +6;
				 l_2 = -12; end
		2016: begin l_1 = -6;
				 l_2 = +12; end
		15539: begin l_1 = -6;
				 l_2 = -12; end
		4128: begin l_1 = +6;
				 l_2 = +13; end
		13555: begin l_1 = +6;
				 l_2 = -13; end
		4064: begin l_1 = -6;
				 l_2 = +13; end
		13491: begin l_1 = -6;
				 l_2 = -13; end
		8224: begin l_1 = +6;
				 l_2 = +14; end
		9459: begin l_1 = +6;
				 l_2 = -14; end
		8160: begin l_1 = -6;
				 l_2 = +14; end
		9395: begin l_1 = -6;
				 l_2 = -14; end
		16416: begin l_1 = +6;
				 l_2 = +15; end
		1267: begin l_1 = +6;
				 l_2 = -15; end
		16352: begin l_1 = -6;
				 l_2 = +15; end
		1203: begin l_1 = -6;
				 l_2 = -15; end
		15181: begin l_1 = +6;
				 l_2 = +16; end
		2502: begin l_1 = +6;
				 l_2 = -16; end
		15117: begin l_1 = -6;
				 l_2 = +16; end
		2438: begin l_1 = -6;
				 l_2 = -16; end
		12711: begin l_1 = +6;
				 l_2 = +17; end
		4972: begin l_1 = +6;
				 l_2 = -17; end
		12647: begin l_1 = -6;
				 l_2 = +17; end
		4908: begin l_1 = -6;
				 l_2 = -17; end
		7771: begin l_1 = +6;
				 l_2 = +18; end
		9912: begin l_1 = +6;
				 l_2 = -18; end
		7707: begin l_1 = -6;
				 l_2 = +18; end
		9848: begin l_1 = -6;
				 l_2 = -18; end
		15510: begin l_1 = +6;
				 l_2 = +19; end
		2173: begin l_1 = +6;
				 l_2 = -19; end
		15446: begin l_1 = -6;
				 l_2 = +19; end
		2109: begin l_1 = -6;
				 l_2 = -19; end
		13369: begin l_1 = +6;
				 l_2 = +20; end
		4314: begin l_1 = +6;
				 l_2 = -20; end
		13305: begin l_1 = -6;
				 l_2 = +20; end
		4250: begin l_1 = -6;
				 l_2 = -20; end
		9087: begin l_1 = +6;
				 l_2 = +21; end
		8596: begin l_1 = +6;
				 l_2 = -21; end
		9023: begin l_1 = -6;
				 l_2 = +21; end
		8532: begin l_1 = -6;
				 l_2 = -21; end
		523: begin l_1 = +6;
				 l_2 = +22; end
		17160: begin l_1 = +6;
				 l_2 = -22; end
		459: begin l_1 = -6;
				 l_2 = +22; end
		17096: begin l_1 = -6;
				 l_2 = -22; end
		1014: begin l_1 = +6;
				 l_2 = +23; end
		16669: begin l_1 = +6;
				 l_2 = -23; end
		950: begin l_1 = -6;
				 l_2 = +23; end
		16605: begin l_1 = -6;
				 l_2 = -23; end
		1996: begin l_1 = +6;
				 l_2 = +24; end
		15687: begin l_1 = +6;
				 l_2 = -24; end
		1932: begin l_1 = -6;
				 l_2 = +24; end
		15623: begin l_1 = -6;
				 l_2 = -24; end
		3960: begin l_1 = +6;
				 l_2 = +25; end
		13723: begin l_1 = +6;
				 l_2 = -25; end
		3896: begin l_1 = -6;
				 l_2 = +25; end
		13659: begin l_1 = -6;
				 l_2 = -25; end
		7888: begin l_1 = +6;
				 l_2 = +26; end
		9795: begin l_1 = +6;
				 l_2 = -26; end
		7824: begin l_1 = -6;
				 l_2 = +26; end
		9731: begin l_1 = -6;
				 l_2 = -26; end
		15744: begin l_1 = +6;
				 l_2 = +27; end
		1939: begin l_1 = +6;
				 l_2 = -27; end
		15680: begin l_1 = -6;
				 l_2 = +27; end
		1875: begin l_1 = -6;
				 l_2 = -27; end
		13837: begin l_1 = +6;
				 l_2 = +28; end
		3846: begin l_1 = +6;
				 l_2 = -28; end
		13773: begin l_1 = -6;
				 l_2 = +28; end
		3782: begin l_1 = -6;
				 l_2 = -28; end
		10023: begin l_1 = +6;
				 l_2 = +29; end
		7660: begin l_1 = +6;
				 l_2 = -29; end
		9959: begin l_1 = -6;
				 l_2 = +29; end
		7596: begin l_1 = -6;
				 l_2 = -29; end
		2395: begin l_1 = +6;
				 l_2 = +30; end
		15288: begin l_1 = +6;
				 l_2 = -30; end
		2331: begin l_1 = -6;
				 l_2 = +30; end
		15224: begin l_1 = -6;
				 l_2 = -30; end
		4758: begin l_1 = +6;
				 l_2 = +31; end
		12925: begin l_1 = +6;
				 l_2 = -31; end
		4694: begin l_1 = -6;
				 l_2 = +31; end
		12861: begin l_1 = -6;
				 l_2 = -31; end
		9484: begin l_1 = +6;
				 l_2 = +32; end
		8199: begin l_1 = +6;
				 l_2 = -32; end
		9420: begin l_1 = -6;
				 l_2 = +32; end
		8135: begin l_1 = -6;
				 l_2 = -32; end
		1317: begin l_1 = +6;
				 l_2 = +33; end
		16366: begin l_1 = +6;
				 l_2 = -33; end
		1253: begin l_1 = -6;
				 l_2 = +33; end
		16302: begin l_1 = -6;
				 l_2 = -33; end
		2602: begin l_1 = +6;
				 l_2 = +34; end
		15081: begin l_1 = +6;
				 l_2 = -34; end
		2538: begin l_1 = -6;
				 l_2 = +34; end
		15017: begin l_1 = -6;
				 l_2 = -34; end
		5172: begin l_1 = +6;
				 l_2 = +35; end
		12511: begin l_1 = +6;
				 l_2 = -35; end
		5108: begin l_1 = -6;
				 l_2 = +35; end
		12447: begin l_1 = -6;
				 l_2 = -35; end
		10312: begin l_1 = +6;
				 l_2 = +36; end
		7371: begin l_1 = +6;
				 l_2 = -36; end
		10248: begin l_1 = -6;
				 l_2 = +36; end
		7307: begin l_1 = -6;
				 l_2 = -36; end
		2973: begin l_1 = +6;
				 l_2 = +37; end
		14710: begin l_1 = +6;
				 l_2 = -37; end
		2909: begin l_1 = -6;
				 l_2 = +37; end
		14646: begin l_1 = -6;
				 l_2 = -37; end
		5914: begin l_1 = +6;
				 l_2 = +38; end
		11769: begin l_1 = +6;
				 l_2 = -38; end
		5850: begin l_1 = -6;
				 l_2 = +38; end
		11705: begin l_1 = -6;
				 l_2 = -38; end
		11796: begin l_1 = +6;
				 l_2 = +39; end
		5887: begin l_1 = +6;
				 l_2 = -39; end
		11732: begin l_1 = -6;
				 l_2 = +39; end
		5823: begin l_1 = -6;
				 l_2 = -39; end
		5941: begin l_1 = +6;
				 l_2 = +40; end
		11742: begin l_1 = +6;
				 l_2 = -40; end
		5877: begin l_1 = -6;
				 l_2 = +40; end
		11678: begin l_1 = -6;
				 l_2 = -40; end
		11850: begin l_1 = +6;
				 l_2 = +41; end
		5833: begin l_1 = +6;
				 l_2 = -41; end
		11786: begin l_1 = -6;
				 l_2 = +41; end
		5769: begin l_1 = -6;
				 l_2 = -41; end
		6049: begin l_1 = +6;
				 l_2 = +42; end
		11634: begin l_1 = +6;
				 l_2 = -42; end
		5985: begin l_1 = -6;
				 l_2 = +42; end
		11570: begin l_1 = -6;
				 l_2 = -42; end
		12066: begin l_1 = +6;
				 l_2 = +43; end
		5617: begin l_1 = +6;
				 l_2 = -43; end
		12002: begin l_1 = -6;
				 l_2 = +43; end
		5553: begin l_1 = -6;
				 l_2 = -43; end
		192: begin l_1 = -7;
				 l_2 = +9; end
		17427: begin l_1 = -7;
				 l_2 = -8; end
		320: begin l_1 = +7;
				 l_2 = +9; end
		17299: begin l_1 = -7;
				 l_2 = -9; end
		576: begin l_1 = +7;
				 l_2 = +10; end
		17171: begin l_1 = +7;
				 l_2 = -10; end
		448: begin l_1 = -7;
				 l_2 = +10; end
		17043: begin l_1 = -7;
				 l_2 = -10; end
		1088: begin l_1 = +7;
				 l_2 = +11; end
		16659: begin l_1 = +7;
				 l_2 = -11; end
		960: begin l_1 = -7;
				 l_2 = +11; end
		16531: begin l_1 = -7;
				 l_2 = -11; end
		2112: begin l_1 = +7;
				 l_2 = +12; end
		15635: begin l_1 = +7;
				 l_2 = -12; end
		1984: begin l_1 = -7;
				 l_2 = +12; end
		15507: begin l_1 = -7;
				 l_2 = -12; end
		4160: begin l_1 = +7;
				 l_2 = +13; end
		13587: begin l_1 = +7;
				 l_2 = -13; end
		4032: begin l_1 = -7;
				 l_2 = +13; end
		13459: begin l_1 = -7;
				 l_2 = -13; end
		8256: begin l_1 = +7;
				 l_2 = +14; end
		9491: begin l_1 = +7;
				 l_2 = -14; end
		8128: begin l_1 = -7;
				 l_2 = +14; end
		9363: begin l_1 = -7;
				 l_2 = -14; end
		16448: begin l_1 = +7;
				 l_2 = +15; end
		1299: begin l_1 = +7;
				 l_2 = -15; end
		16320: begin l_1 = -7;
				 l_2 = +15; end
		1171: begin l_1 = -7;
				 l_2 = -15; end
		15213: begin l_1 = +7;
				 l_2 = +16; end
		2534: begin l_1 = +7;
				 l_2 = -16; end
		15085: begin l_1 = -7;
				 l_2 = +16; end
		2406: begin l_1 = -7;
				 l_2 = -16; end
		12743: begin l_1 = +7;
				 l_2 = +17; end
		5004: begin l_1 = +7;
				 l_2 = -17; end
		12615: begin l_1 = -7;
				 l_2 = +17; end
		4876: begin l_1 = -7;
				 l_2 = -17; end
		7803: begin l_1 = +7;
				 l_2 = +18; end
		9944: begin l_1 = +7;
				 l_2 = -18; end
		7675: begin l_1 = -7;
				 l_2 = +18; end
		9816: begin l_1 = -7;
				 l_2 = -18; end
		15542: begin l_1 = +7;
				 l_2 = +19; end
		2205: begin l_1 = +7;
				 l_2 = -19; end
		15414: begin l_1 = -7;
				 l_2 = +19; end
		2077: begin l_1 = -7;
				 l_2 = -19; end
		13401: begin l_1 = +7;
				 l_2 = +20; end
		4346: begin l_1 = +7;
				 l_2 = -20; end
		13273: begin l_1 = -7;
				 l_2 = +20; end
		4218: begin l_1 = -7;
				 l_2 = -20; end
		9119: begin l_1 = +7;
				 l_2 = +21; end
		8628: begin l_1 = +7;
				 l_2 = -21; end
		8991: begin l_1 = -7;
				 l_2 = +21; end
		8500: begin l_1 = -7;
				 l_2 = -21; end
		555: begin l_1 = +7;
				 l_2 = +22; end
		17192: begin l_1 = +7;
				 l_2 = -22; end
		427: begin l_1 = -7;
				 l_2 = +22; end
		17064: begin l_1 = -7;
				 l_2 = -22; end
		1046: begin l_1 = +7;
				 l_2 = +23; end
		16701: begin l_1 = +7;
				 l_2 = -23; end
		918: begin l_1 = -7;
				 l_2 = +23; end
		16573: begin l_1 = -7;
				 l_2 = -23; end
		2028: begin l_1 = +7;
				 l_2 = +24; end
		15719: begin l_1 = +7;
				 l_2 = -24; end
		1900: begin l_1 = -7;
				 l_2 = +24; end
		15591: begin l_1 = -7;
				 l_2 = -24; end
		3992: begin l_1 = +7;
				 l_2 = +25; end
		13755: begin l_1 = +7;
				 l_2 = -25; end
		3864: begin l_1 = -7;
				 l_2 = +25; end
		13627: begin l_1 = -7;
				 l_2 = -25; end
		7920: begin l_1 = +7;
				 l_2 = +26; end
		9827: begin l_1 = +7;
				 l_2 = -26; end
		7792: begin l_1 = -7;
				 l_2 = +26; end
		9699: begin l_1 = -7;
				 l_2 = -26; end
		15776: begin l_1 = +7;
				 l_2 = +27; end
		1971: begin l_1 = +7;
				 l_2 = -27; end
		15648: begin l_1 = -7;
				 l_2 = +27; end
		1843: begin l_1 = -7;
				 l_2 = -27; end
		13869: begin l_1 = +7;
				 l_2 = +28; end
		3878: begin l_1 = +7;
				 l_2 = -28; end
		13741: begin l_1 = -7;
				 l_2 = +28; end
		3750: begin l_1 = -7;
				 l_2 = -28; end
		10055: begin l_1 = +7;
				 l_2 = +29; end
		7692: begin l_1 = +7;
				 l_2 = -29; end
		9927: begin l_1 = -7;
				 l_2 = +29; end
		7564: begin l_1 = -7;
				 l_2 = -29; end
		2427: begin l_1 = +7;
				 l_2 = +30; end
		15320: begin l_1 = +7;
				 l_2 = -30; end
		2299: begin l_1 = -7;
				 l_2 = +30; end
		15192: begin l_1 = -7;
				 l_2 = -30; end
		4790: begin l_1 = +7;
				 l_2 = +31; end
		12957: begin l_1 = +7;
				 l_2 = -31; end
		4662: begin l_1 = -7;
				 l_2 = +31; end
		12829: begin l_1 = -7;
				 l_2 = -31; end
		9516: begin l_1 = +7;
				 l_2 = +32; end
		8231: begin l_1 = +7;
				 l_2 = -32; end
		9388: begin l_1 = -7;
				 l_2 = +32; end
		8103: begin l_1 = -7;
				 l_2 = -32; end
		1349: begin l_1 = +7;
				 l_2 = +33; end
		16398: begin l_1 = +7;
				 l_2 = -33; end
		1221: begin l_1 = -7;
				 l_2 = +33; end
		16270: begin l_1 = -7;
				 l_2 = -33; end
		2634: begin l_1 = +7;
				 l_2 = +34; end
		15113: begin l_1 = +7;
				 l_2 = -34; end
		2506: begin l_1 = -7;
				 l_2 = +34; end
		14985: begin l_1 = -7;
				 l_2 = -34; end
		5204: begin l_1 = +7;
				 l_2 = +35; end
		12543: begin l_1 = +7;
				 l_2 = -35; end
		5076: begin l_1 = -7;
				 l_2 = +35; end
		12415: begin l_1 = -7;
				 l_2 = -35; end
		10344: begin l_1 = +7;
				 l_2 = +36; end
		7403: begin l_1 = +7;
				 l_2 = -36; end
		10216: begin l_1 = -7;
				 l_2 = +36; end
		7275: begin l_1 = -7;
				 l_2 = -36; end
		3005: begin l_1 = +7;
				 l_2 = +37; end
		14742: begin l_1 = +7;
				 l_2 = -37; end
		2877: begin l_1 = -7;
				 l_2 = +37; end
		14614: begin l_1 = -7;
				 l_2 = -37; end
		5946: begin l_1 = +7;
				 l_2 = +38; end
		11801: begin l_1 = +7;
				 l_2 = -38; end
		5818: begin l_1 = -7;
				 l_2 = +38; end
		11673: begin l_1 = -7;
				 l_2 = -38; end
		11828: begin l_1 = +7;
				 l_2 = +39; end
		5919: begin l_1 = +7;
				 l_2 = -39; end
		11700: begin l_1 = -7;
				 l_2 = +39; end
		5791: begin l_1 = -7;
				 l_2 = -39; end
		5973: begin l_1 = +7;
				 l_2 = +40; end
		11774: begin l_1 = +7;
				 l_2 = -40; end
		5845: begin l_1 = -7;
				 l_2 = +40; end
		11646: begin l_1 = -7;
				 l_2 = -40; end
		11882: begin l_1 = +7;
				 l_2 = +41; end
		5865: begin l_1 = +7;
				 l_2 = -41; end
		11754: begin l_1 = -7;
				 l_2 = +41; end
		5737: begin l_1 = -7;
				 l_2 = -41; end
		6081: begin l_1 = +7;
				 l_2 = +42; end
		11666: begin l_1 = +7;
				 l_2 = -42; end
		5953: begin l_1 = -7;
				 l_2 = +42; end
		11538: begin l_1 = -7;
				 l_2 = -42; end
		12098: begin l_1 = +7;
				 l_2 = +43; end
		5649: begin l_1 = +7;
				 l_2 = -43; end
		11970: begin l_1 = -7;
				 l_2 = +43; end
		5521: begin l_1 = -7;
				 l_2 = -43; end
		384: begin l_1 = -8;
				 l_2 = +10; end
		17235: begin l_1 = -8;
				 l_2 = -9; end
		640: begin l_1 = +8;
				 l_2 = +10; end
		16979: begin l_1 = -8;
				 l_2 = -10; end
		1152: begin l_1 = +8;
				 l_2 = +11; end
		16723: begin l_1 = +8;
				 l_2 = -11; end
		896: begin l_1 = -8;
				 l_2 = +11; end
		16467: begin l_1 = -8;
				 l_2 = -11; end
		2176: begin l_1 = +8;
				 l_2 = +12; end
		15699: begin l_1 = +8;
				 l_2 = -12; end
		1920: begin l_1 = -8;
				 l_2 = +12; end
		15443: begin l_1 = -8;
				 l_2 = -12; end
		4224: begin l_1 = +8;
				 l_2 = +13; end
		13651: begin l_1 = +8;
				 l_2 = -13; end
		3968: begin l_1 = -8;
				 l_2 = +13; end
		13395: begin l_1 = -8;
				 l_2 = -13; end
		8320: begin l_1 = +8;
				 l_2 = +14; end
		9555: begin l_1 = +8;
				 l_2 = -14; end
		8064: begin l_1 = -8;
				 l_2 = +14; end
		9299: begin l_1 = -8;
				 l_2 = -14; end
		16512: begin l_1 = +8;
				 l_2 = +15; end
		1363: begin l_1 = +8;
				 l_2 = -15; end
		16256: begin l_1 = -8;
				 l_2 = +15; end
		1107: begin l_1 = -8;
				 l_2 = -15; end
		15277: begin l_1 = +8;
				 l_2 = +16; end
		2598: begin l_1 = +8;
				 l_2 = -16; end
		15021: begin l_1 = -8;
				 l_2 = +16; end
		2342: begin l_1 = -8;
				 l_2 = -16; end
		12807: begin l_1 = +8;
				 l_2 = +17; end
		5068: begin l_1 = +8;
				 l_2 = -17; end
		12551: begin l_1 = -8;
				 l_2 = +17; end
		4812: begin l_1 = -8;
				 l_2 = -17; end
		7867: begin l_1 = +8;
				 l_2 = +18; end
		10008: begin l_1 = +8;
				 l_2 = -18; end
		7611: begin l_1 = -8;
				 l_2 = +18; end
		9752: begin l_1 = -8;
				 l_2 = -18; end
		15606: begin l_1 = +8;
				 l_2 = +19; end
		2269: begin l_1 = +8;
				 l_2 = -19; end
		15350: begin l_1 = -8;
				 l_2 = +19; end
		2013: begin l_1 = -8;
				 l_2 = -19; end
		13465: begin l_1 = +8;
				 l_2 = +20; end
		4410: begin l_1 = +8;
				 l_2 = -20; end
		13209: begin l_1 = -8;
				 l_2 = +20; end
		4154: begin l_1 = -8;
				 l_2 = -20; end
		9183: begin l_1 = +8;
				 l_2 = +21; end
		8692: begin l_1 = +8;
				 l_2 = -21; end
		8927: begin l_1 = -8;
				 l_2 = +21; end
		8436: begin l_1 = -8;
				 l_2 = -21; end
		619: begin l_1 = +8;
				 l_2 = +22; end
		17256: begin l_1 = +8;
				 l_2 = -22; end
		363: begin l_1 = -8;
				 l_2 = +22; end
		17000: begin l_1 = -8;
				 l_2 = -22; end
		1110: begin l_1 = +8;
				 l_2 = +23; end
		16765: begin l_1 = +8;
				 l_2 = -23; end
		854: begin l_1 = -8;
				 l_2 = +23; end
		16509: begin l_1 = -8;
				 l_2 = -23; end
		2092: begin l_1 = +8;
				 l_2 = +24; end
		15783: begin l_1 = +8;
				 l_2 = -24; end
		1836: begin l_1 = -8;
				 l_2 = +24; end
		15527: begin l_1 = -8;
				 l_2 = -24; end
		4056: begin l_1 = +8;
				 l_2 = +25; end
		13819: begin l_1 = +8;
				 l_2 = -25; end
		3800: begin l_1 = -8;
				 l_2 = +25; end
		13563: begin l_1 = -8;
				 l_2 = -25; end
		7984: begin l_1 = +8;
				 l_2 = +26; end
		9891: begin l_1 = +8;
				 l_2 = -26; end
		7728: begin l_1 = -8;
				 l_2 = +26; end
		9635: begin l_1 = -8;
				 l_2 = -26; end
		15840: begin l_1 = +8;
				 l_2 = +27; end
		2035: begin l_1 = +8;
				 l_2 = -27; end
		15584: begin l_1 = -8;
				 l_2 = +27; end
		1779: begin l_1 = -8;
				 l_2 = -27; end
		13933: begin l_1 = +8;
				 l_2 = +28; end
		3942: begin l_1 = +8;
				 l_2 = -28; end
		13677: begin l_1 = -8;
				 l_2 = +28; end
		3686: begin l_1 = -8;
				 l_2 = -28; end
		10119: begin l_1 = +8;
				 l_2 = +29; end
		7756: begin l_1 = +8;
				 l_2 = -29; end
		9863: begin l_1 = -8;
				 l_2 = +29; end
		7500: begin l_1 = -8;
				 l_2 = -29; end
		2491: begin l_1 = +8;
				 l_2 = +30; end
		15384: begin l_1 = +8;
				 l_2 = -30; end
		2235: begin l_1 = -8;
				 l_2 = +30; end
		15128: begin l_1 = -8;
				 l_2 = -30; end
		4854: begin l_1 = +8;
				 l_2 = +31; end
		13021: begin l_1 = +8;
				 l_2 = -31; end
		4598: begin l_1 = -8;
				 l_2 = +31; end
		12765: begin l_1 = -8;
				 l_2 = -31; end
		9580: begin l_1 = +8;
				 l_2 = +32; end
		8295: begin l_1 = +8;
				 l_2 = -32; end
		9324: begin l_1 = -8;
				 l_2 = +32; end
		8039: begin l_1 = -8;
				 l_2 = -32; end
		1413: begin l_1 = +8;
				 l_2 = +33; end
		16462: begin l_1 = +8;
				 l_2 = -33; end
		1157: begin l_1 = -8;
				 l_2 = +33; end
		16206: begin l_1 = -8;
				 l_2 = -33; end
		2698: begin l_1 = +8;
				 l_2 = +34; end
		15177: begin l_1 = +8;
				 l_2 = -34; end
		2442: begin l_1 = -8;
				 l_2 = +34; end
		14921: begin l_1 = -8;
				 l_2 = -34; end
		5268: begin l_1 = +8;
				 l_2 = +35; end
		12607: begin l_1 = +8;
				 l_2 = -35; end
		5012: begin l_1 = -8;
				 l_2 = +35; end
		12351: begin l_1 = -8;
				 l_2 = -35; end
		10408: begin l_1 = +8;
				 l_2 = +36; end
		7467: begin l_1 = +8;
				 l_2 = -36; end
		10152: begin l_1 = -8;
				 l_2 = +36; end
		7211: begin l_1 = -8;
				 l_2 = -36; end
		3069: begin l_1 = +8;
				 l_2 = +37; end
		14806: begin l_1 = +8;
				 l_2 = -37; end
		2813: begin l_1 = -8;
				 l_2 = +37; end
		14550: begin l_1 = -8;
				 l_2 = -37; end
		6010: begin l_1 = +8;
				 l_2 = +38; end
		11865: begin l_1 = +8;
				 l_2 = -38; end
		5754: begin l_1 = -8;
				 l_2 = +38; end
		11609: begin l_1 = -8;
				 l_2 = -38; end
		11892: begin l_1 = +8;
				 l_2 = +39; end
		5983: begin l_1 = +8;
				 l_2 = -39; end
		11636: begin l_1 = -8;
				 l_2 = +39; end
		5727: begin l_1 = -8;
				 l_2 = -39; end
		6037: begin l_1 = +8;
				 l_2 = +40; end
		11838: begin l_1 = +8;
				 l_2 = -40; end
		5781: begin l_1 = -8;
				 l_2 = +40; end
		11582: begin l_1 = -8;
				 l_2 = -40; end
		11946: begin l_1 = +8;
				 l_2 = +41; end
		5929: begin l_1 = +8;
				 l_2 = -41; end
		11690: begin l_1 = -8;
				 l_2 = +41; end
		5673: begin l_1 = -8;
				 l_2 = -41; end
		6145: begin l_1 = +8;
				 l_2 = +42; end
		11730: begin l_1 = +8;
				 l_2 = -42; end
		5889: begin l_1 = -8;
				 l_2 = +42; end
		11474: begin l_1 = -8;
				 l_2 = -42; end
		12162: begin l_1 = +8;
				 l_2 = +43; end
		5713: begin l_1 = +8;
				 l_2 = -43; end
		11906: begin l_1 = -8;
				 l_2 = +43; end
		5457: begin l_1 = -8;
				 l_2 = -43; end
		768: begin l_1 = -9;
				 l_2 = +11; end
		16851: begin l_1 = -9;
				 l_2 = -10; end
		1280: begin l_1 = +9;
				 l_2 = +11; end
		16339: begin l_1 = -9;
				 l_2 = -11; end
		2304: begin l_1 = +9;
				 l_2 = +12; end
		15827: begin l_1 = +9;
				 l_2 = -12; end
		1792: begin l_1 = -9;
				 l_2 = +12; end
		15315: begin l_1 = -9;
				 l_2 = -12; end
		4352: begin l_1 = +9;
				 l_2 = +13; end
		13779: begin l_1 = +9;
				 l_2 = -13; end
		3840: begin l_1 = -9;
				 l_2 = +13; end
		13267: begin l_1 = -9;
				 l_2 = -13; end
		8448: begin l_1 = +9;
				 l_2 = +14; end
		9683: begin l_1 = +9;
				 l_2 = -14; end
		7936: begin l_1 = -9;
				 l_2 = +14; end
		9171: begin l_1 = -9;
				 l_2 = -14; end
		16640: begin l_1 = +9;
				 l_2 = +15; end
		1491: begin l_1 = +9;
				 l_2 = -15; end
		16128: begin l_1 = -9;
				 l_2 = +15; end
		979: begin l_1 = -9;
				 l_2 = -15; end
		15405: begin l_1 = +9;
				 l_2 = +16; end
		2726: begin l_1 = +9;
				 l_2 = -16; end
		14893: begin l_1 = -9;
				 l_2 = +16; end
		2214: begin l_1 = -9;
				 l_2 = -16; end
		12935: begin l_1 = +9;
				 l_2 = +17; end
		5196: begin l_1 = +9;
				 l_2 = -17; end
		12423: begin l_1 = -9;
				 l_2 = +17; end
		4684: begin l_1 = -9;
				 l_2 = -17; end
		7995: begin l_1 = +9;
				 l_2 = +18; end
		10136: begin l_1 = +9;
				 l_2 = -18; end
		7483: begin l_1 = -9;
				 l_2 = +18; end
		9624: begin l_1 = -9;
				 l_2 = -18; end
		15734: begin l_1 = +9;
				 l_2 = +19; end
		2397: begin l_1 = +9;
				 l_2 = -19; end
		15222: begin l_1 = -9;
				 l_2 = +19; end
		1885: begin l_1 = -9;
				 l_2 = -19; end
		13593: begin l_1 = +9;
				 l_2 = +20; end
		4538: begin l_1 = +9;
				 l_2 = -20; end
		13081: begin l_1 = -9;
				 l_2 = +20; end
		4026: begin l_1 = -9;
				 l_2 = -20; end
		9311: begin l_1 = +9;
				 l_2 = +21; end
		8820: begin l_1 = +9;
				 l_2 = -21; end
		8799: begin l_1 = -9;
				 l_2 = +21; end
		8308: begin l_1 = -9;
				 l_2 = -21; end
		747: begin l_1 = +9;
				 l_2 = +22; end
		17384: begin l_1 = +9;
				 l_2 = -22; end
		235: begin l_1 = -9;
				 l_2 = +22; end
		16872: begin l_1 = -9;
				 l_2 = -22; end
		1238: begin l_1 = +9;
				 l_2 = +23; end
		16893: begin l_1 = +9;
				 l_2 = -23; end
		726: begin l_1 = -9;
				 l_2 = +23; end
		16381: begin l_1 = -9;
				 l_2 = -23; end
		2220: begin l_1 = +9;
				 l_2 = +24; end
		15911: begin l_1 = +9;
				 l_2 = -24; end
		1708: begin l_1 = -9;
				 l_2 = +24; end
		15399: begin l_1 = -9;
				 l_2 = -24; end
		4184: begin l_1 = +9;
				 l_2 = +25; end
		13947: begin l_1 = +9;
				 l_2 = -25; end
		3672: begin l_1 = -9;
				 l_2 = +25; end
		13435: begin l_1 = -9;
				 l_2 = -25; end
		8112: begin l_1 = +9;
				 l_2 = +26; end
		10019: begin l_1 = +9;
				 l_2 = -26; end
		7600: begin l_1 = -9;
				 l_2 = +26; end
		9507: begin l_1 = -9;
				 l_2 = -26; end
		15968: begin l_1 = +9;
				 l_2 = +27; end
		2163: begin l_1 = +9;
				 l_2 = -27; end
		15456: begin l_1 = -9;
				 l_2 = +27; end
		1651: begin l_1 = -9;
				 l_2 = -27; end
		14061: begin l_1 = +9;
				 l_2 = +28; end
		4070: begin l_1 = +9;
				 l_2 = -28; end
		13549: begin l_1 = -9;
				 l_2 = +28; end
		3558: begin l_1 = -9;
				 l_2 = -28; end
		10247: begin l_1 = +9;
				 l_2 = +29; end
		7884: begin l_1 = +9;
				 l_2 = -29; end
		9735: begin l_1 = -9;
				 l_2 = +29; end
		7372: begin l_1 = -9;
				 l_2 = -29; end
		2619: begin l_1 = +9;
				 l_2 = +30; end
		15512: begin l_1 = +9;
				 l_2 = -30; end
		2107: begin l_1 = -9;
				 l_2 = +30; end
		15000: begin l_1 = -9;
				 l_2 = -30; end
		4982: begin l_1 = +9;
				 l_2 = +31; end
		13149: begin l_1 = +9;
				 l_2 = -31; end
		4470: begin l_1 = -9;
				 l_2 = +31; end
		12637: begin l_1 = -9;
				 l_2 = -31; end
		9708: begin l_1 = +9;
				 l_2 = +32; end
		8423: begin l_1 = +9;
				 l_2 = -32; end
		9196: begin l_1 = -9;
				 l_2 = +32; end
		7911: begin l_1 = -9;
				 l_2 = -32; end
		1541: begin l_1 = +9;
				 l_2 = +33; end
		16590: begin l_1 = +9;
				 l_2 = -33; end
		1029: begin l_1 = -9;
				 l_2 = +33; end
		16078: begin l_1 = -9;
				 l_2 = -33; end
		2826: begin l_1 = +9;
				 l_2 = +34; end
		15305: begin l_1 = +9;
				 l_2 = -34; end
		2314: begin l_1 = -9;
				 l_2 = +34; end
		14793: begin l_1 = -9;
				 l_2 = -34; end
		5396: begin l_1 = +9;
				 l_2 = +35; end
		12735: begin l_1 = +9;
				 l_2 = -35; end
		4884: begin l_1 = -9;
				 l_2 = +35; end
		12223: begin l_1 = -9;
				 l_2 = -35; end
		10536: begin l_1 = +9;
				 l_2 = +36; end
		7595: begin l_1 = +9;
				 l_2 = -36; end
		10024: begin l_1 = -9;
				 l_2 = +36; end
		7083: begin l_1 = -9;
				 l_2 = -36; end
		3197: begin l_1 = +9;
				 l_2 = +37; end
		14934: begin l_1 = +9;
				 l_2 = -37; end
		2685: begin l_1 = -9;
				 l_2 = +37; end
		14422: begin l_1 = -9;
				 l_2 = -37; end
		6138: begin l_1 = +9;
				 l_2 = +38; end
		11993: begin l_1 = +9;
				 l_2 = -38; end
		5626: begin l_1 = -9;
				 l_2 = +38; end
		11481: begin l_1 = -9;
				 l_2 = -38; end
		12020: begin l_1 = +9;
				 l_2 = +39; end
		6111: begin l_1 = +9;
				 l_2 = -39; end
		11508: begin l_1 = -9;
				 l_2 = +39; end
		5599: begin l_1 = -9;
				 l_2 = -39; end
		6165: begin l_1 = +9;
				 l_2 = +40; end
		11966: begin l_1 = +9;
				 l_2 = -40; end
		5653: begin l_1 = -9;
				 l_2 = +40; end
		11454: begin l_1 = -9;
				 l_2 = -40; end
		12074: begin l_1 = +9;
				 l_2 = +41; end
		6057: begin l_1 = +9;
				 l_2 = -41; end
		11562: begin l_1 = -9;
				 l_2 = +41; end
		5545: begin l_1 = -9;
				 l_2 = -41; end
		6273: begin l_1 = +9;
				 l_2 = +42; end
		11858: begin l_1 = +9;
				 l_2 = -42; end
		5761: begin l_1 = -9;
				 l_2 = +42; end
		11346: begin l_1 = -9;
				 l_2 = -42; end
		12290: begin l_1 = +9;
				 l_2 = +43; end
		5841: begin l_1 = +9;
				 l_2 = -43; end
		11778: begin l_1 = -9;
				 l_2 = +43; end
		5329: begin l_1 = -9;
				 l_2 = -43; end
		1536: begin l_1 = -10;
				 l_2 = +12; end
		16083: begin l_1 = -10;
				 l_2 = -11; end
		2560: begin l_1 = +10;
				 l_2 = +12; end
		15059: begin l_1 = -10;
				 l_2 = -12; end
		4608: begin l_1 = +10;
				 l_2 = +13; end
		14035: begin l_1 = +10;
				 l_2 = -13; end
		3584: begin l_1 = -10;
				 l_2 = +13; end
		13011: begin l_1 = -10;
				 l_2 = -13; end
		8704: begin l_1 = +10;
				 l_2 = +14; end
		9939: begin l_1 = +10;
				 l_2 = -14; end
		7680: begin l_1 = -10;
				 l_2 = +14; end
		8915: begin l_1 = -10;
				 l_2 = -14; end
		16896: begin l_1 = +10;
				 l_2 = +15; end
		1747: begin l_1 = +10;
				 l_2 = -15; end
		15872: begin l_1 = -10;
				 l_2 = +15; end
		723: begin l_1 = -10;
				 l_2 = -15; end
		15661: begin l_1 = +10;
				 l_2 = +16; end
		2982: begin l_1 = +10;
				 l_2 = -16; end
		14637: begin l_1 = -10;
				 l_2 = +16; end
		1958: begin l_1 = -10;
				 l_2 = -16; end
		13191: begin l_1 = +10;
				 l_2 = +17; end
		5452: begin l_1 = +10;
				 l_2 = -17; end
		12167: begin l_1 = -10;
				 l_2 = +17; end
		4428: begin l_1 = -10;
				 l_2 = -17; end
		8251: begin l_1 = +10;
				 l_2 = +18; end
		10392: begin l_1 = +10;
				 l_2 = -18; end
		7227: begin l_1 = -10;
				 l_2 = +18; end
		9368: begin l_1 = -10;
				 l_2 = -18; end
		15990: begin l_1 = +10;
				 l_2 = +19; end
		2653: begin l_1 = +10;
				 l_2 = -19; end
		14966: begin l_1 = -10;
				 l_2 = +19; end
		1629: begin l_1 = -10;
				 l_2 = -19; end
		13849: begin l_1 = +10;
				 l_2 = +20; end
		4794: begin l_1 = +10;
				 l_2 = -20; end
		12825: begin l_1 = -10;
				 l_2 = +20; end
		3770: begin l_1 = -10;
				 l_2 = -20; end
		9567: begin l_1 = +10;
				 l_2 = +21; end
		9076: begin l_1 = +10;
				 l_2 = -21; end
		8543: begin l_1 = -10;
				 l_2 = +21; end
		8052: begin l_1 = -10;
				 l_2 = -21; end
		1003: begin l_1 = +10;
				 l_2 = +22; end
		21: begin l_1 = +10;
				 l_2 = -22; end
		17598: begin l_1 = -10;
				 l_2 = +22; end
		16616: begin l_1 = -10;
				 l_2 = -22; end
		1494: begin l_1 = +10;
				 l_2 = +23; end
		17149: begin l_1 = +10;
				 l_2 = -23; end
		470: begin l_1 = -10;
				 l_2 = +23; end
		16125: begin l_1 = -10;
				 l_2 = -23; end
		2476: begin l_1 = +10;
				 l_2 = +24; end
		16167: begin l_1 = +10;
				 l_2 = -24; end
		1452: begin l_1 = -10;
				 l_2 = +24; end
		15143: begin l_1 = -10;
				 l_2 = -24; end
		4440: begin l_1 = +10;
				 l_2 = +25; end
		14203: begin l_1 = +10;
				 l_2 = -25; end
		3416: begin l_1 = -10;
				 l_2 = +25; end
		13179: begin l_1 = -10;
				 l_2 = -25; end
		8368: begin l_1 = +10;
				 l_2 = +26; end
		10275: begin l_1 = +10;
				 l_2 = -26; end
		7344: begin l_1 = -10;
				 l_2 = +26; end
		9251: begin l_1 = -10;
				 l_2 = -26; end
		16224: begin l_1 = +10;
				 l_2 = +27; end
		2419: begin l_1 = +10;
				 l_2 = -27; end
		15200: begin l_1 = -10;
				 l_2 = +27; end
		1395: begin l_1 = -10;
				 l_2 = -27; end
		14317: begin l_1 = +10;
				 l_2 = +28; end
		4326: begin l_1 = +10;
				 l_2 = -28; end
		13293: begin l_1 = -10;
				 l_2 = +28; end
		3302: begin l_1 = -10;
				 l_2 = -28; end
		10503: begin l_1 = +10;
				 l_2 = +29; end
		8140: begin l_1 = +10;
				 l_2 = -29; end
		9479: begin l_1 = -10;
				 l_2 = +29; end
		7116: begin l_1 = -10;
				 l_2 = -29; end
		2875: begin l_1 = +10;
				 l_2 = +30; end
		15768: begin l_1 = +10;
				 l_2 = -30; end
		1851: begin l_1 = -10;
				 l_2 = +30; end
		14744: begin l_1 = -10;
				 l_2 = -30; end
		5238: begin l_1 = +10;
				 l_2 = +31; end
		13405: begin l_1 = +10;
				 l_2 = -31; end
		4214: begin l_1 = -10;
				 l_2 = +31; end
		12381: begin l_1 = -10;
				 l_2 = -31; end
		9964: begin l_1 = +10;
				 l_2 = +32; end
		8679: begin l_1 = +10;
				 l_2 = -32; end
		8940: begin l_1 = -10;
				 l_2 = +32; end
		7655: begin l_1 = -10;
				 l_2 = -32; end
		1797: begin l_1 = +10;
				 l_2 = +33; end
		16846: begin l_1 = +10;
				 l_2 = -33; end
		773: begin l_1 = -10;
				 l_2 = +33; end
		15822: begin l_1 = -10;
				 l_2 = -33; end
		3082: begin l_1 = +10;
				 l_2 = +34; end
		15561: begin l_1 = +10;
				 l_2 = -34; end
		2058: begin l_1 = -10;
				 l_2 = +34; end
		14537: begin l_1 = -10;
				 l_2 = -34; end
		5652: begin l_1 = +10;
				 l_2 = +35; end
		12991: begin l_1 = +10;
				 l_2 = -35; end
		4628: begin l_1 = -10;
				 l_2 = +35; end
		11967: begin l_1 = -10;
				 l_2 = -35; end
		10792: begin l_1 = +10;
				 l_2 = +36; end
		7851: begin l_1 = +10;
				 l_2 = -36; end
		9768: begin l_1 = -10;
				 l_2 = +36; end
		6827: begin l_1 = -10;
				 l_2 = -36; end
		3453: begin l_1 = +10;
				 l_2 = +37; end
		15190: begin l_1 = +10;
				 l_2 = -37; end
		2429: begin l_1 = -10;
				 l_2 = +37; end
		14166: begin l_1 = -10;
				 l_2 = -37; end
		6394: begin l_1 = +10;
				 l_2 = +38; end
		12249: begin l_1 = +10;
				 l_2 = -38; end
		5370: begin l_1 = -10;
				 l_2 = +38; end
		11225: begin l_1 = -10;
				 l_2 = -38; end
		12276: begin l_1 = +10;
				 l_2 = +39; end
		6367: begin l_1 = +10;
				 l_2 = -39; end
		11252: begin l_1 = -10;
				 l_2 = +39; end
		5343: begin l_1 = -10;
				 l_2 = -39; end
		6421: begin l_1 = +10;
				 l_2 = +40; end
		12222: begin l_1 = +10;
				 l_2 = -40; end
		5397: begin l_1 = -10;
				 l_2 = +40; end
		11198: begin l_1 = -10;
				 l_2 = -40; end
		12330: begin l_1 = +10;
				 l_2 = +41; end
		6313: begin l_1 = +10;
				 l_2 = -41; end
		11306: begin l_1 = -10;
				 l_2 = +41; end
		5289: begin l_1 = -10;
				 l_2 = -41; end
		6529: begin l_1 = +10;
				 l_2 = +42; end
		12114: begin l_1 = +10;
				 l_2 = -42; end
		5505: begin l_1 = -10;
				 l_2 = +42; end
		11090: begin l_1 = -10;
				 l_2 = -42; end
		12546: begin l_1 = +10;
				 l_2 = +43; end
		6097: begin l_1 = +10;
				 l_2 = -43; end
		11522: begin l_1 = -10;
				 l_2 = +43; end
		5073: begin l_1 = -10;
				 l_2 = -43; end
		3072: begin l_1 = -11;
				 l_2 = +13; end
		14547: begin l_1 = -11;
				 l_2 = -12; end
		5120: begin l_1 = +11;
				 l_2 = +13; end
		12499: begin l_1 = -11;
				 l_2 = -13; end
		9216: begin l_1 = +11;
				 l_2 = +14; end
		10451: begin l_1 = +11;
				 l_2 = -14; end
		7168: begin l_1 = -11;
				 l_2 = +14; end
		8403: begin l_1 = -11;
				 l_2 = -14; end
		17408: begin l_1 = +11;
				 l_2 = +15; end
		2259: begin l_1 = +11;
				 l_2 = -15; end
		15360: begin l_1 = -11;
				 l_2 = +15; end
		211: begin l_1 = -11;
				 l_2 = -15; end
		16173: begin l_1 = +11;
				 l_2 = +16; end
		3494: begin l_1 = +11;
				 l_2 = -16; end
		14125: begin l_1 = -11;
				 l_2 = +16; end
		1446: begin l_1 = -11;
				 l_2 = -16; end
		13703: begin l_1 = +11;
				 l_2 = +17; end
		5964: begin l_1 = +11;
				 l_2 = -17; end
		11655: begin l_1 = -11;
				 l_2 = +17; end
		3916: begin l_1 = -11;
				 l_2 = -17; end
		8763: begin l_1 = +11;
				 l_2 = +18; end
		10904: begin l_1 = +11;
				 l_2 = -18; end
		6715: begin l_1 = -11;
				 l_2 = +18; end
		8856: begin l_1 = -11;
				 l_2 = -18; end
		16502: begin l_1 = +11;
				 l_2 = +19; end
		3165: begin l_1 = +11;
				 l_2 = -19; end
		14454: begin l_1 = -11;
				 l_2 = +19; end
		1117: begin l_1 = -11;
				 l_2 = -19; end
		14361: begin l_1 = +11;
				 l_2 = +20; end
		5306: begin l_1 = +11;
				 l_2 = -20; end
		12313: begin l_1 = -11;
				 l_2 = +20; end
		3258: begin l_1 = -11;
				 l_2 = -20; end
		10079: begin l_1 = +11;
				 l_2 = +21; end
		9588: begin l_1 = +11;
				 l_2 = -21; end
		8031: begin l_1 = -11;
				 l_2 = +21; end
		7540: begin l_1 = -11;
				 l_2 = -21; end
		1515: begin l_1 = +11;
				 l_2 = +22; end
		533: begin l_1 = +11;
				 l_2 = -22; end
		17086: begin l_1 = -11;
				 l_2 = +22; end
		16104: begin l_1 = -11;
				 l_2 = -22; end
		2006: begin l_1 = +11;
				 l_2 = +23; end
		42: begin l_1 = +11;
				 l_2 = -23; end
		17577: begin l_1 = -11;
				 l_2 = +23; end
		15613: begin l_1 = -11;
				 l_2 = -23; end
		2988: begin l_1 = +11;
				 l_2 = +24; end
		16679: begin l_1 = +11;
				 l_2 = -24; end
		940: begin l_1 = -11;
				 l_2 = +24; end
		14631: begin l_1 = -11;
				 l_2 = -24; end
		4952: begin l_1 = +11;
				 l_2 = +25; end
		14715: begin l_1 = +11;
				 l_2 = -25; end
		2904: begin l_1 = -11;
				 l_2 = +25; end
		12667: begin l_1 = -11;
				 l_2 = -25; end
		8880: begin l_1 = +11;
				 l_2 = +26; end
		10787: begin l_1 = +11;
				 l_2 = -26; end
		6832: begin l_1 = -11;
				 l_2 = +26; end
		8739: begin l_1 = -11;
				 l_2 = -26; end
		16736: begin l_1 = +11;
				 l_2 = +27; end
		2931: begin l_1 = +11;
				 l_2 = -27; end
		14688: begin l_1 = -11;
				 l_2 = +27; end
		883: begin l_1 = -11;
				 l_2 = -27; end
		14829: begin l_1 = +11;
				 l_2 = +28; end
		4838: begin l_1 = +11;
				 l_2 = -28; end
		12781: begin l_1 = -11;
				 l_2 = +28; end
		2790: begin l_1 = -11;
				 l_2 = -28; end
		11015: begin l_1 = +11;
				 l_2 = +29; end
		8652: begin l_1 = +11;
				 l_2 = -29; end
		8967: begin l_1 = -11;
				 l_2 = +29; end
		6604: begin l_1 = -11;
				 l_2 = -29; end
		3387: begin l_1 = +11;
				 l_2 = +30; end
		16280: begin l_1 = +11;
				 l_2 = -30; end
		1339: begin l_1 = -11;
				 l_2 = +30; end
		14232: begin l_1 = -11;
				 l_2 = -30; end
		5750: begin l_1 = +11;
				 l_2 = +31; end
		13917: begin l_1 = +11;
				 l_2 = -31; end
		3702: begin l_1 = -11;
				 l_2 = +31; end
		11869: begin l_1 = -11;
				 l_2 = -31; end
		10476: begin l_1 = +11;
				 l_2 = +32; end
		9191: begin l_1 = +11;
				 l_2 = -32; end
		8428: begin l_1 = -11;
				 l_2 = +32; end
		7143: begin l_1 = -11;
				 l_2 = -32; end
		2309: begin l_1 = +11;
				 l_2 = +33; end
		17358: begin l_1 = +11;
				 l_2 = -33; end
		261: begin l_1 = -11;
				 l_2 = +33; end
		15310: begin l_1 = -11;
				 l_2 = -33; end
		3594: begin l_1 = +11;
				 l_2 = +34; end
		16073: begin l_1 = +11;
				 l_2 = -34; end
		1546: begin l_1 = -11;
				 l_2 = +34; end
		14025: begin l_1 = -11;
				 l_2 = -34; end
		6164: begin l_1 = +11;
				 l_2 = +35; end
		13503: begin l_1 = +11;
				 l_2 = -35; end
		4116: begin l_1 = -11;
				 l_2 = +35; end
		11455: begin l_1 = -11;
				 l_2 = -35; end
		11304: begin l_1 = +11;
				 l_2 = +36; end
		8363: begin l_1 = +11;
				 l_2 = -36; end
		9256: begin l_1 = -11;
				 l_2 = +36; end
		6315: begin l_1 = -11;
				 l_2 = -36; end
		3965: begin l_1 = +11;
				 l_2 = +37; end
		15702: begin l_1 = +11;
				 l_2 = -37; end
		1917: begin l_1 = -11;
				 l_2 = +37; end
		13654: begin l_1 = -11;
				 l_2 = -37; end
		6906: begin l_1 = +11;
				 l_2 = +38; end
		12761: begin l_1 = +11;
				 l_2 = -38; end
		4858: begin l_1 = -11;
				 l_2 = +38; end
		10713: begin l_1 = -11;
				 l_2 = -38; end
		12788: begin l_1 = +11;
				 l_2 = +39; end
		6879: begin l_1 = +11;
				 l_2 = -39; end
		10740: begin l_1 = -11;
				 l_2 = +39; end
		4831: begin l_1 = -11;
				 l_2 = -39; end
		6933: begin l_1 = +11;
				 l_2 = +40; end
		12734: begin l_1 = +11;
				 l_2 = -40; end
		4885: begin l_1 = -11;
				 l_2 = +40; end
		10686: begin l_1 = -11;
				 l_2 = -40; end
		12842: begin l_1 = +11;
				 l_2 = +41; end
		6825: begin l_1 = +11;
				 l_2 = -41; end
		10794: begin l_1 = -11;
				 l_2 = +41; end
		4777: begin l_1 = -11;
				 l_2 = -41; end
		7041: begin l_1 = +11;
				 l_2 = +42; end
		12626: begin l_1 = +11;
				 l_2 = -42; end
		4993: begin l_1 = -11;
				 l_2 = +42; end
		10578: begin l_1 = -11;
				 l_2 = -42; end
		13058: begin l_1 = +11;
				 l_2 = +43; end
		6609: begin l_1 = +11;
				 l_2 = -43; end
		11010: begin l_1 = -11;
				 l_2 = +43; end
		4561: begin l_1 = -11;
				 l_2 = -43; end
		6144: begin l_1 = -12;
				 l_2 = +14; end
		11475: begin l_1 = -12;
				 l_2 = -13; end
		10240: begin l_1 = +12;
				 l_2 = +14; end
		7379: begin l_1 = -12;
				 l_2 = -14; end
		813: begin l_1 = +12;
				 l_2 = +15; end
		3283: begin l_1 = +12;
				 l_2 = -15; end
		14336: begin l_1 = -12;
				 l_2 = +15; end
		16806: begin l_1 = -12;
				 l_2 = -15; end
		17197: begin l_1 = +12;
				 l_2 = +16; end
		4518: begin l_1 = +12;
				 l_2 = -16; end
		13101: begin l_1 = -12;
				 l_2 = +16; end
		422: begin l_1 = -12;
				 l_2 = -16; end
		14727: begin l_1 = +12;
				 l_2 = +17; end
		6988: begin l_1 = +12;
				 l_2 = -17; end
		10631: begin l_1 = -12;
				 l_2 = +17; end
		2892: begin l_1 = -12;
				 l_2 = -17; end
		9787: begin l_1 = +12;
				 l_2 = +18; end
		11928: begin l_1 = +12;
				 l_2 = -18; end
		5691: begin l_1 = -12;
				 l_2 = +18; end
		7832: begin l_1 = -12;
				 l_2 = -18; end
		17526: begin l_1 = +12;
				 l_2 = +19; end
		4189: begin l_1 = +12;
				 l_2 = -19; end
		13430: begin l_1 = -12;
				 l_2 = +19; end
		93: begin l_1 = -12;
				 l_2 = -19; end
		15385: begin l_1 = +12;
				 l_2 = +20; end
		6330: begin l_1 = +12;
				 l_2 = -20; end
		11289: begin l_1 = -12;
				 l_2 = +20; end
		2234: begin l_1 = -12;
				 l_2 = -20; end
		11103: begin l_1 = +12;
				 l_2 = +21; end
		10612: begin l_1 = +12;
				 l_2 = -21; end
		7007: begin l_1 = -12;
				 l_2 = +21; end
		6516: begin l_1 = -12;
				 l_2 = -21; end
		2539: begin l_1 = +12;
				 l_2 = +22; end
		1557: begin l_1 = +12;
				 l_2 = -22; end
		16062: begin l_1 = -12;
				 l_2 = +22; end
		15080: begin l_1 = -12;
				 l_2 = -22; end
		3030: begin l_1 = +12;
				 l_2 = +23; end
		1066: begin l_1 = +12;
				 l_2 = -23; end
		16553: begin l_1 = -12;
				 l_2 = +23; end
		14589: begin l_1 = -12;
				 l_2 = -23; end
		4012: begin l_1 = +12;
				 l_2 = +24; end
		84: begin l_1 = +12;
				 l_2 = -24; end
		17535: begin l_1 = -12;
				 l_2 = +24; end
		13607: begin l_1 = -12;
				 l_2 = -24; end
		5976: begin l_1 = +12;
				 l_2 = +25; end
		15739: begin l_1 = +12;
				 l_2 = -25; end
		1880: begin l_1 = -12;
				 l_2 = +25; end
		11643: begin l_1 = -12;
				 l_2 = -25; end
		9904: begin l_1 = +12;
				 l_2 = +26; end
		11811: begin l_1 = +12;
				 l_2 = -26; end
		5808: begin l_1 = -12;
				 l_2 = +26; end
		7715: begin l_1 = -12;
				 l_2 = -26; end
		141: begin l_1 = +12;
				 l_2 = +27; end
		3955: begin l_1 = +12;
				 l_2 = -27; end
		13664: begin l_1 = -12;
				 l_2 = +27; end
		17478: begin l_1 = -12;
				 l_2 = -27; end
		15853: begin l_1 = +12;
				 l_2 = +28; end
		5862: begin l_1 = +12;
				 l_2 = -28; end
		11757: begin l_1 = -12;
				 l_2 = +28; end
		1766: begin l_1 = -12;
				 l_2 = -28; end
		12039: begin l_1 = +12;
				 l_2 = +29; end
		9676: begin l_1 = +12;
				 l_2 = -29; end
		7943: begin l_1 = -12;
				 l_2 = +29; end
		5580: begin l_1 = -12;
				 l_2 = -29; end
		4411: begin l_1 = +12;
				 l_2 = +30; end
		17304: begin l_1 = +12;
				 l_2 = -30; end
		315: begin l_1 = -12;
				 l_2 = +30; end
		13208: begin l_1 = -12;
				 l_2 = -30; end
		6774: begin l_1 = +12;
				 l_2 = +31; end
		14941: begin l_1 = +12;
				 l_2 = -31; end
		2678: begin l_1 = -12;
				 l_2 = +31; end
		10845: begin l_1 = -12;
				 l_2 = -31; end
		11500: begin l_1 = +12;
				 l_2 = +32; end
		10215: begin l_1 = +12;
				 l_2 = -32; end
		7404: begin l_1 = -12;
				 l_2 = +32; end
		6119: begin l_1 = -12;
				 l_2 = -32; end
		3333: begin l_1 = +12;
				 l_2 = +33; end
		763: begin l_1 = +12;
				 l_2 = -33; end
		16856: begin l_1 = -12;
				 l_2 = +33; end
		14286: begin l_1 = -12;
				 l_2 = -33; end
		4618: begin l_1 = +12;
				 l_2 = +34; end
		17097: begin l_1 = +12;
				 l_2 = -34; end
		522: begin l_1 = -12;
				 l_2 = +34; end
		13001: begin l_1 = -12;
				 l_2 = -34; end
		7188: begin l_1 = +12;
				 l_2 = +35; end
		14527: begin l_1 = +12;
				 l_2 = -35; end
		3092: begin l_1 = -12;
				 l_2 = +35; end
		10431: begin l_1 = -12;
				 l_2 = -35; end
		12328: begin l_1 = +12;
				 l_2 = +36; end
		9387: begin l_1 = +12;
				 l_2 = -36; end
		8232: begin l_1 = -12;
				 l_2 = +36; end
		5291: begin l_1 = -12;
				 l_2 = -36; end
		4989: begin l_1 = +12;
				 l_2 = +37; end
		16726: begin l_1 = +12;
				 l_2 = -37; end
		893: begin l_1 = -12;
				 l_2 = +37; end
		12630: begin l_1 = -12;
				 l_2 = -37; end
		7930: begin l_1 = +12;
				 l_2 = +38; end
		13785: begin l_1 = +12;
				 l_2 = -38; end
		3834: begin l_1 = -12;
				 l_2 = +38; end
		9689: begin l_1 = -12;
				 l_2 = -38; end
		13812: begin l_1 = +12;
				 l_2 = +39; end
		7903: begin l_1 = +12;
				 l_2 = -39; end
		9716: begin l_1 = -12;
				 l_2 = +39; end
		3807: begin l_1 = -12;
				 l_2 = -39; end
		7957: begin l_1 = +12;
				 l_2 = +40; end
		13758: begin l_1 = +12;
				 l_2 = -40; end
		3861: begin l_1 = -12;
				 l_2 = +40; end
		9662: begin l_1 = -12;
				 l_2 = -40; end
		13866: begin l_1 = +12;
				 l_2 = +41; end
		7849: begin l_1 = +12;
				 l_2 = -41; end
		9770: begin l_1 = -12;
				 l_2 = +41; end
		3753: begin l_1 = -12;
				 l_2 = -41; end
		8065: begin l_1 = +12;
				 l_2 = +42; end
		13650: begin l_1 = +12;
				 l_2 = -42; end
		3969: begin l_1 = -12;
				 l_2 = +42; end
		9554: begin l_1 = -12;
				 l_2 = -42; end
		14082: begin l_1 = +12;
				 l_2 = +43; end
		7633: begin l_1 = +12;
				 l_2 = -43; end
		9986: begin l_1 = -12;
				 l_2 = +43; end
		3537: begin l_1 = -12;
				 l_2 = -43; end
		12288: begin l_1 = -13;
				 l_2 = +15; end
		5331: begin l_1 = -13;
				 l_2 = -14; end
		2861: begin l_1 = +13;
				 l_2 = +15; end
		14758: begin l_1 = -13;
				 l_2 = -15; end
		1626: begin l_1 = +13;
				 l_2 = +16; end
		6566: begin l_1 = +13;
				 l_2 = -16; end
		11053: begin l_1 = -13;
				 l_2 = +16; end
		15993: begin l_1 = -13;
				 l_2 = -16; end
		16775: begin l_1 = +13;
				 l_2 = +17; end
		9036: begin l_1 = +13;
				 l_2 = -17; end
		8583: begin l_1 = -13;
				 l_2 = +17; end
		844: begin l_1 = -13;
				 l_2 = -17; end
		11835: begin l_1 = +13;
				 l_2 = +18; end
		13976: begin l_1 = +13;
				 l_2 = -18; end
		3643: begin l_1 = -13;
				 l_2 = +18; end
		5784: begin l_1 = -13;
				 l_2 = -18; end
		1955: begin l_1 = +13;
				 l_2 = +19; end
		6237: begin l_1 = +13;
				 l_2 = -19; end
		11382: begin l_1 = -13;
				 l_2 = +19; end
		15664: begin l_1 = -13;
				 l_2 = -19; end
		17433: begin l_1 = +13;
				 l_2 = +20; end
		8378: begin l_1 = +13;
				 l_2 = -20; end
		9241: begin l_1 = -13;
				 l_2 = +20; end
		186: begin l_1 = -13;
				 l_2 = -20; end
		13151: begin l_1 = +13;
				 l_2 = +21; end
		12660: begin l_1 = +13;
				 l_2 = -21; end
		4959: begin l_1 = -13;
				 l_2 = +21; end
		4468: begin l_1 = -13;
				 l_2 = -21; end
		4587: begin l_1 = +13;
				 l_2 = +22; end
		3605: begin l_1 = +13;
				 l_2 = -22; end
		14014: begin l_1 = -13;
				 l_2 = +22; end
		13032: begin l_1 = -13;
				 l_2 = -22; end
		5078: begin l_1 = +13;
				 l_2 = +23; end
		3114: begin l_1 = +13;
				 l_2 = -23; end
		14505: begin l_1 = -13;
				 l_2 = +23; end
		12541: begin l_1 = -13;
				 l_2 = -23; end
		6060: begin l_1 = +13;
				 l_2 = +24; end
		2132: begin l_1 = +13;
				 l_2 = -24; end
		15487: begin l_1 = -13;
				 l_2 = +24; end
		11559: begin l_1 = -13;
				 l_2 = -24; end
		8024: begin l_1 = +13;
				 l_2 = +25; end
		168: begin l_1 = +13;
				 l_2 = -25; end
		17451: begin l_1 = -13;
				 l_2 = +25; end
		9595: begin l_1 = -13;
				 l_2 = -25; end
		11952: begin l_1 = +13;
				 l_2 = +26; end
		13859: begin l_1 = +13;
				 l_2 = -26; end
		3760: begin l_1 = -13;
				 l_2 = +26; end
		5667: begin l_1 = -13;
				 l_2 = -26; end
		2189: begin l_1 = +13;
				 l_2 = +27; end
		6003: begin l_1 = +13;
				 l_2 = -27; end
		11616: begin l_1 = -13;
				 l_2 = +27; end
		15430: begin l_1 = -13;
				 l_2 = -27; end
		282: begin l_1 = +13;
				 l_2 = +28; end
		7910: begin l_1 = +13;
				 l_2 = -28; end
		9709: begin l_1 = -13;
				 l_2 = +28; end
		17337: begin l_1 = -13;
				 l_2 = -28; end
		14087: begin l_1 = +13;
				 l_2 = +29; end
		11724: begin l_1 = +13;
				 l_2 = -29; end
		5895: begin l_1 = -13;
				 l_2 = +29; end
		3532: begin l_1 = -13;
				 l_2 = -29; end
		6459: begin l_1 = +13;
				 l_2 = +30; end
		1733: begin l_1 = +13;
				 l_2 = -30; end
		15886: begin l_1 = -13;
				 l_2 = +30; end
		11160: begin l_1 = -13;
				 l_2 = -30; end
		8822: begin l_1 = +13;
				 l_2 = +31; end
		16989: begin l_1 = +13;
				 l_2 = -31; end
		630: begin l_1 = -13;
				 l_2 = +31; end
		8797: begin l_1 = -13;
				 l_2 = -31; end
		13548: begin l_1 = +13;
				 l_2 = +32; end
		12263: begin l_1 = +13;
				 l_2 = -32; end
		5356: begin l_1 = -13;
				 l_2 = +32; end
		4071: begin l_1 = -13;
				 l_2 = -32; end
		5381: begin l_1 = +13;
				 l_2 = +33; end
		2811: begin l_1 = +13;
				 l_2 = -33; end
		14808: begin l_1 = -13;
				 l_2 = +33; end
		12238: begin l_1 = -13;
				 l_2 = -33; end
		6666: begin l_1 = +13;
				 l_2 = +34; end
		1526: begin l_1 = +13;
				 l_2 = -34; end
		16093: begin l_1 = -13;
				 l_2 = +34; end
		10953: begin l_1 = -13;
				 l_2 = -34; end
		9236: begin l_1 = +13;
				 l_2 = +35; end
		16575: begin l_1 = +13;
				 l_2 = -35; end
		1044: begin l_1 = -13;
				 l_2 = +35; end
		8383: begin l_1 = -13;
				 l_2 = -35; end
		14376: begin l_1 = +13;
				 l_2 = +36; end
		11435: begin l_1 = +13;
				 l_2 = -36; end
		6184: begin l_1 = -13;
				 l_2 = +36; end
		3243: begin l_1 = -13;
				 l_2 = -36; end
		7037: begin l_1 = +13;
				 l_2 = +37; end
		1155: begin l_1 = +13;
				 l_2 = -37; end
		16464: begin l_1 = -13;
				 l_2 = +37; end
		10582: begin l_1 = -13;
				 l_2 = -37; end
		9978: begin l_1 = +13;
				 l_2 = +38; end
		15833: begin l_1 = +13;
				 l_2 = -38; end
		1786: begin l_1 = -13;
				 l_2 = +38; end
		7641: begin l_1 = -13;
				 l_2 = -38; end
		15860: begin l_1 = +13;
				 l_2 = +39; end
		9951: begin l_1 = +13;
				 l_2 = -39; end
		7668: begin l_1 = -13;
				 l_2 = +39; end
		1759: begin l_1 = -13;
				 l_2 = -39; end
		10005: begin l_1 = +13;
				 l_2 = +40; end
		15806: begin l_1 = +13;
				 l_2 = -40; end
		1813: begin l_1 = -13;
				 l_2 = +40; end
		7614: begin l_1 = -13;
				 l_2 = -40; end
		15914: begin l_1 = +13;
				 l_2 = +41; end
		9897: begin l_1 = +13;
				 l_2 = -41; end
		7722: begin l_1 = -13;
				 l_2 = +41; end
		1705: begin l_1 = -13;
				 l_2 = -41; end
		10113: begin l_1 = +13;
				 l_2 = +42; end
		15698: begin l_1 = +13;
				 l_2 = -42; end
		1921: begin l_1 = -13;
				 l_2 = +42; end
		7506: begin l_1 = -13;
				 l_2 = -42; end
		16130: begin l_1 = +13;
				 l_2 = +43; end
		9681: begin l_1 = +13;
				 l_2 = -43; end
		7938: begin l_1 = -13;
				 l_2 = +43; end
		1489: begin l_1 = -13;
				 l_2 = -43; end
		6957: begin l_1 = -14;
				 l_2 = +16; end
		10662: begin l_1 = -14;
				 l_2 = -15; end
		5722: begin l_1 = +14;
				 l_2 = +16; end
		11897: begin l_1 = -14;
				 l_2 = -16; end
		3252: begin l_1 = +14;
				 l_2 = +17; end
		13132: begin l_1 = +14;
				 l_2 = -17; end
		4487: begin l_1 = -14;
				 l_2 = +17; end
		14367: begin l_1 = -14;
				 l_2 = -17; end
		15931: begin l_1 = +14;
				 l_2 = +18; end
		453: begin l_1 = +14;
				 l_2 = -18; end
		17166: begin l_1 = -14;
				 l_2 = +18; end
		1688: begin l_1 = -14;
				 l_2 = -18; end
		6051: begin l_1 = +14;
				 l_2 = +19; end
		10333: begin l_1 = +14;
				 l_2 = -19; end
		7286: begin l_1 = -14;
				 l_2 = +19; end
		11568: begin l_1 = -14;
				 l_2 = -19; end
		3910: begin l_1 = +14;
				 l_2 = +20; end
		12474: begin l_1 = +14;
				 l_2 = -20; end
		5145: begin l_1 = -14;
				 l_2 = +20; end
		13709: begin l_1 = -14;
				 l_2 = -20; end
		17247: begin l_1 = +14;
				 l_2 = +21; end
		16756: begin l_1 = +14;
				 l_2 = -21; end
		863: begin l_1 = -14;
				 l_2 = +21; end
		372: begin l_1 = -14;
				 l_2 = -21; end
		8683: begin l_1 = +14;
				 l_2 = +22; end
		7701: begin l_1 = +14;
				 l_2 = -22; end
		9918: begin l_1 = -14;
				 l_2 = +22; end
		8936: begin l_1 = -14;
				 l_2 = -22; end
		9174: begin l_1 = +14;
				 l_2 = +23; end
		7210: begin l_1 = +14;
				 l_2 = -23; end
		10409: begin l_1 = -14;
				 l_2 = +23; end
		8445: begin l_1 = -14;
				 l_2 = -23; end
		10156: begin l_1 = +14;
				 l_2 = +24; end
		6228: begin l_1 = +14;
				 l_2 = -24; end
		11391: begin l_1 = -14;
				 l_2 = +24; end
		7463: begin l_1 = -14;
				 l_2 = -24; end
		12120: begin l_1 = +14;
				 l_2 = +25; end
		4264: begin l_1 = +14;
				 l_2 = -25; end
		13355: begin l_1 = -14;
				 l_2 = +25; end
		5499: begin l_1 = -14;
				 l_2 = -25; end
		16048: begin l_1 = +14;
				 l_2 = +26; end
		336: begin l_1 = +14;
				 l_2 = -26; end
		17283: begin l_1 = -14;
				 l_2 = +26; end
		1571: begin l_1 = -14;
				 l_2 = -26; end
		6285: begin l_1 = +14;
				 l_2 = +27; end
		10099: begin l_1 = +14;
				 l_2 = -27; end
		7520: begin l_1 = -14;
				 l_2 = +27; end
		11334: begin l_1 = -14;
				 l_2 = -27; end
		4378: begin l_1 = +14;
				 l_2 = +28; end
		12006: begin l_1 = +14;
				 l_2 = -28; end
		5613: begin l_1 = -14;
				 l_2 = +28; end
		13241: begin l_1 = -14;
				 l_2 = -28; end
		564: begin l_1 = +14;
				 l_2 = +29; end
		15820: begin l_1 = +14;
				 l_2 = -29; end
		1799: begin l_1 = -14;
				 l_2 = +29; end
		17055: begin l_1 = -14;
				 l_2 = -29; end
		10555: begin l_1 = +14;
				 l_2 = +30; end
		5829: begin l_1 = +14;
				 l_2 = -30; end
		11790: begin l_1 = -14;
				 l_2 = +30; end
		7064: begin l_1 = -14;
				 l_2 = -30; end
		12918: begin l_1 = +14;
				 l_2 = +31; end
		3466: begin l_1 = +14;
				 l_2 = -31; end
		14153: begin l_1 = -14;
				 l_2 = +31; end
		4701: begin l_1 = -14;
				 l_2 = -31; end
		25: begin l_1 = +14;
				 l_2 = +32; end
		16359: begin l_1 = +14;
				 l_2 = -32; end
		1260: begin l_1 = -14;
				 l_2 = +32; end
		17594: begin l_1 = -14;
				 l_2 = -32; end
		9477: begin l_1 = +14;
				 l_2 = +33; end
		6907: begin l_1 = +14;
				 l_2 = -33; end
		10712: begin l_1 = -14;
				 l_2 = +33; end
		8142: begin l_1 = -14;
				 l_2 = -33; end
		10762: begin l_1 = +14;
				 l_2 = +34; end
		5622: begin l_1 = +14;
				 l_2 = -34; end
		11997: begin l_1 = -14;
				 l_2 = +34; end
		6857: begin l_1 = -14;
				 l_2 = -34; end
		13332: begin l_1 = +14;
				 l_2 = +35; end
		3052: begin l_1 = +14;
				 l_2 = -35; end
		14567: begin l_1 = -14;
				 l_2 = +35; end
		4287: begin l_1 = -14;
				 l_2 = -35; end
		853: begin l_1 = +14;
				 l_2 = +36; end
		15531: begin l_1 = +14;
				 l_2 = -36; end
		2088: begin l_1 = -14;
				 l_2 = +36; end
		16766: begin l_1 = -14;
				 l_2 = -36; end
		11133: begin l_1 = +14;
				 l_2 = +37; end
		5251: begin l_1 = +14;
				 l_2 = -37; end
		12368: begin l_1 = -14;
				 l_2 = +37; end
		6486: begin l_1 = -14;
				 l_2 = -37; end
		14074: begin l_1 = +14;
				 l_2 = +38; end
		2310: begin l_1 = +14;
				 l_2 = -38; end
		15309: begin l_1 = -14;
				 l_2 = +38; end
		3545: begin l_1 = -14;
				 l_2 = -38; end
		2337: begin l_1 = +14;
				 l_2 = +39; end
		14047: begin l_1 = +14;
				 l_2 = -39; end
		3572: begin l_1 = -14;
				 l_2 = +39; end
		15282: begin l_1 = -14;
				 l_2 = -39; end
		14101: begin l_1 = +14;
				 l_2 = +40; end
		2283: begin l_1 = +14;
				 l_2 = -40; end
		15336: begin l_1 = -14;
				 l_2 = +40; end
		3518: begin l_1 = -14;
				 l_2 = -40; end
		2391: begin l_1 = +14;
				 l_2 = +41; end
		13993: begin l_1 = +14;
				 l_2 = -41; end
		3626: begin l_1 = -14;
				 l_2 = +41; end
		15228: begin l_1 = -14;
				 l_2 = -41; end
		14209: begin l_1 = +14;
				 l_2 = +42; end
		2175: begin l_1 = +14;
				 l_2 = -42; end
		15444: begin l_1 = -14;
				 l_2 = +42; end
		3410: begin l_1 = -14;
				 l_2 = -42; end
		2607: begin l_1 = +14;
				 l_2 = +43; end
		13777: begin l_1 = +14;
				 l_2 = -43; end
		3842: begin l_1 = -14;
				 l_2 = +43; end
		15012: begin l_1 = -14;
				 l_2 = -43; end
		13914: begin l_1 = -15;
				 l_2 = +17; end
		3705: begin l_1 = -15;
				 l_2 = -16; end
		11444: begin l_1 = +15;
				 l_2 = +17; end
		6175: begin l_1 = -15;
				 l_2 = -17; end
		6504: begin l_1 = +15;
				 l_2 = +18; end
		8645: begin l_1 = +15;
				 l_2 = -18; end
		8974: begin l_1 = -15;
				 l_2 = +18; end
		11115: begin l_1 = -15;
				 l_2 = -18; end
		14243: begin l_1 = +15;
				 l_2 = +19; end
		906: begin l_1 = +15;
				 l_2 = -19; end
		16713: begin l_1 = -15;
				 l_2 = +19; end
		3376: begin l_1 = -15;
				 l_2 = -19; end
		12102: begin l_1 = +15;
				 l_2 = +20; end
		3047: begin l_1 = +15;
				 l_2 = -20; end
		14572: begin l_1 = -15;
				 l_2 = +20; end
		5517: begin l_1 = -15;
				 l_2 = -20; end
		7820: begin l_1 = +15;
				 l_2 = +21; end
		7329: begin l_1 = +15;
				 l_2 = -21; end
		10290: begin l_1 = -15;
				 l_2 = +21; end
		9799: begin l_1 = -15;
				 l_2 = -21; end
		16875: begin l_1 = +15;
				 l_2 = +22; end
		15893: begin l_1 = +15;
				 l_2 = -22; end
		1726: begin l_1 = -15;
				 l_2 = +22; end
		744: begin l_1 = -15;
				 l_2 = -22; end
		17366: begin l_1 = +15;
				 l_2 = +23; end
		15402: begin l_1 = +15;
				 l_2 = -23; end
		2217: begin l_1 = -15;
				 l_2 = +23; end
		253: begin l_1 = -15;
				 l_2 = -23; end
		729: begin l_1 = +15;
				 l_2 = +24; end
		14420: begin l_1 = +15;
				 l_2 = -24; end
		3199: begin l_1 = -15;
				 l_2 = +24; end
		16890: begin l_1 = -15;
				 l_2 = -24; end
		2693: begin l_1 = +15;
				 l_2 = +25; end
		12456: begin l_1 = +15;
				 l_2 = -25; end
		5163: begin l_1 = -15;
				 l_2 = +25; end
		14926: begin l_1 = -15;
				 l_2 = -25; end
		6621: begin l_1 = +15;
				 l_2 = +26; end
		8528: begin l_1 = +15;
				 l_2 = -26; end
		9091: begin l_1 = -15;
				 l_2 = +26; end
		10998: begin l_1 = -15;
				 l_2 = -26; end
		14477: begin l_1 = +15;
				 l_2 = +27; end
		672: begin l_1 = +15;
				 l_2 = -27; end
		16947: begin l_1 = -15;
				 l_2 = +27; end
		3142: begin l_1 = -15;
				 l_2 = -27; end
		12570: begin l_1 = +15;
				 l_2 = +28; end
		2579: begin l_1 = +15;
				 l_2 = -28; end
		15040: begin l_1 = -15;
				 l_2 = +28; end
		5049: begin l_1 = -15;
				 l_2 = -28; end
		8756: begin l_1 = +15;
				 l_2 = +29; end
		6393: begin l_1 = +15;
				 l_2 = -29; end
		11226: begin l_1 = -15;
				 l_2 = +29; end
		8863: begin l_1 = -15;
				 l_2 = -29; end
		1128: begin l_1 = +15;
				 l_2 = +30; end
		14021: begin l_1 = +15;
				 l_2 = -30; end
		3598: begin l_1 = -15;
				 l_2 = +30; end
		16491: begin l_1 = -15;
				 l_2 = -30; end
		3491: begin l_1 = +15;
				 l_2 = +31; end
		11658: begin l_1 = +15;
				 l_2 = -31; end
		5961: begin l_1 = -15;
				 l_2 = +31; end
		14128: begin l_1 = -15;
				 l_2 = -31; end
		8217: begin l_1 = +15;
				 l_2 = +32; end
		6932: begin l_1 = +15;
				 l_2 = -32; end
		10687: begin l_1 = -15;
				 l_2 = +32; end
		9402: begin l_1 = -15;
				 l_2 = -32; end
		50: begin l_1 = +15;
				 l_2 = +33; end
		15099: begin l_1 = +15;
				 l_2 = -33; end
		2520: begin l_1 = -15;
				 l_2 = +33; end
		17569: begin l_1 = -15;
				 l_2 = -33; end
		1335: begin l_1 = +15;
				 l_2 = +34; end
		13814: begin l_1 = +15;
				 l_2 = -34; end
		3805: begin l_1 = -15;
				 l_2 = +34; end
		16284: begin l_1 = -15;
				 l_2 = -34; end
		3905: begin l_1 = +15;
				 l_2 = +35; end
		11244: begin l_1 = +15;
				 l_2 = -35; end
		6375: begin l_1 = -15;
				 l_2 = +35; end
		13714: begin l_1 = -15;
				 l_2 = -35; end
		9045: begin l_1 = +15;
				 l_2 = +36; end
		6104: begin l_1 = +15;
				 l_2 = -36; end
		11515: begin l_1 = -15;
				 l_2 = +36; end
		8574: begin l_1 = -15;
				 l_2 = -36; end
		1706: begin l_1 = +15;
				 l_2 = +37; end
		13443: begin l_1 = +15;
				 l_2 = -37; end
		4176: begin l_1 = -15;
				 l_2 = +37; end
		15913: begin l_1 = -15;
				 l_2 = -37; end
		4647: begin l_1 = +15;
				 l_2 = +38; end
		10502: begin l_1 = +15;
				 l_2 = -38; end
		7117: begin l_1 = -15;
				 l_2 = +38; end
		12972: begin l_1 = -15;
				 l_2 = -38; end
		10529: begin l_1 = +15;
				 l_2 = +39; end
		4620: begin l_1 = +15;
				 l_2 = -39; end
		12999: begin l_1 = -15;
				 l_2 = +39; end
		7090: begin l_1 = -15;
				 l_2 = -39; end
		4674: begin l_1 = +15;
				 l_2 = +40; end
		10475: begin l_1 = +15;
				 l_2 = -40; end
		7144: begin l_1 = -15;
				 l_2 = +40; end
		12945: begin l_1 = -15;
				 l_2 = -40; end
		10583: begin l_1 = +15;
				 l_2 = +41; end
		4566: begin l_1 = +15;
				 l_2 = -41; end
		13053: begin l_1 = -15;
				 l_2 = +41; end
		7036: begin l_1 = -15;
				 l_2 = -41; end
		4782: begin l_1 = +15;
				 l_2 = +42; end
		10367: begin l_1 = +15;
				 l_2 = -42; end
		7252: begin l_1 = -15;
				 l_2 = +42; end
		12837: begin l_1 = -15;
				 l_2 = -42; end
		10799: begin l_1 = +15;
				 l_2 = +43; end
		4350: begin l_1 = +15;
				 l_2 = -43; end
		13269: begin l_1 = -15;
				 l_2 = +43; end
		6820: begin l_1 = -15;
				 l_2 = -43; end
		10209: begin l_1 = -16;
				 l_2 = +18; end
		7410: begin l_1 = -16;
				 l_2 = -17; end
		5269: begin l_1 = +16;
				 l_2 = +18; end
		12350: begin l_1 = -16;
				 l_2 = -18; end
		13008: begin l_1 = +16;
				 l_2 = +19; end
		17290: begin l_1 = +16;
				 l_2 = -19; end
		329: begin l_1 = -16;
				 l_2 = +19; end
		4611: begin l_1 = -16;
				 l_2 = -19; end
		10867: begin l_1 = +16;
				 l_2 = +20; end
		1812: begin l_1 = +16;
				 l_2 = -20; end
		15807: begin l_1 = -16;
				 l_2 = +20; end
		6752: begin l_1 = -16;
				 l_2 = -20; end
		6585: begin l_1 = +16;
				 l_2 = +21; end
		6094: begin l_1 = +16;
				 l_2 = -21; end
		11525: begin l_1 = -16;
				 l_2 = +21; end
		11034: begin l_1 = -16;
				 l_2 = -21; end
		15640: begin l_1 = +16;
				 l_2 = +22; end
		14658: begin l_1 = +16;
				 l_2 = -22; end
		2961: begin l_1 = -16;
				 l_2 = +22; end
		1979: begin l_1 = -16;
				 l_2 = -22; end
		16131: begin l_1 = +16;
				 l_2 = +23; end
		14167: begin l_1 = +16;
				 l_2 = -23; end
		3452: begin l_1 = -16;
				 l_2 = +23; end
		1488: begin l_1 = -16;
				 l_2 = -23; end
		17113: begin l_1 = +16;
				 l_2 = +24; end
		13185: begin l_1 = +16;
				 l_2 = -24; end
		4434: begin l_1 = -16;
				 l_2 = +24; end
		506: begin l_1 = -16;
				 l_2 = -24; end
		1458: begin l_1 = +16;
				 l_2 = +25; end
		11221: begin l_1 = +16;
				 l_2 = -25; end
		6398: begin l_1 = -16;
				 l_2 = +25; end
		16161: begin l_1 = -16;
				 l_2 = -25; end
		5386: begin l_1 = +16;
				 l_2 = +26; end
		7293: begin l_1 = +16;
				 l_2 = -26; end
		10326: begin l_1 = -16;
				 l_2 = +26; end
		12233: begin l_1 = -16;
				 l_2 = -26; end
		13242: begin l_1 = +16;
				 l_2 = +27; end
		17056: begin l_1 = +16;
				 l_2 = -27; end
		563: begin l_1 = -16;
				 l_2 = +27; end
		4377: begin l_1 = -16;
				 l_2 = -27; end
		11335: begin l_1 = +16;
				 l_2 = +28; end
		1344: begin l_1 = +16;
				 l_2 = -28; end
		16275: begin l_1 = -16;
				 l_2 = +28; end
		6284: begin l_1 = -16;
				 l_2 = -28; end
		7521: begin l_1 = +16;
				 l_2 = +29; end
		5158: begin l_1 = +16;
				 l_2 = -29; end
		12461: begin l_1 = -16;
				 l_2 = +29; end
		10098: begin l_1 = -16;
				 l_2 = -29; end
		17512: begin l_1 = +16;
				 l_2 = +30; end
		12786: begin l_1 = +16;
				 l_2 = -30; end
		4833: begin l_1 = -16;
				 l_2 = +30; end
		107: begin l_1 = -16;
				 l_2 = -30; end
		2256: begin l_1 = +16;
				 l_2 = +31; end
		10423: begin l_1 = +16;
				 l_2 = -31; end
		7196: begin l_1 = -16;
				 l_2 = +31; end
		15363: begin l_1 = -16;
				 l_2 = -31; end
		6982: begin l_1 = +16;
				 l_2 = +32; end
		5697: begin l_1 = +16;
				 l_2 = -32; end
		11922: begin l_1 = -16;
				 l_2 = +32; end
		10637: begin l_1 = -16;
				 l_2 = -32; end
		16434: begin l_1 = +16;
				 l_2 = +33; end
		13864: begin l_1 = +16;
				 l_2 = -33; end
		3755: begin l_1 = -16;
				 l_2 = +33; end
		1185: begin l_1 = -16;
				 l_2 = -33; end
		100: begin l_1 = +16;
				 l_2 = +34; end
		12579: begin l_1 = +16;
				 l_2 = -34; end
		5040: begin l_1 = -16;
				 l_2 = +34; end
		17519: begin l_1 = -16;
				 l_2 = -34; end
		2670: begin l_1 = +16;
				 l_2 = +35; end
		10009: begin l_1 = +16;
				 l_2 = -35; end
		7610: begin l_1 = -16;
				 l_2 = +35; end
		14949: begin l_1 = -16;
				 l_2 = -35; end
		7810: begin l_1 = +16;
				 l_2 = +36; end
		4869: begin l_1 = +16;
				 l_2 = -36; end
		12750: begin l_1 = -16;
				 l_2 = +36; end
		9809: begin l_1 = -16;
				 l_2 = -36; end
		471: begin l_1 = +16;
				 l_2 = +37; end
		12208: begin l_1 = +16;
				 l_2 = -37; end
		5411: begin l_1 = -16;
				 l_2 = +37; end
		17148: begin l_1 = -16;
				 l_2 = -37; end
		3412: begin l_1 = +16;
				 l_2 = +38; end
		9267: begin l_1 = +16;
				 l_2 = -38; end
		8352: begin l_1 = -16;
				 l_2 = +38; end
		14207: begin l_1 = -16;
				 l_2 = -38; end
		9294: begin l_1 = +16;
				 l_2 = +39; end
		3385: begin l_1 = +16;
				 l_2 = -39; end
		14234: begin l_1 = -16;
				 l_2 = +39; end
		8325: begin l_1 = -16;
				 l_2 = -39; end
		3439: begin l_1 = +16;
				 l_2 = +40; end
		9240: begin l_1 = +16;
				 l_2 = -40; end
		8379: begin l_1 = -16;
				 l_2 = +40; end
		14180: begin l_1 = -16;
				 l_2 = -40; end
		9348: begin l_1 = +16;
				 l_2 = +41; end
		3331: begin l_1 = +16;
				 l_2 = -41; end
		14288: begin l_1 = -16;
				 l_2 = +41; end
		8271: begin l_1 = -16;
				 l_2 = -41; end
		3547: begin l_1 = +16;
				 l_2 = +42; end
		9132: begin l_1 = +16;
				 l_2 = -42; end
		8487: begin l_1 = -16;
				 l_2 = +42; end
		14072: begin l_1 = -16;
				 l_2 = -42; end
		9564: begin l_1 = +16;
				 l_2 = +43; end
		3115: begin l_1 = +16;
				 l_2 = -43; end
		14504: begin l_1 = -16;
				 l_2 = +43; end
		8055: begin l_1 = -16;
				 l_2 = -43; end
		2799: begin l_1 = -17;
				 l_2 = +19; end
		14820: begin l_1 = -17;
				 l_2 = -18; end
		10538: begin l_1 = +17;
				 l_2 = +19; end
		7081: begin l_1 = -17;
				 l_2 = -19; end
		8397: begin l_1 = +17;
				 l_2 = +20; end
		16961: begin l_1 = +17;
				 l_2 = -20; end
		658: begin l_1 = -17;
				 l_2 = +20; end
		9222: begin l_1 = -17;
				 l_2 = -20; end
		4115: begin l_1 = +17;
				 l_2 = +21; end
		3624: begin l_1 = +17;
				 l_2 = -21; end
		13995: begin l_1 = -17;
				 l_2 = +21; end
		13504: begin l_1 = -17;
				 l_2 = -21; end
		13170: begin l_1 = +17;
				 l_2 = +22; end
		12188: begin l_1 = +17;
				 l_2 = -22; end
		5431: begin l_1 = -17;
				 l_2 = +22; end
		4449: begin l_1 = -17;
				 l_2 = -22; end
		13661: begin l_1 = +17;
				 l_2 = +23; end
		11697: begin l_1 = +17;
				 l_2 = -23; end
		5922: begin l_1 = -17;
				 l_2 = +23; end
		3958: begin l_1 = -17;
				 l_2 = -23; end
		14643: begin l_1 = +17;
				 l_2 = +24; end
		10715: begin l_1 = +17;
				 l_2 = -24; end
		6904: begin l_1 = -17;
				 l_2 = +24; end
		2976: begin l_1 = -17;
				 l_2 = -24; end
		16607: begin l_1 = +17;
				 l_2 = +25; end
		8751: begin l_1 = +17;
				 l_2 = -25; end
		8868: begin l_1 = -17;
				 l_2 = +25; end
		1012: begin l_1 = -17;
				 l_2 = -25; end
		2916: begin l_1 = +17;
				 l_2 = +26; end
		4823: begin l_1 = +17;
				 l_2 = -26; end
		12796: begin l_1 = -17;
				 l_2 = +26; end
		14703: begin l_1 = -17;
				 l_2 = -26; end
		10772: begin l_1 = +17;
				 l_2 = +27; end
		14586: begin l_1 = +17;
				 l_2 = -27; end
		3033: begin l_1 = -17;
				 l_2 = +27; end
		6847: begin l_1 = -17;
				 l_2 = -27; end
		8865: begin l_1 = +17;
				 l_2 = +28; end
		16493: begin l_1 = +17;
				 l_2 = -28; end
		1126: begin l_1 = -17;
				 l_2 = +28; end
		8754: begin l_1 = -17;
				 l_2 = -28; end
		5051: begin l_1 = +17;
				 l_2 = +29; end
		2688: begin l_1 = +17;
				 l_2 = -29; end
		14931: begin l_1 = -17;
				 l_2 = +29; end
		12568: begin l_1 = -17;
				 l_2 = -29; end
		15042: begin l_1 = +17;
				 l_2 = +30; end
		10316: begin l_1 = +17;
				 l_2 = -30; end
		7303: begin l_1 = -17;
				 l_2 = +30; end
		2577: begin l_1 = -17;
				 l_2 = -30; end
		17405: begin l_1 = +17;
				 l_2 = +31; end
		7953: begin l_1 = +17;
				 l_2 = -31; end
		9666: begin l_1 = -17;
				 l_2 = +31; end
		214: begin l_1 = -17;
				 l_2 = -31; end
		4512: begin l_1 = +17;
				 l_2 = +32; end
		3227: begin l_1 = +17;
				 l_2 = -32; end
		14392: begin l_1 = -17;
				 l_2 = +32; end
		13107: begin l_1 = -17;
				 l_2 = -32; end
		13964: begin l_1 = +17;
				 l_2 = +33; end
		11394: begin l_1 = +17;
				 l_2 = -33; end
		6225: begin l_1 = -17;
				 l_2 = +33; end
		3655: begin l_1 = -17;
				 l_2 = -33; end
		15249: begin l_1 = +17;
				 l_2 = +34; end
		10109: begin l_1 = +17;
				 l_2 = -34; end
		7510: begin l_1 = -17;
				 l_2 = +34; end
		2370: begin l_1 = -17;
				 l_2 = -34; end
		200: begin l_1 = +17;
				 l_2 = +35; end
		7539: begin l_1 = +17;
				 l_2 = -35; end
		10080: begin l_1 = -17;
				 l_2 = +35; end
		17419: begin l_1 = -17;
				 l_2 = -35; end
		5340: begin l_1 = +17;
				 l_2 = +36; end
		2399: begin l_1 = +17;
				 l_2 = -36; end
		15220: begin l_1 = -17;
				 l_2 = +36; end
		12279: begin l_1 = -17;
				 l_2 = -36; end
		15620: begin l_1 = +17;
				 l_2 = +37; end
		9738: begin l_1 = +17;
				 l_2 = -37; end
		7881: begin l_1 = -17;
				 l_2 = +37; end
		1999: begin l_1 = -17;
				 l_2 = -37; end
		942: begin l_1 = +17;
				 l_2 = +38; end
		6797: begin l_1 = +17;
				 l_2 = -38; end
		10822: begin l_1 = -17;
				 l_2 = +38; end
		16677: begin l_1 = -17;
				 l_2 = -38; end
		6824: begin l_1 = +17;
				 l_2 = +39; end
		915: begin l_1 = +17;
				 l_2 = -39; end
		16704: begin l_1 = -17;
				 l_2 = +39; end
		10795: begin l_1 = -17;
				 l_2 = -39; end
		969: begin l_1 = +17;
				 l_2 = +40; end
		6770: begin l_1 = +17;
				 l_2 = -40; end
		10849: begin l_1 = -17;
				 l_2 = +40; end
		16650: begin l_1 = -17;
				 l_2 = -40; end
		6878: begin l_1 = +17;
				 l_2 = +41; end
		861: begin l_1 = +17;
				 l_2 = -41; end
		16758: begin l_1 = -17;
				 l_2 = +41; end
		10741: begin l_1 = -17;
				 l_2 = -41; end
		1077: begin l_1 = +17;
				 l_2 = +42; end
		6662: begin l_1 = +17;
				 l_2 = -42; end
		10957: begin l_1 = -17;
				 l_2 = +42; end
		16542: begin l_1 = -17;
				 l_2 = -42; end
		7094: begin l_1 = +17;
				 l_2 = +43; end
		645: begin l_1 = +17;
				 l_2 = -43; end
		16974: begin l_1 = -17;
				 l_2 = +43; end
		10525: begin l_1 = -17;
				 l_2 = -43; end
		5598: begin l_1 = -18;
				 l_2 = +20; end
		12021: begin l_1 = -18;
				 l_2 = -19; end
		3457: begin l_1 = +18;
				 l_2 = +20; end
		14162: begin l_1 = -18;
				 l_2 = -20; end
		16794: begin l_1 = +18;
				 l_2 = +21; end
		16303: begin l_1 = +18;
				 l_2 = -21; end
		1316: begin l_1 = -18;
				 l_2 = +21; end
		825: begin l_1 = -18;
				 l_2 = -21; end
		8230: begin l_1 = +18;
				 l_2 = +22; end
		7248: begin l_1 = +18;
				 l_2 = -22; end
		10371: begin l_1 = -18;
				 l_2 = +22; end
		9389: begin l_1 = -18;
				 l_2 = -22; end
		8721: begin l_1 = +18;
				 l_2 = +23; end
		6757: begin l_1 = +18;
				 l_2 = -23; end
		10862: begin l_1 = -18;
				 l_2 = +23; end
		8898: begin l_1 = -18;
				 l_2 = -23; end
		9703: begin l_1 = +18;
				 l_2 = +24; end
		5775: begin l_1 = +18;
				 l_2 = -24; end
		11844: begin l_1 = -18;
				 l_2 = +24; end
		7916: begin l_1 = -18;
				 l_2 = -24; end
		11667: begin l_1 = +18;
				 l_2 = +25; end
		3811: begin l_1 = +18;
				 l_2 = -25; end
		13808: begin l_1 = -18;
				 l_2 = +25; end
		5952: begin l_1 = -18;
				 l_2 = -25; end
		15595: begin l_1 = +18;
				 l_2 = +26; end
		17502: begin l_1 = +18;
				 l_2 = -26; end
		117: begin l_1 = -18;
				 l_2 = +26; end
		2024: begin l_1 = -18;
				 l_2 = -26; end
		5832: begin l_1 = +18;
				 l_2 = +27; end
		9646: begin l_1 = +18;
				 l_2 = -27; end
		7973: begin l_1 = -18;
				 l_2 = +27; end
		11787: begin l_1 = -18;
				 l_2 = -27; end
		3925: begin l_1 = +18;
				 l_2 = +28; end
		11553: begin l_1 = +18;
				 l_2 = -28; end
		6066: begin l_1 = -18;
				 l_2 = +28; end
		13694: begin l_1 = -18;
				 l_2 = -28; end
		111: begin l_1 = +18;
				 l_2 = +29; end
		15367: begin l_1 = +18;
				 l_2 = -29; end
		2252: begin l_1 = -18;
				 l_2 = +29; end
		17508: begin l_1 = -18;
				 l_2 = -29; end
		10102: begin l_1 = +18;
				 l_2 = +30; end
		5376: begin l_1 = +18;
				 l_2 = -30; end
		12243: begin l_1 = -18;
				 l_2 = +30; end
		7517: begin l_1 = -18;
				 l_2 = -30; end
		12465: begin l_1 = +18;
				 l_2 = +31; end
		3013: begin l_1 = +18;
				 l_2 = -31; end
		14606: begin l_1 = -18;
				 l_2 = +31; end
		5154: begin l_1 = -18;
				 l_2 = -31; end
		17191: begin l_1 = +18;
				 l_2 = +32; end
		15906: begin l_1 = +18;
				 l_2 = -32; end
		1713: begin l_1 = -18;
				 l_2 = +32; end
		428: begin l_1 = -18;
				 l_2 = -32; end
		9024: begin l_1 = +18;
				 l_2 = +33; end
		6454: begin l_1 = +18;
				 l_2 = -33; end
		11165: begin l_1 = -18;
				 l_2 = +33; end
		8595: begin l_1 = -18;
				 l_2 = -33; end
		10309: begin l_1 = +18;
				 l_2 = +34; end
		5169: begin l_1 = +18;
				 l_2 = -34; end
		12450: begin l_1 = -18;
				 l_2 = +34; end
		7310: begin l_1 = -18;
				 l_2 = -34; end
		12879: begin l_1 = +18;
				 l_2 = +35; end
		2599: begin l_1 = +18;
				 l_2 = -35; end
		15020: begin l_1 = -18;
				 l_2 = +35; end
		4740: begin l_1 = -18;
				 l_2 = -35; end
		400: begin l_1 = +18;
				 l_2 = +36; end
		15078: begin l_1 = +18;
				 l_2 = -36; end
		2541: begin l_1 = -18;
				 l_2 = +36; end
		17219: begin l_1 = -18;
				 l_2 = -36; end
		10680: begin l_1 = +18;
				 l_2 = +37; end
		4798: begin l_1 = +18;
				 l_2 = -37; end
		12821: begin l_1 = -18;
				 l_2 = +37; end
		6939: begin l_1 = -18;
				 l_2 = -37; end
		13621: begin l_1 = +18;
				 l_2 = +38; end
		1857: begin l_1 = +18;
				 l_2 = -38; end
		15762: begin l_1 = -18;
				 l_2 = +38; end
		3998: begin l_1 = -18;
				 l_2 = -38; end
		1884: begin l_1 = +18;
				 l_2 = +39; end
		13594: begin l_1 = +18;
				 l_2 = -39; end
		4025: begin l_1 = -18;
				 l_2 = +39; end
		15735: begin l_1 = -18;
				 l_2 = -39; end
		13648: begin l_1 = +18;
				 l_2 = +40; end
		1830: begin l_1 = +18;
				 l_2 = -40; end
		15789: begin l_1 = -18;
				 l_2 = +40; end
		3971: begin l_1 = -18;
				 l_2 = -40; end
		1938: begin l_1 = +18;
				 l_2 = +41; end
		13540: begin l_1 = +18;
				 l_2 = -41; end
		4079: begin l_1 = -18;
				 l_2 = +41; end
		15681: begin l_1 = -18;
				 l_2 = -41; end
		13756: begin l_1 = +18;
				 l_2 = +42; end
		1722: begin l_1 = +18;
				 l_2 = -42; end
		15897: begin l_1 = -18;
				 l_2 = +42; end
		3863: begin l_1 = -18;
				 l_2 = -42; end
		2154: begin l_1 = +18;
				 l_2 = +43; end
		13324: begin l_1 = +18;
				 l_2 = -43; end
		4295: begin l_1 = -18;
				 l_2 = +43; end
		15465: begin l_1 = -18;
				 l_2 = -43; end
		11196: begin l_1 = -19;
				 l_2 = +21; end
		6423: begin l_1 = -19;
				 l_2 = -20; end
		6914: begin l_1 = +19;
				 l_2 = +21; end
		10705: begin l_1 = -19;
				 l_2 = -21; end
		15969: begin l_1 = +19;
				 l_2 = +22; end
		14987: begin l_1 = +19;
				 l_2 = -22; end
		2632: begin l_1 = -19;
				 l_2 = +22; end
		1650: begin l_1 = -19;
				 l_2 = -22; end
		16460: begin l_1 = +19;
				 l_2 = +23; end
		14496: begin l_1 = +19;
				 l_2 = -23; end
		3123: begin l_1 = -19;
				 l_2 = +23; end
		1159: begin l_1 = -19;
				 l_2 = -23; end
		17442: begin l_1 = +19;
				 l_2 = +24; end
		13514: begin l_1 = +19;
				 l_2 = -24; end
		4105: begin l_1 = -19;
				 l_2 = +24; end
		177: begin l_1 = -19;
				 l_2 = -24; end
		1787: begin l_1 = +19;
				 l_2 = +25; end
		11550: begin l_1 = +19;
				 l_2 = -25; end
		6069: begin l_1 = -19;
				 l_2 = +25; end
		15832: begin l_1 = -19;
				 l_2 = -25; end
		5715: begin l_1 = +19;
				 l_2 = +26; end
		7622: begin l_1 = +19;
				 l_2 = -26; end
		9997: begin l_1 = -19;
				 l_2 = +26; end
		11904: begin l_1 = -19;
				 l_2 = -26; end
		13571: begin l_1 = +19;
				 l_2 = +27; end
		17385: begin l_1 = +19;
				 l_2 = -27; end
		234: begin l_1 = -19;
				 l_2 = +27; end
		4048: begin l_1 = -19;
				 l_2 = -27; end
		11664: begin l_1 = +19;
				 l_2 = +28; end
		1673: begin l_1 = +19;
				 l_2 = -28; end
		15946: begin l_1 = -19;
				 l_2 = +28; end
		5955: begin l_1 = -19;
				 l_2 = -28; end
		7850: begin l_1 = +19;
				 l_2 = +29; end
		5487: begin l_1 = +19;
				 l_2 = -29; end
		12132: begin l_1 = -19;
				 l_2 = +29; end
		9769: begin l_1 = -19;
				 l_2 = -29; end
		222: begin l_1 = +19;
				 l_2 = +30; end
		13115: begin l_1 = +19;
				 l_2 = -30; end
		4504: begin l_1 = -19;
				 l_2 = +30; end
		17397: begin l_1 = -19;
				 l_2 = -30; end
		2585: begin l_1 = +19;
				 l_2 = +31; end
		10752: begin l_1 = +19;
				 l_2 = -31; end
		6867: begin l_1 = -19;
				 l_2 = +31; end
		15034: begin l_1 = -19;
				 l_2 = -31; end
		7311: begin l_1 = +19;
				 l_2 = +32; end
		6026: begin l_1 = +19;
				 l_2 = -32; end
		11593: begin l_1 = -19;
				 l_2 = +32; end
		10308: begin l_1 = -19;
				 l_2 = -32; end
		16763: begin l_1 = +19;
				 l_2 = +33; end
		14193: begin l_1 = +19;
				 l_2 = -33; end
		3426: begin l_1 = -19;
				 l_2 = +33; end
		856: begin l_1 = -19;
				 l_2 = -33; end
		429: begin l_1 = +19;
				 l_2 = +34; end
		12908: begin l_1 = +19;
				 l_2 = -34; end
		4711: begin l_1 = -19;
				 l_2 = +34; end
		17190: begin l_1 = -19;
				 l_2 = -34; end
		2999: begin l_1 = +19;
				 l_2 = +35; end
		10338: begin l_1 = +19;
				 l_2 = -35; end
		7281: begin l_1 = -19;
				 l_2 = +35; end
		14620: begin l_1 = -19;
				 l_2 = -35; end
		8139: begin l_1 = +19;
				 l_2 = +36; end
		5198: begin l_1 = +19;
				 l_2 = -36; end
		12421: begin l_1 = -19;
				 l_2 = +36; end
		9480: begin l_1 = -19;
				 l_2 = -36; end
		800: begin l_1 = +19;
				 l_2 = +37; end
		12537: begin l_1 = +19;
				 l_2 = -37; end
		5082: begin l_1 = -19;
				 l_2 = +37; end
		16819: begin l_1 = -19;
				 l_2 = -37; end
		3741: begin l_1 = +19;
				 l_2 = +38; end
		9596: begin l_1 = +19;
				 l_2 = -38; end
		8023: begin l_1 = -19;
				 l_2 = +38; end
		13878: begin l_1 = -19;
				 l_2 = -38; end
		9623: begin l_1 = +19;
				 l_2 = +39; end
		3714: begin l_1 = +19;
				 l_2 = -39; end
		13905: begin l_1 = -19;
				 l_2 = +39; end
		7996: begin l_1 = -19;
				 l_2 = -39; end
		3768: begin l_1 = +19;
				 l_2 = +40; end
		9569: begin l_1 = +19;
				 l_2 = -40; end
		8050: begin l_1 = -19;
				 l_2 = +40; end
		13851: begin l_1 = -19;
				 l_2 = -40; end
		9677: begin l_1 = +19;
				 l_2 = +41; end
		3660: begin l_1 = +19;
				 l_2 = -41; end
		13959: begin l_1 = -19;
				 l_2 = +41; end
		7942: begin l_1 = -19;
				 l_2 = -41; end
		3876: begin l_1 = +19;
				 l_2 = +42; end
		9461: begin l_1 = +19;
				 l_2 = -42; end
		8158: begin l_1 = -19;
				 l_2 = +42; end
		13743: begin l_1 = -19;
				 l_2 = -42; end
		9893: begin l_1 = +19;
				 l_2 = +43; end
		3444: begin l_1 = +19;
				 l_2 = -43; end
		14175: begin l_1 = -19;
				 l_2 = +43; end
		7726: begin l_1 = -19;
				 l_2 = -43; end
		4773: begin l_1 = -20;
				 l_2 = +22; end
		12846: begin l_1 = -20;
				 l_2 = -21; end
		13828: begin l_1 = +20;
				 l_2 = +22; end
		3791: begin l_1 = -20;
				 l_2 = -22; end
		14319: begin l_1 = +20;
				 l_2 = +23; end
		12355: begin l_1 = +20;
				 l_2 = -23; end
		5264: begin l_1 = -20;
				 l_2 = +23; end
		3300: begin l_1 = -20;
				 l_2 = -23; end
		15301: begin l_1 = +20;
				 l_2 = +24; end
		11373: begin l_1 = +20;
				 l_2 = -24; end
		6246: begin l_1 = -20;
				 l_2 = +24; end
		2318: begin l_1 = -20;
				 l_2 = -24; end
		17265: begin l_1 = +20;
				 l_2 = +25; end
		9409: begin l_1 = +20;
				 l_2 = -25; end
		8210: begin l_1 = -20;
				 l_2 = +25; end
		354: begin l_1 = -20;
				 l_2 = -25; end
		3574: begin l_1 = +20;
				 l_2 = +26; end
		5481: begin l_1 = +20;
				 l_2 = -26; end
		12138: begin l_1 = -20;
				 l_2 = +26; end
		14045: begin l_1 = -20;
				 l_2 = -26; end
		11430: begin l_1 = +20;
				 l_2 = +27; end
		15244: begin l_1 = +20;
				 l_2 = -27; end
		2375: begin l_1 = -20;
				 l_2 = +27; end
		6189: begin l_1 = -20;
				 l_2 = -27; end
		9523: begin l_1 = +20;
				 l_2 = +28; end
		17151: begin l_1 = +20;
				 l_2 = -28; end
		468: begin l_1 = -20;
				 l_2 = +28; end
		8096: begin l_1 = -20;
				 l_2 = -28; end
		5709: begin l_1 = +20;
				 l_2 = +29; end
		3346: begin l_1 = +20;
				 l_2 = -29; end
		14273: begin l_1 = -20;
				 l_2 = +29; end
		11910: begin l_1 = -20;
				 l_2 = -29; end
		15700: begin l_1 = +20;
				 l_2 = +30; end
		10974: begin l_1 = +20;
				 l_2 = -30; end
		6645: begin l_1 = -20;
				 l_2 = +30; end
		1919: begin l_1 = -20;
				 l_2 = -30; end
		444: begin l_1 = +20;
				 l_2 = +31; end
		8611: begin l_1 = +20;
				 l_2 = -31; end
		9008: begin l_1 = -20;
				 l_2 = +31; end
		17175: begin l_1 = -20;
				 l_2 = -31; end
		5170: begin l_1 = +20;
				 l_2 = +32; end
		3885: begin l_1 = +20;
				 l_2 = -32; end
		13734: begin l_1 = -20;
				 l_2 = +32; end
		12449: begin l_1 = -20;
				 l_2 = -32; end
		14622: begin l_1 = +20;
				 l_2 = +33; end
		12052: begin l_1 = +20;
				 l_2 = -33; end
		5567: begin l_1 = -20;
				 l_2 = +33; end
		2997: begin l_1 = -20;
				 l_2 = -33; end
		15907: begin l_1 = +20;
				 l_2 = +34; end
		10767: begin l_1 = +20;
				 l_2 = -34; end
		6852: begin l_1 = -20;
				 l_2 = +34; end
		1712: begin l_1 = -20;
				 l_2 = -34; end
		858: begin l_1 = +20;
				 l_2 = +35; end
		8197: begin l_1 = +20;
				 l_2 = -35; end
		9422: begin l_1 = -20;
				 l_2 = +35; end
		16761: begin l_1 = -20;
				 l_2 = -35; end
		5998: begin l_1 = +20;
				 l_2 = +36; end
		3057: begin l_1 = +20;
				 l_2 = -36; end
		14562: begin l_1 = -20;
				 l_2 = +36; end
		11621: begin l_1 = -20;
				 l_2 = -36; end
		16278: begin l_1 = +20;
				 l_2 = +37; end
		10396: begin l_1 = +20;
				 l_2 = -37; end
		7223: begin l_1 = -20;
				 l_2 = +37; end
		1341: begin l_1 = -20;
				 l_2 = -37; end
		1600: begin l_1 = +20;
				 l_2 = +38; end
		7455: begin l_1 = +20;
				 l_2 = -38; end
		10164: begin l_1 = -20;
				 l_2 = +38; end
		16019: begin l_1 = -20;
				 l_2 = -38; end
		7482: begin l_1 = +20;
				 l_2 = +39; end
		1573: begin l_1 = +20;
				 l_2 = -39; end
		16046: begin l_1 = -20;
				 l_2 = +39; end
		10137: begin l_1 = -20;
				 l_2 = -39; end
		1627: begin l_1 = +20;
				 l_2 = +40; end
		7428: begin l_1 = +20;
				 l_2 = -40; end
		10191: begin l_1 = -20;
				 l_2 = +40; end
		15992: begin l_1 = -20;
				 l_2 = -40; end
		7536: begin l_1 = +20;
				 l_2 = +41; end
		1519: begin l_1 = +20;
				 l_2 = -41; end
		16100: begin l_1 = -20;
				 l_2 = +41; end
		10083: begin l_1 = -20;
				 l_2 = -41; end
		1735: begin l_1 = +20;
				 l_2 = +42; end
		7320: begin l_1 = +20;
				 l_2 = -42; end
		10299: begin l_1 = -20;
				 l_2 = +42; end
		15884: begin l_1 = -20;
				 l_2 = -42; end
		7752: begin l_1 = +20;
				 l_2 = +43; end
		1303: begin l_1 = +20;
				 l_2 = -43; end
		16316: begin l_1 = -20;
				 l_2 = +43; end
		9867: begin l_1 = -20;
				 l_2 = -43; end
		9546: begin l_1 = -21;
				 l_2 = +23; end
		8073: begin l_1 = -21;
				 l_2 = -22; end
		10037: begin l_1 = +21;
				 l_2 = +23; end
		7582: begin l_1 = -21;
				 l_2 = -23; end
		11019: begin l_1 = +21;
				 l_2 = +24; end
		7091: begin l_1 = +21;
				 l_2 = -24; end
		10528: begin l_1 = -21;
				 l_2 = +24; end
		6600: begin l_1 = -21;
				 l_2 = -24; end
		12983: begin l_1 = +21;
				 l_2 = +25; end
		5127: begin l_1 = +21;
				 l_2 = -25; end
		12492: begin l_1 = -21;
				 l_2 = +25; end
		4636: begin l_1 = -21;
				 l_2 = -25; end
		16911: begin l_1 = +21;
				 l_2 = +26; end
		1199: begin l_1 = +21;
				 l_2 = -26; end
		16420: begin l_1 = -21;
				 l_2 = +26; end
		708: begin l_1 = -21;
				 l_2 = -26; end
		7148: begin l_1 = +21;
				 l_2 = +27; end
		10962: begin l_1 = +21;
				 l_2 = -27; end
		6657: begin l_1 = -21;
				 l_2 = +27; end
		10471: begin l_1 = -21;
				 l_2 = -27; end
		5241: begin l_1 = +21;
				 l_2 = +28; end
		12869: begin l_1 = +21;
				 l_2 = -28; end
		4750: begin l_1 = -21;
				 l_2 = +28; end
		12378: begin l_1 = -21;
				 l_2 = -28; end
		1427: begin l_1 = +21;
				 l_2 = +29; end
		16683: begin l_1 = +21;
				 l_2 = -29; end
		936: begin l_1 = -21;
				 l_2 = +29; end
		16192: begin l_1 = -21;
				 l_2 = -29; end
		11418: begin l_1 = +21;
				 l_2 = +30; end
		6692: begin l_1 = +21;
				 l_2 = -30; end
		10927: begin l_1 = -21;
				 l_2 = +30; end
		6201: begin l_1 = -21;
				 l_2 = -30; end
		13781: begin l_1 = +21;
				 l_2 = +31; end
		4329: begin l_1 = +21;
				 l_2 = -31; end
		13290: begin l_1 = -21;
				 l_2 = +31; end
		3838: begin l_1 = -21;
				 l_2 = -31; end
		888: begin l_1 = +21;
				 l_2 = +32; end
		17222: begin l_1 = +21;
				 l_2 = -32; end
		397: begin l_1 = -21;
				 l_2 = +32; end
		16731: begin l_1 = -21;
				 l_2 = -32; end
		10340: begin l_1 = +21;
				 l_2 = +33; end
		7770: begin l_1 = +21;
				 l_2 = -33; end
		9849: begin l_1 = -21;
				 l_2 = +33; end
		7279: begin l_1 = -21;
				 l_2 = -33; end
		11625: begin l_1 = +21;
				 l_2 = +34; end
		6485: begin l_1 = +21;
				 l_2 = -34; end
		11134: begin l_1 = -21;
				 l_2 = +34; end
		5994: begin l_1 = -21;
				 l_2 = -34; end
		14195: begin l_1 = +21;
				 l_2 = +35; end
		3915: begin l_1 = +21;
				 l_2 = -35; end
		13704: begin l_1 = -21;
				 l_2 = +35; end
		3424: begin l_1 = -21;
				 l_2 = -35; end
		1716: begin l_1 = +21;
				 l_2 = +36; end
		16394: begin l_1 = +21;
				 l_2 = -36; end
		1225: begin l_1 = -21;
				 l_2 = +36; end
		15903: begin l_1 = -21;
				 l_2 = -36; end
		11996: begin l_1 = +21;
				 l_2 = +37; end
		6114: begin l_1 = +21;
				 l_2 = -37; end
		11505: begin l_1 = -21;
				 l_2 = +37; end
		5623: begin l_1 = -21;
				 l_2 = -37; end
		14937: begin l_1 = +21;
				 l_2 = +38; end
		3173: begin l_1 = +21;
				 l_2 = -38; end
		14446: begin l_1 = -21;
				 l_2 = +38; end
		2682: begin l_1 = -21;
				 l_2 = -38; end
		3200: begin l_1 = +21;
				 l_2 = +39; end
		14910: begin l_1 = +21;
				 l_2 = -39; end
		2709: begin l_1 = -21;
				 l_2 = +39; end
		14419: begin l_1 = -21;
				 l_2 = -39; end
		14964: begin l_1 = +21;
				 l_2 = +40; end
		3146: begin l_1 = +21;
				 l_2 = -40; end
		14473: begin l_1 = -21;
				 l_2 = +40; end
		2655: begin l_1 = -21;
				 l_2 = -40; end
		3254: begin l_1 = +21;
				 l_2 = +41; end
		14856: begin l_1 = +21;
				 l_2 = -41; end
		2763: begin l_1 = -21;
				 l_2 = +41; end
		14365: begin l_1 = -21;
				 l_2 = -41; end
		15072: begin l_1 = +21;
				 l_2 = +42; end
		3038: begin l_1 = +21;
				 l_2 = -42; end
		14581: begin l_1 = -21;
				 l_2 = +42; end
		2547: begin l_1 = -21;
				 l_2 = -42; end
		3470: begin l_1 = +21;
				 l_2 = +43; end
		14640: begin l_1 = +21;
				 l_2 = -43; end
		2979: begin l_1 = -21;
				 l_2 = +43; end
		14149: begin l_1 = -21;
				 l_2 = -43; end
		1473: begin l_1 = -22;
				 l_2 = +24; end
		16146: begin l_1 = -22;
				 l_2 = -23; end
		2455: begin l_1 = +22;
				 l_2 = +24; end
		15164: begin l_1 = -22;
				 l_2 = -24; end
		4419: begin l_1 = +22;
				 l_2 = +25; end
		14182: begin l_1 = +22;
				 l_2 = -25; end
		3437: begin l_1 = -22;
				 l_2 = +25; end
		13200: begin l_1 = -22;
				 l_2 = -25; end
		8347: begin l_1 = +22;
				 l_2 = +26; end
		10254: begin l_1 = +22;
				 l_2 = -26; end
		7365: begin l_1 = -22;
				 l_2 = +26; end
		9272: begin l_1 = -22;
				 l_2 = -26; end
		16203: begin l_1 = +22;
				 l_2 = +27; end
		2398: begin l_1 = +22;
				 l_2 = -27; end
		15221: begin l_1 = -22;
				 l_2 = +27; end
		1416: begin l_1 = -22;
				 l_2 = -27; end
		14296: begin l_1 = +22;
				 l_2 = +28; end
		4305: begin l_1 = +22;
				 l_2 = -28; end
		13314: begin l_1 = -22;
				 l_2 = +28; end
		3323: begin l_1 = -22;
				 l_2 = -28; end
		10482: begin l_1 = +22;
				 l_2 = +29; end
		8119: begin l_1 = +22;
				 l_2 = -29; end
		9500: begin l_1 = -22;
				 l_2 = +29; end
		7137: begin l_1 = -22;
				 l_2 = -29; end
		2854: begin l_1 = +22;
				 l_2 = +30; end
		15747: begin l_1 = +22;
				 l_2 = -30; end
		1872: begin l_1 = -22;
				 l_2 = +30; end
		14765: begin l_1 = -22;
				 l_2 = -30; end
		5217: begin l_1 = +22;
				 l_2 = +31; end
		13384: begin l_1 = +22;
				 l_2 = -31; end
		4235: begin l_1 = -22;
				 l_2 = +31; end
		12402: begin l_1 = -22;
				 l_2 = -31; end
		9943: begin l_1 = +22;
				 l_2 = +32; end
		8658: begin l_1 = +22;
				 l_2 = -32; end
		8961: begin l_1 = -22;
				 l_2 = +32; end
		7676: begin l_1 = -22;
				 l_2 = -32; end
		1776: begin l_1 = +22;
				 l_2 = +33; end
		16825: begin l_1 = +22;
				 l_2 = -33; end
		794: begin l_1 = -22;
				 l_2 = +33; end
		15843: begin l_1 = -22;
				 l_2 = -33; end
		3061: begin l_1 = +22;
				 l_2 = +34; end
		15540: begin l_1 = +22;
				 l_2 = -34; end
		2079: begin l_1 = -22;
				 l_2 = +34; end
		14558: begin l_1 = -22;
				 l_2 = -34; end
		5631: begin l_1 = +22;
				 l_2 = +35; end
		12970: begin l_1 = +22;
				 l_2 = -35; end
		4649: begin l_1 = -22;
				 l_2 = +35; end
		11988: begin l_1 = -22;
				 l_2 = -35; end
		10771: begin l_1 = +22;
				 l_2 = +36; end
		7830: begin l_1 = +22;
				 l_2 = -36; end
		9789: begin l_1 = -22;
				 l_2 = +36; end
		6848: begin l_1 = -22;
				 l_2 = -36; end
		3432: begin l_1 = +22;
				 l_2 = +37; end
		15169: begin l_1 = +22;
				 l_2 = -37; end
		2450: begin l_1 = -22;
				 l_2 = +37; end
		14187: begin l_1 = -22;
				 l_2 = -37; end
		6373: begin l_1 = +22;
				 l_2 = +38; end
		12228: begin l_1 = +22;
				 l_2 = -38; end
		5391: begin l_1 = -22;
				 l_2 = +38; end
		11246: begin l_1 = -22;
				 l_2 = -38; end
		12255: begin l_1 = +22;
				 l_2 = +39; end
		6346: begin l_1 = +22;
				 l_2 = -39; end
		11273: begin l_1 = -22;
				 l_2 = +39; end
		5364: begin l_1 = -22;
				 l_2 = -39; end
		6400: begin l_1 = +22;
				 l_2 = +40; end
		12201: begin l_1 = +22;
				 l_2 = -40; end
		5418: begin l_1 = -22;
				 l_2 = +40; end
		11219: begin l_1 = -22;
				 l_2 = -40; end
		12309: begin l_1 = +22;
				 l_2 = +41; end
		6292: begin l_1 = +22;
				 l_2 = -41; end
		11327: begin l_1 = -22;
				 l_2 = +41; end
		5310: begin l_1 = -22;
				 l_2 = -41; end
		6508: begin l_1 = +22;
				 l_2 = +42; end
		12093: begin l_1 = +22;
				 l_2 = -42; end
		5526: begin l_1 = -22;
				 l_2 = +42; end
		11111: begin l_1 = -22;
				 l_2 = -42; end
		12525: begin l_1 = +22;
				 l_2 = +43; end
		6076: begin l_1 = +22;
				 l_2 = -43; end
		11543: begin l_1 = -22;
				 l_2 = +43; end
		5094: begin l_1 = -22;
				 l_2 = -43; end
		2946: begin l_1 = -23;
				 l_2 = +25; end
		14673: begin l_1 = -23;
				 l_2 = -24; end
		4910: begin l_1 = +23;
				 l_2 = +25; end
		12709: begin l_1 = -23;
				 l_2 = -25; end
		8838: begin l_1 = +23;
				 l_2 = +26; end
		10745: begin l_1 = +23;
				 l_2 = -26; end
		6874: begin l_1 = -23;
				 l_2 = +26; end
		8781: begin l_1 = -23;
				 l_2 = -26; end
		16694: begin l_1 = +23;
				 l_2 = +27; end
		2889: begin l_1 = +23;
				 l_2 = -27; end
		14730: begin l_1 = -23;
				 l_2 = +27; end
		925: begin l_1 = -23;
				 l_2 = -27; end
		14787: begin l_1 = +23;
				 l_2 = +28; end
		4796: begin l_1 = +23;
				 l_2 = -28; end
		12823: begin l_1 = -23;
				 l_2 = +28; end
		2832: begin l_1 = -23;
				 l_2 = -28; end
		10973: begin l_1 = +23;
				 l_2 = +29; end
		8610: begin l_1 = +23;
				 l_2 = -29; end
		9009: begin l_1 = -23;
				 l_2 = +29; end
		6646: begin l_1 = -23;
				 l_2 = -29; end
		3345: begin l_1 = +23;
				 l_2 = +30; end
		16238: begin l_1 = +23;
				 l_2 = -30; end
		1381: begin l_1 = -23;
				 l_2 = +30; end
		14274: begin l_1 = -23;
				 l_2 = -30; end
		5708: begin l_1 = +23;
				 l_2 = +31; end
		13875: begin l_1 = +23;
				 l_2 = -31; end
		3744: begin l_1 = -23;
				 l_2 = +31; end
		11911: begin l_1 = -23;
				 l_2 = -31; end
		10434: begin l_1 = +23;
				 l_2 = +32; end
		9149: begin l_1 = +23;
				 l_2 = -32; end
		8470: begin l_1 = -23;
				 l_2 = +32; end
		7185: begin l_1 = -23;
				 l_2 = -32; end
		2267: begin l_1 = +23;
				 l_2 = +33; end
		17316: begin l_1 = +23;
				 l_2 = -33; end
		303: begin l_1 = -23;
				 l_2 = +33; end
		15352: begin l_1 = -23;
				 l_2 = -33; end
		3552: begin l_1 = +23;
				 l_2 = +34; end
		16031: begin l_1 = +23;
				 l_2 = -34; end
		1588: begin l_1 = -23;
				 l_2 = +34; end
		14067: begin l_1 = -23;
				 l_2 = -34; end
		6122: begin l_1 = +23;
				 l_2 = +35; end
		13461: begin l_1 = +23;
				 l_2 = -35; end
		4158: begin l_1 = -23;
				 l_2 = +35; end
		11497: begin l_1 = -23;
				 l_2 = -35; end
		11262: begin l_1 = +23;
				 l_2 = +36; end
		8321: begin l_1 = +23;
				 l_2 = -36; end
		9298: begin l_1 = -23;
				 l_2 = +36; end
		6357: begin l_1 = -23;
				 l_2 = -36; end
		3923: begin l_1 = +23;
				 l_2 = +37; end
		15660: begin l_1 = +23;
				 l_2 = -37; end
		1959: begin l_1 = -23;
				 l_2 = +37; end
		13696: begin l_1 = -23;
				 l_2 = -37; end
		6864: begin l_1 = +23;
				 l_2 = +38; end
		12719: begin l_1 = +23;
				 l_2 = -38; end
		4900: begin l_1 = -23;
				 l_2 = +38; end
		10755: begin l_1 = -23;
				 l_2 = -38; end
		12746: begin l_1 = +23;
				 l_2 = +39; end
		6837: begin l_1 = +23;
				 l_2 = -39; end
		10782: begin l_1 = -23;
				 l_2 = +39; end
		4873: begin l_1 = -23;
				 l_2 = -39; end
		6891: begin l_1 = +23;
				 l_2 = +40; end
		12692: begin l_1 = +23;
				 l_2 = -40; end
		4927: begin l_1 = -23;
				 l_2 = +40; end
		10728: begin l_1 = -23;
				 l_2 = -40; end
		12800: begin l_1 = +23;
				 l_2 = +41; end
		6783: begin l_1 = +23;
				 l_2 = -41; end
		10836: begin l_1 = -23;
				 l_2 = +41; end
		4819: begin l_1 = -23;
				 l_2 = -41; end
		6999: begin l_1 = +23;
				 l_2 = +42; end
		12584: begin l_1 = +23;
				 l_2 = -42; end
		5035: begin l_1 = -23;
				 l_2 = +42; end
		10620: begin l_1 = -23;
				 l_2 = -42; end
		13016: begin l_1 = +23;
				 l_2 = +43; end
		6567: begin l_1 = +23;
				 l_2 = -43; end
		11052: begin l_1 = -23;
				 l_2 = +43; end
		4603: begin l_1 = -23;
				 l_2 = -43; end
		5892: begin l_1 = -24;
				 l_2 = +26; end
		11727: begin l_1 = -24;
				 l_2 = -25; end
		9820: begin l_1 = +24;
				 l_2 = +26; end
		7799: begin l_1 = -24;
				 l_2 = -26; end
		57: begin l_1 = +24;
				 l_2 = +27; end
		3871: begin l_1 = +24;
				 l_2 = -27; end
		13748: begin l_1 = -24;
				 l_2 = +27; end
		17562: begin l_1 = -24;
				 l_2 = -27; end
		15769: begin l_1 = +24;
				 l_2 = +28; end
		5778: begin l_1 = +24;
				 l_2 = -28; end
		11841: begin l_1 = -24;
				 l_2 = +28; end
		1850: begin l_1 = -24;
				 l_2 = -28; end
		11955: begin l_1 = +24;
				 l_2 = +29; end
		9592: begin l_1 = +24;
				 l_2 = -29; end
		8027: begin l_1 = -24;
				 l_2 = +29; end
		5664: begin l_1 = -24;
				 l_2 = -29; end
		4327: begin l_1 = +24;
				 l_2 = +30; end
		17220: begin l_1 = +24;
				 l_2 = -30; end
		399: begin l_1 = -24;
				 l_2 = +30; end
		13292: begin l_1 = -24;
				 l_2 = -30; end
		6690: begin l_1 = +24;
				 l_2 = +31; end
		14857: begin l_1 = +24;
				 l_2 = -31; end
		2762: begin l_1 = -24;
				 l_2 = +31; end
		10929: begin l_1 = -24;
				 l_2 = -31; end
		11416: begin l_1 = +24;
				 l_2 = +32; end
		10131: begin l_1 = +24;
				 l_2 = -32; end
		7488: begin l_1 = -24;
				 l_2 = +32; end
		6203: begin l_1 = -24;
				 l_2 = -32; end
		3249: begin l_1 = +24;
				 l_2 = +33; end
		679: begin l_1 = +24;
				 l_2 = -33; end
		16940: begin l_1 = -24;
				 l_2 = +33; end
		14370: begin l_1 = -24;
				 l_2 = -33; end
		4534: begin l_1 = +24;
				 l_2 = +34; end
		17013: begin l_1 = +24;
				 l_2 = -34; end
		606: begin l_1 = -24;
				 l_2 = +34; end
		13085: begin l_1 = -24;
				 l_2 = -34; end
		7104: begin l_1 = +24;
				 l_2 = +35; end
		14443: begin l_1 = +24;
				 l_2 = -35; end
		3176: begin l_1 = -24;
				 l_2 = +35; end
		10515: begin l_1 = -24;
				 l_2 = -35; end
		12244: begin l_1 = +24;
				 l_2 = +36; end
		9303: begin l_1 = +24;
				 l_2 = -36; end
		8316: begin l_1 = -24;
				 l_2 = +36; end
		5375: begin l_1 = -24;
				 l_2 = -36; end
		4905: begin l_1 = +24;
				 l_2 = +37; end
		16642: begin l_1 = +24;
				 l_2 = -37; end
		977: begin l_1 = -24;
				 l_2 = +37; end
		12714: begin l_1 = -24;
				 l_2 = -37; end
		7846: begin l_1 = +24;
				 l_2 = +38; end
		13701: begin l_1 = +24;
				 l_2 = -38; end
		3918: begin l_1 = -24;
				 l_2 = +38; end
		9773: begin l_1 = -24;
				 l_2 = -38; end
		13728: begin l_1 = +24;
				 l_2 = +39; end
		7819: begin l_1 = +24;
				 l_2 = -39; end
		9800: begin l_1 = -24;
				 l_2 = +39; end
		3891: begin l_1 = -24;
				 l_2 = -39; end
		7873: begin l_1 = +24;
				 l_2 = +40; end
		13674: begin l_1 = +24;
				 l_2 = -40; end
		3945: begin l_1 = -24;
				 l_2 = +40; end
		9746: begin l_1 = -24;
				 l_2 = -40; end
		13782: begin l_1 = +24;
				 l_2 = +41; end
		7765: begin l_1 = +24;
				 l_2 = -41; end
		9854: begin l_1 = -24;
				 l_2 = +41; end
		3837: begin l_1 = -24;
				 l_2 = -41; end
		7981: begin l_1 = +24;
				 l_2 = +42; end
		13566: begin l_1 = +24;
				 l_2 = -42; end
		4053: begin l_1 = -24;
				 l_2 = +42; end
		9638: begin l_1 = -24;
				 l_2 = -42; end
		13998: begin l_1 = +24;
				 l_2 = +43; end
		7549: begin l_1 = +24;
				 l_2 = -43; end
		10070: begin l_1 = -24;
				 l_2 = +43; end
		3621: begin l_1 = -24;
				 l_2 = -43; end
		11784: begin l_1 = -25;
				 l_2 = +27; end
		5835: begin l_1 = -25;
				 l_2 = -26; end
		2021: begin l_1 = +25;
				 l_2 = +27; end
		15598: begin l_1 = -25;
				 l_2 = -27; end
		114: begin l_1 = +25;
				 l_2 = +28; end
		7742: begin l_1 = +25;
				 l_2 = -28; end
		9877: begin l_1 = -25;
				 l_2 = +28; end
		17505: begin l_1 = -25;
				 l_2 = -28; end
		13919: begin l_1 = +25;
				 l_2 = +29; end
		11556: begin l_1 = +25;
				 l_2 = -29; end
		6063: begin l_1 = -25;
				 l_2 = +29; end
		3700: begin l_1 = -25;
				 l_2 = -29; end
		6291: begin l_1 = +25;
				 l_2 = +30; end
		1565: begin l_1 = +25;
				 l_2 = -30; end
		16054: begin l_1 = -25;
				 l_2 = +30; end
		11328: begin l_1 = -25;
				 l_2 = -30; end
		8654: begin l_1 = +25;
				 l_2 = +31; end
		16821: begin l_1 = +25;
				 l_2 = -31; end
		798: begin l_1 = -25;
				 l_2 = +31; end
		8965: begin l_1 = -25;
				 l_2 = -31; end
		13380: begin l_1 = +25;
				 l_2 = +32; end
		12095: begin l_1 = +25;
				 l_2 = -32; end
		5524: begin l_1 = -25;
				 l_2 = +32; end
		4239: begin l_1 = -25;
				 l_2 = -32; end
		5213: begin l_1 = +25;
				 l_2 = +33; end
		2643: begin l_1 = +25;
				 l_2 = -33; end
		14976: begin l_1 = -25;
				 l_2 = +33; end
		12406: begin l_1 = -25;
				 l_2 = -33; end
		6498: begin l_1 = +25;
				 l_2 = +34; end
		1358: begin l_1 = +25;
				 l_2 = -34; end
		16261: begin l_1 = -25;
				 l_2 = +34; end
		11121: begin l_1 = -25;
				 l_2 = -34; end
		9068: begin l_1 = +25;
				 l_2 = +35; end
		16407: begin l_1 = +25;
				 l_2 = -35; end
		1212: begin l_1 = -25;
				 l_2 = +35; end
		8551: begin l_1 = -25;
				 l_2 = -35; end
		14208: begin l_1 = +25;
				 l_2 = +36; end
		11267: begin l_1 = +25;
				 l_2 = -36; end
		6352: begin l_1 = -25;
				 l_2 = +36; end
		3411: begin l_1 = -25;
				 l_2 = -36; end
		6869: begin l_1 = +25;
				 l_2 = +37; end
		987: begin l_1 = +25;
				 l_2 = -37; end
		16632: begin l_1 = -25;
				 l_2 = +37; end
		10750: begin l_1 = -25;
				 l_2 = -37; end
		9810: begin l_1 = +25;
				 l_2 = +38; end
		15665: begin l_1 = +25;
				 l_2 = -38; end
		1954: begin l_1 = -25;
				 l_2 = +38; end
		7809: begin l_1 = -25;
				 l_2 = -38; end
		15692: begin l_1 = +25;
				 l_2 = +39; end
		9783: begin l_1 = +25;
				 l_2 = -39; end
		7836: begin l_1 = -25;
				 l_2 = +39; end
		1927: begin l_1 = -25;
				 l_2 = -39; end
		9837: begin l_1 = +25;
				 l_2 = +40; end
		15638: begin l_1 = +25;
				 l_2 = -40; end
		1981: begin l_1 = -25;
				 l_2 = +40; end
		7782: begin l_1 = -25;
				 l_2 = -40; end
		15746: begin l_1 = +25;
				 l_2 = +41; end
		9729: begin l_1 = +25;
				 l_2 = -41; end
		7890: begin l_1 = -25;
				 l_2 = +41; end
		1873: begin l_1 = -25;
				 l_2 = -41; end
		9945: begin l_1 = +25;
				 l_2 = +42; end
		15530: begin l_1 = +25;
				 l_2 = -42; end
		2089: begin l_1 = -25;
				 l_2 = +42; end
		7674: begin l_1 = -25;
				 l_2 = -42; end
		15962: begin l_1 = +25;
				 l_2 = +43; end
		9513: begin l_1 = +25;
				 l_2 = -43; end
		8106: begin l_1 = -25;
				 l_2 = +43; end
		1657: begin l_1 = -25;
				 l_2 = -43; end
		5949: begin l_1 = -26;
				 l_2 = +28; end
		11670: begin l_1 = -26;
				 l_2 = -27; end
		4042: begin l_1 = +26;
				 l_2 = +28; end
		13577: begin l_1 = -26;
				 l_2 = -28; end
		228: begin l_1 = +26;
				 l_2 = +29; end
		15484: begin l_1 = +26;
				 l_2 = -29; end
		2135: begin l_1 = -26;
				 l_2 = +29; end
		17391: begin l_1 = -26;
				 l_2 = -29; end
		10219: begin l_1 = +26;
				 l_2 = +30; end
		5493: begin l_1 = +26;
				 l_2 = -30; end
		12126: begin l_1 = -26;
				 l_2 = +30; end
		7400: begin l_1 = -26;
				 l_2 = -30; end
		12582: begin l_1 = +26;
				 l_2 = +31; end
		3130: begin l_1 = +26;
				 l_2 = -31; end
		14489: begin l_1 = -26;
				 l_2 = +31; end
		5037: begin l_1 = -26;
				 l_2 = -31; end
		17308: begin l_1 = +26;
				 l_2 = +32; end
		16023: begin l_1 = +26;
				 l_2 = -32; end
		1596: begin l_1 = -26;
				 l_2 = +32; end
		311: begin l_1 = -26;
				 l_2 = -32; end
		9141: begin l_1 = +26;
				 l_2 = +33; end
		6571: begin l_1 = +26;
				 l_2 = -33; end
		11048: begin l_1 = -26;
				 l_2 = +33; end
		8478: begin l_1 = -26;
				 l_2 = -33; end
		10426: begin l_1 = +26;
				 l_2 = +34; end
		5286: begin l_1 = +26;
				 l_2 = -34; end
		12333: begin l_1 = -26;
				 l_2 = +34; end
		7193: begin l_1 = -26;
				 l_2 = -34; end
		12996: begin l_1 = +26;
				 l_2 = +35; end
		2716: begin l_1 = +26;
				 l_2 = -35; end
		14903: begin l_1 = -26;
				 l_2 = +35; end
		4623: begin l_1 = -26;
				 l_2 = -35; end
		517: begin l_1 = +26;
				 l_2 = +36; end
		15195: begin l_1 = +26;
				 l_2 = -36; end
		2424: begin l_1 = -26;
				 l_2 = +36; end
		17102: begin l_1 = -26;
				 l_2 = -36; end
		10797: begin l_1 = +26;
				 l_2 = +37; end
		4915: begin l_1 = +26;
				 l_2 = -37; end
		12704: begin l_1 = -26;
				 l_2 = +37; end
		6822: begin l_1 = -26;
				 l_2 = -37; end
		13738: begin l_1 = +26;
				 l_2 = +38; end
		1974: begin l_1 = +26;
				 l_2 = -38; end
		15645: begin l_1 = -26;
				 l_2 = +38; end
		3881: begin l_1 = -26;
				 l_2 = -38; end
		2001: begin l_1 = +26;
				 l_2 = +39; end
		13711: begin l_1 = +26;
				 l_2 = -39; end
		3908: begin l_1 = -26;
				 l_2 = +39; end
		15618: begin l_1 = -26;
				 l_2 = -39; end
		13765: begin l_1 = +26;
				 l_2 = +40; end
		1947: begin l_1 = +26;
				 l_2 = -40; end
		15672: begin l_1 = -26;
				 l_2 = +40; end
		3854: begin l_1 = -26;
				 l_2 = -40; end
		2055: begin l_1 = +26;
				 l_2 = +41; end
		13657: begin l_1 = +26;
				 l_2 = -41; end
		3962: begin l_1 = -26;
				 l_2 = +41; end
		15564: begin l_1 = -26;
				 l_2 = -41; end
		13873: begin l_1 = +26;
				 l_2 = +42; end
		1839: begin l_1 = +26;
				 l_2 = -42; end
		15780: begin l_1 = -26;
				 l_2 = +42; end
		3746: begin l_1 = -26;
				 l_2 = -42; end
		2271: begin l_1 = +26;
				 l_2 = +43; end
		13441: begin l_1 = +26;
				 l_2 = -43; end
		4178: begin l_1 = -26;
				 l_2 = +43; end
		15348: begin l_1 = -26;
				 l_2 = -43; end
		11898: begin l_1 = -27;
				 l_2 = +29; end
		5721: begin l_1 = -27;
				 l_2 = -28; end
		8084: begin l_1 = +27;
				 l_2 = +29; end
		9535: begin l_1 = -27;
				 l_2 = -29; end
		456: begin l_1 = +27;
				 l_2 = +30; end
		13349: begin l_1 = +27;
				 l_2 = -30; end
		4270: begin l_1 = -27;
				 l_2 = +30; end
		17163: begin l_1 = -27;
				 l_2 = -30; end
		2819: begin l_1 = +27;
				 l_2 = +31; end
		10986: begin l_1 = +27;
				 l_2 = -31; end
		6633: begin l_1 = -27;
				 l_2 = +31; end
		14800: begin l_1 = -27;
				 l_2 = -31; end
		7545: begin l_1 = +27;
				 l_2 = +32; end
		6260: begin l_1 = +27;
				 l_2 = -32; end
		11359: begin l_1 = -27;
				 l_2 = +32; end
		10074: begin l_1 = -27;
				 l_2 = -32; end
		16997: begin l_1 = +27;
				 l_2 = +33; end
		14427: begin l_1 = +27;
				 l_2 = -33; end
		3192: begin l_1 = -27;
				 l_2 = +33; end
		622: begin l_1 = -27;
				 l_2 = -33; end
		663: begin l_1 = +27;
				 l_2 = +34; end
		13142: begin l_1 = +27;
				 l_2 = -34; end
		4477: begin l_1 = -27;
				 l_2 = +34; end
		16956: begin l_1 = -27;
				 l_2 = -34; end
		3233: begin l_1 = +27;
				 l_2 = +35; end
		10572: begin l_1 = +27;
				 l_2 = -35; end
		7047: begin l_1 = -27;
				 l_2 = +35; end
		14386: begin l_1 = -27;
				 l_2 = -35; end
		8373: begin l_1 = +27;
				 l_2 = +36; end
		5432: begin l_1 = +27;
				 l_2 = -36; end
		12187: begin l_1 = -27;
				 l_2 = +36; end
		9246: begin l_1 = -27;
				 l_2 = -36; end
		1034: begin l_1 = +27;
				 l_2 = +37; end
		12771: begin l_1 = +27;
				 l_2 = -37; end
		4848: begin l_1 = -27;
				 l_2 = +37; end
		16585: begin l_1 = -27;
				 l_2 = -37; end
		3975: begin l_1 = +27;
				 l_2 = +38; end
		9830: begin l_1 = +27;
				 l_2 = -38; end
		7789: begin l_1 = -27;
				 l_2 = +38; end
		13644: begin l_1 = -27;
				 l_2 = -38; end
		9857: begin l_1 = +27;
				 l_2 = +39; end
		3948: begin l_1 = +27;
				 l_2 = -39; end
		13671: begin l_1 = -27;
				 l_2 = +39; end
		7762: begin l_1 = -27;
				 l_2 = -39; end
		4002: begin l_1 = +27;
				 l_2 = +40; end
		9803: begin l_1 = +27;
				 l_2 = -40; end
		7816: begin l_1 = -27;
				 l_2 = +40; end
		13617: begin l_1 = -27;
				 l_2 = -40; end
		9911: begin l_1 = +27;
				 l_2 = +41; end
		3894: begin l_1 = +27;
				 l_2 = -41; end
		13725: begin l_1 = -27;
				 l_2 = +41; end
		7708: begin l_1 = -27;
				 l_2 = -41; end
		4110: begin l_1 = +27;
				 l_2 = +42; end
		9695: begin l_1 = +27;
				 l_2 = -42; end
		7924: begin l_1 = -27;
				 l_2 = +42; end
		13509: begin l_1 = -27;
				 l_2 = -42; end
		10127: begin l_1 = +27;
				 l_2 = +43; end
		3678: begin l_1 = +27;
				 l_2 = -43; end
		13941: begin l_1 = -27;
				 l_2 = +43; end
		7492: begin l_1 = -27;
				 l_2 = -43; end
		6177: begin l_1 = -28;
				 l_2 = +30; end
		11442: begin l_1 = -28;
				 l_2 = -29; end
		16168: begin l_1 = +28;
				 l_2 = +30; end
		1451: begin l_1 = -28;
				 l_2 = -30; end
		912: begin l_1 = +28;
				 l_2 = +31; end
		9079: begin l_1 = +28;
				 l_2 = -31; end
		8540: begin l_1 = -28;
				 l_2 = +31; end
		16707: begin l_1 = -28;
				 l_2 = -31; end
		5638: begin l_1 = +28;
				 l_2 = +32; end
		4353: begin l_1 = +28;
				 l_2 = -32; end
		13266: begin l_1 = -28;
				 l_2 = +32; end
		11981: begin l_1 = -28;
				 l_2 = -32; end
		15090: begin l_1 = +28;
				 l_2 = +33; end
		12520: begin l_1 = +28;
				 l_2 = -33; end
		5099: begin l_1 = -28;
				 l_2 = +33; end
		2529: begin l_1 = -28;
				 l_2 = -33; end
		16375: begin l_1 = +28;
				 l_2 = +34; end
		11235: begin l_1 = +28;
				 l_2 = -34; end
		6384: begin l_1 = -28;
				 l_2 = +34; end
		1244: begin l_1 = -28;
				 l_2 = -34; end
		1326: begin l_1 = +28;
				 l_2 = +35; end
		8665: begin l_1 = +28;
				 l_2 = -35; end
		8954: begin l_1 = -28;
				 l_2 = +35; end
		16293: begin l_1 = -28;
				 l_2 = -35; end
		6466: begin l_1 = +28;
				 l_2 = +36; end
		3525: begin l_1 = +28;
				 l_2 = -36; end
		14094: begin l_1 = -28;
				 l_2 = +36; end
		11153: begin l_1 = -28;
				 l_2 = -36; end
		16746: begin l_1 = +28;
				 l_2 = +37; end
		10864: begin l_1 = +28;
				 l_2 = -37; end
		6755: begin l_1 = -28;
				 l_2 = +37; end
		873: begin l_1 = -28;
				 l_2 = -37; end
		2068: begin l_1 = +28;
				 l_2 = +38; end
		7923: begin l_1 = +28;
				 l_2 = -38; end
		9696: begin l_1 = -28;
				 l_2 = +38; end
		15551: begin l_1 = -28;
				 l_2 = -38; end
		7950: begin l_1 = +28;
				 l_2 = +39; end
		2041: begin l_1 = +28;
				 l_2 = -39; end
		15578: begin l_1 = -28;
				 l_2 = +39; end
		9669: begin l_1 = -28;
				 l_2 = -39; end
		2095: begin l_1 = +28;
				 l_2 = +40; end
		7896: begin l_1 = +28;
				 l_2 = -40; end
		9723: begin l_1 = -28;
				 l_2 = +40; end
		15524: begin l_1 = -28;
				 l_2 = -40; end
		8004: begin l_1 = +28;
				 l_2 = +41; end
		1987: begin l_1 = +28;
				 l_2 = -41; end
		15632: begin l_1 = -28;
				 l_2 = +41; end
		9615: begin l_1 = -28;
				 l_2 = -41; end
		2203: begin l_1 = +28;
				 l_2 = +42; end
		7788: begin l_1 = +28;
				 l_2 = -42; end
		9831: begin l_1 = -28;
				 l_2 = +42; end
		15416: begin l_1 = -28;
				 l_2 = -42; end
		8220: begin l_1 = +28;
				 l_2 = +43; end
		1771: begin l_1 = +28;
				 l_2 = -43; end
		15848: begin l_1 = -28;
				 l_2 = +43; end
		9399: begin l_1 = -28;
				 l_2 = -43; end
		12354: begin l_1 = -29;
				 l_2 = +31; end
		5265: begin l_1 = -29;
				 l_2 = -30; end
		14717: begin l_1 = +29;
				 l_2 = +31; end
		2902: begin l_1 = -29;
				 l_2 = -31; end
		1824: begin l_1 = +29;
				 l_2 = +32; end
		539: begin l_1 = +29;
				 l_2 = -32; end
		17080: begin l_1 = -29;
				 l_2 = +32; end
		15795: begin l_1 = -29;
				 l_2 = -32; end
		11276: begin l_1 = +29;
				 l_2 = +33; end
		8706: begin l_1 = +29;
				 l_2 = -33; end
		8913: begin l_1 = -29;
				 l_2 = +33; end
		6343: begin l_1 = -29;
				 l_2 = -33; end
		12561: begin l_1 = +29;
				 l_2 = +34; end
		7421: begin l_1 = +29;
				 l_2 = -34; end
		10198: begin l_1 = -29;
				 l_2 = +34; end
		5058: begin l_1 = -29;
				 l_2 = -34; end
		15131: begin l_1 = +29;
				 l_2 = +35; end
		4851: begin l_1 = +29;
				 l_2 = -35; end
		12768: begin l_1 = -29;
				 l_2 = +35; end
		2488: begin l_1 = -29;
				 l_2 = -35; end
		2652: begin l_1 = +29;
				 l_2 = +36; end
		17330: begin l_1 = +29;
				 l_2 = -36; end
		289: begin l_1 = -29;
				 l_2 = +36; end
		14967: begin l_1 = -29;
				 l_2 = -36; end
		12932: begin l_1 = +29;
				 l_2 = +37; end
		7050: begin l_1 = +29;
				 l_2 = -37; end
		10569: begin l_1 = -29;
				 l_2 = +37; end
		4687: begin l_1 = -29;
				 l_2 = -37; end
		15873: begin l_1 = +29;
				 l_2 = +38; end
		4109: begin l_1 = +29;
				 l_2 = -38; end
		13510: begin l_1 = -29;
				 l_2 = +38; end
		1746: begin l_1 = -29;
				 l_2 = -38; end
		4136: begin l_1 = +29;
				 l_2 = +39; end
		15846: begin l_1 = +29;
				 l_2 = -39; end
		1773: begin l_1 = -29;
				 l_2 = +39; end
		13483: begin l_1 = -29;
				 l_2 = -39; end
		15900: begin l_1 = +29;
				 l_2 = +40; end
		4082: begin l_1 = +29;
				 l_2 = -40; end
		13537: begin l_1 = -29;
				 l_2 = +40; end
		1719: begin l_1 = -29;
				 l_2 = -40; end
		4190: begin l_1 = +29;
				 l_2 = +41; end
		15792: begin l_1 = +29;
				 l_2 = -41; end
		1827: begin l_1 = -29;
				 l_2 = +41; end
		13429: begin l_1 = -29;
				 l_2 = -41; end
		16008: begin l_1 = +29;
				 l_2 = +42; end
		3974: begin l_1 = +29;
				 l_2 = -42; end
		13645: begin l_1 = -29;
				 l_2 = +42; end
		1611: begin l_1 = -29;
				 l_2 = -42; end
		4406: begin l_1 = +29;
				 l_2 = +43; end
		15576: begin l_1 = +29;
				 l_2 = -43; end
		2043: begin l_1 = -29;
				 l_2 = +43; end
		13213: begin l_1 = -29;
				 l_2 = -43; end
		7089: begin l_1 = -30;
				 l_2 = +32; end
		10530: begin l_1 = -30;
				 l_2 = -31; end
		11815: begin l_1 = +30;
				 l_2 = +32; end
		5804: begin l_1 = -30;
				 l_2 = -32; end
		3648: begin l_1 = +30;
				 l_2 = +33; end
		1078: begin l_1 = +30;
				 l_2 = -33; end
		16541: begin l_1 = -30;
				 l_2 = +33; end
		13971: begin l_1 = -30;
				 l_2 = -33; end
		4933: begin l_1 = +30;
				 l_2 = +34; end
		17412: begin l_1 = +30;
				 l_2 = -34; end
		207: begin l_1 = -30;
				 l_2 = +34; end
		12686: begin l_1 = -30;
				 l_2 = -34; end
		7503: begin l_1 = +30;
				 l_2 = +35; end
		14842: begin l_1 = +30;
				 l_2 = -35; end
		2777: begin l_1 = -30;
				 l_2 = +35; end
		10116: begin l_1 = -30;
				 l_2 = -35; end
		12643: begin l_1 = +30;
				 l_2 = +36; end
		9702: begin l_1 = +30;
				 l_2 = -36; end
		7917: begin l_1 = -30;
				 l_2 = +36; end
		4976: begin l_1 = -30;
				 l_2 = -36; end
		5304: begin l_1 = +30;
				 l_2 = +37; end
		17041: begin l_1 = +30;
				 l_2 = -37; end
		578: begin l_1 = -30;
				 l_2 = +37; end
		12315: begin l_1 = -30;
				 l_2 = -37; end
		8245: begin l_1 = +30;
				 l_2 = +38; end
		14100: begin l_1 = +30;
				 l_2 = -38; end
		3519: begin l_1 = -30;
				 l_2 = +38; end
		9374: begin l_1 = -30;
				 l_2 = -38; end
		14127: begin l_1 = +30;
				 l_2 = +39; end
		8218: begin l_1 = +30;
				 l_2 = -39; end
		9401: begin l_1 = -30;
				 l_2 = +39; end
		3492: begin l_1 = -30;
				 l_2 = -39; end
		8272: begin l_1 = +30;
				 l_2 = +40; end
		14073: begin l_1 = +30;
				 l_2 = -40; end
		3546: begin l_1 = -30;
				 l_2 = +40; end
		9347: begin l_1 = -30;
				 l_2 = -40; end
		14181: begin l_1 = +30;
				 l_2 = +41; end
		8164: begin l_1 = +30;
				 l_2 = -41; end
		9455: begin l_1 = -30;
				 l_2 = +41; end
		3438: begin l_1 = -30;
				 l_2 = -41; end
		8380: begin l_1 = +30;
				 l_2 = +42; end
		13965: begin l_1 = +30;
				 l_2 = -42; end
		3654: begin l_1 = -30;
				 l_2 = +42; end
		9239: begin l_1 = -30;
				 l_2 = -42; end
		14397: begin l_1 = +30;
				 l_2 = +43; end
		7948: begin l_1 = +30;
				 l_2 = -43; end
		9671: begin l_1 = -30;
				 l_2 = +43; end
		3222: begin l_1 = -30;
				 l_2 = -43; end
		14178: begin l_1 = -31;
				 l_2 = +33; end
		3441: begin l_1 = -31;
				 l_2 = -32; end
		6011: begin l_1 = +31;
				 l_2 = +33; end
		11608: begin l_1 = -31;
				 l_2 = -33; end
		7296: begin l_1 = +31;
				 l_2 = +34; end
		2156: begin l_1 = +31;
				 l_2 = -34; end
		15463: begin l_1 = -31;
				 l_2 = +34; end
		10323: begin l_1 = -31;
				 l_2 = -34; end
		9866: begin l_1 = +31;
				 l_2 = +35; end
		17205: begin l_1 = +31;
				 l_2 = -35; end
		414: begin l_1 = -31;
				 l_2 = +35; end
		7753: begin l_1 = -31;
				 l_2 = -35; end
		15006: begin l_1 = +31;
				 l_2 = +36; end
		12065: begin l_1 = +31;
				 l_2 = -36; end
		5554: begin l_1 = -31;
				 l_2 = +36; end
		2613: begin l_1 = -31;
				 l_2 = -36; end
		7667: begin l_1 = +31;
				 l_2 = +37; end
		1785: begin l_1 = +31;
				 l_2 = -37; end
		15834: begin l_1 = -31;
				 l_2 = +37; end
		9952: begin l_1 = -31;
				 l_2 = -37; end
		10608: begin l_1 = +31;
				 l_2 = +38; end
		16463: begin l_1 = +31;
				 l_2 = -38; end
		1156: begin l_1 = -31;
				 l_2 = +38; end
		7011: begin l_1 = -31;
				 l_2 = -38; end
		16490: begin l_1 = +31;
				 l_2 = +39; end
		10581: begin l_1 = +31;
				 l_2 = -39; end
		7038: begin l_1 = -31;
				 l_2 = +39; end
		1129: begin l_1 = -31;
				 l_2 = -39; end
		10635: begin l_1 = +31;
				 l_2 = +40; end
		16436: begin l_1 = +31;
				 l_2 = -40; end
		1183: begin l_1 = -31;
				 l_2 = +40; end
		6984: begin l_1 = -31;
				 l_2 = -40; end
		16544: begin l_1 = +31;
				 l_2 = +41; end
		10527: begin l_1 = +31;
				 l_2 = -41; end
		7092: begin l_1 = -31;
				 l_2 = +41; end
		1075: begin l_1 = -31;
				 l_2 = -41; end
		10743: begin l_1 = +31;
				 l_2 = +42; end
		16328: begin l_1 = +31;
				 l_2 = -42; end
		1291: begin l_1 = -31;
				 l_2 = +42; end
		6876: begin l_1 = -31;
				 l_2 = -42; end
		16760: begin l_1 = +31;
				 l_2 = +43; end
		10311: begin l_1 = +31;
				 l_2 = -43; end
		7308: begin l_1 = -31;
				 l_2 = +43; end
		859: begin l_1 = -31;
				 l_2 = -43; end
		10737: begin l_1 = -32;
				 l_2 = +34; end
		6882: begin l_1 = -32;
				 l_2 = -33; end
		12022: begin l_1 = +32;
				 l_2 = +34; end
		5597: begin l_1 = -32;
				 l_2 = -34; end
		14592: begin l_1 = +32;
				 l_2 = +35; end
		4312: begin l_1 = +32;
				 l_2 = -35; end
		13307: begin l_1 = -32;
				 l_2 = +35; end
		3027: begin l_1 = -32;
				 l_2 = -35; end
		2113: begin l_1 = +32;
				 l_2 = +36; end
		16791: begin l_1 = +32;
				 l_2 = -36; end
		828: begin l_1 = -32;
				 l_2 = +36; end
		15506: begin l_1 = -32;
				 l_2 = -36; end
		12393: begin l_1 = +32;
				 l_2 = +37; end
		6511: begin l_1 = +32;
				 l_2 = -37; end
		11108: begin l_1 = -32;
				 l_2 = +37; end
		5226: begin l_1 = -32;
				 l_2 = -37; end
		15334: begin l_1 = +32;
				 l_2 = +38; end
		3570: begin l_1 = +32;
				 l_2 = -38; end
		14049: begin l_1 = -32;
				 l_2 = +38; end
		2285: begin l_1 = -32;
				 l_2 = -38; end
		3597: begin l_1 = +32;
				 l_2 = +39; end
		15307: begin l_1 = +32;
				 l_2 = -39; end
		2312: begin l_1 = -32;
				 l_2 = +39; end
		14022: begin l_1 = -32;
				 l_2 = -39; end
		15361: begin l_1 = +32;
				 l_2 = +40; end
		3543: begin l_1 = +32;
				 l_2 = -40; end
		14076: begin l_1 = -32;
				 l_2 = +40; end
		2258: begin l_1 = -32;
				 l_2 = -40; end
		3651: begin l_1 = +32;
				 l_2 = +41; end
		15253: begin l_1 = +32;
				 l_2 = -41; end
		2366: begin l_1 = -32;
				 l_2 = +41; end
		13968: begin l_1 = -32;
				 l_2 = -41; end
		15469: begin l_1 = +32;
				 l_2 = +42; end
		3435: begin l_1 = +32;
				 l_2 = -42; end
		14184: begin l_1 = -32;
				 l_2 = +42; end
		2150: begin l_1 = -32;
				 l_2 = -42; end
		3867: begin l_1 = +32;
				 l_2 = +43; end
		15037: begin l_1 = +32;
				 l_2 = -43; end
		2582: begin l_1 = -32;
				 l_2 = +43; end
		13752: begin l_1 = -32;
				 l_2 = -43; end
		3855: begin l_1 = -33;
				 l_2 = +35; end
		13764: begin l_1 = -33;
				 l_2 = -34; end
		6425: begin l_1 = +33;
				 l_2 = +35; end
		11194: begin l_1 = -33;
				 l_2 = -35; end
		11565: begin l_1 = +33;
				 l_2 = +36; end
		8624: begin l_1 = +33;
				 l_2 = -36; end
		8995: begin l_1 = -33;
				 l_2 = +36; end
		6054: begin l_1 = -33;
				 l_2 = -36; end
		4226: begin l_1 = +33;
				 l_2 = +37; end
		15963: begin l_1 = +33;
				 l_2 = -37; end
		1656: begin l_1 = -33;
				 l_2 = +37; end
		13393: begin l_1 = -33;
				 l_2 = -37; end
		7167: begin l_1 = +33;
				 l_2 = +38; end
		13022: begin l_1 = +33;
				 l_2 = -38; end
		4597: begin l_1 = -33;
				 l_2 = +38; end
		10452: begin l_1 = -33;
				 l_2 = -38; end
		13049: begin l_1 = +33;
				 l_2 = +39; end
		7140: begin l_1 = +33;
				 l_2 = -39; end
		10479: begin l_1 = -33;
				 l_2 = +39; end
		4570: begin l_1 = -33;
				 l_2 = -39; end
		7194: begin l_1 = +33;
				 l_2 = +40; end
		12995: begin l_1 = +33;
				 l_2 = -40; end
		4624: begin l_1 = -33;
				 l_2 = +40; end
		10425: begin l_1 = -33;
				 l_2 = -40; end
		13103: begin l_1 = +33;
				 l_2 = +41; end
		7086: begin l_1 = +33;
				 l_2 = -41; end
		10533: begin l_1 = -33;
				 l_2 = +41; end
		4516: begin l_1 = -33;
				 l_2 = -41; end
		7302: begin l_1 = +33;
				 l_2 = +42; end
		12887: begin l_1 = +33;
				 l_2 = -42; end
		4732: begin l_1 = -33;
				 l_2 = +42; end
		10317: begin l_1 = -33;
				 l_2 = -42; end
		13319: begin l_1 = +33;
				 l_2 = +43; end
		6870: begin l_1 = +33;
				 l_2 = -43; end
		10749: begin l_1 = -33;
				 l_2 = +43; end
		4300: begin l_1 = -33;
				 l_2 = -43; end
		7710: begin l_1 = -34;
				 l_2 = +36; end
		9909: begin l_1 = -34;
				 l_2 = -35; end
		12850: begin l_1 = +34;
				 l_2 = +36; end
		4769: begin l_1 = -34;
				 l_2 = -36; end
		5511: begin l_1 = +34;
				 l_2 = +37; end
		17248: begin l_1 = +34;
				 l_2 = -37; end
		371: begin l_1 = -34;
				 l_2 = +37; end
		12108: begin l_1 = -34;
				 l_2 = -37; end
		8452: begin l_1 = +34;
				 l_2 = +38; end
		14307: begin l_1 = +34;
				 l_2 = -38; end
		3312: begin l_1 = -34;
				 l_2 = +38; end
		9167: begin l_1 = -34;
				 l_2 = -38; end
		14334: begin l_1 = +34;
				 l_2 = +39; end
		8425: begin l_1 = +34;
				 l_2 = -39; end
		9194: begin l_1 = -34;
				 l_2 = +39; end
		3285: begin l_1 = -34;
				 l_2 = -39; end
		8479: begin l_1 = +34;
				 l_2 = +40; end
		14280: begin l_1 = +34;
				 l_2 = -40; end
		3339: begin l_1 = -34;
				 l_2 = +40; end
		9140: begin l_1 = -34;
				 l_2 = -40; end
		14388: begin l_1 = +34;
				 l_2 = +41; end
		8371: begin l_1 = +34;
				 l_2 = -41; end
		9248: begin l_1 = -34;
				 l_2 = +41; end
		3231: begin l_1 = -34;
				 l_2 = -41; end
		8587: begin l_1 = +34;
				 l_2 = +42; end
		14172: begin l_1 = +34;
				 l_2 = -42; end
		3447: begin l_1 = -34;
				 l_2 = +42; end
		9032: begin l_1 = -34;
				 l_2 = -42; end
		14604: begin l_1 = +34;
				 l_2 = +43; end
		8155: begin l_1 = +34;
				 l_2 = -43; end
		9464: begin l_1 = -34;
				 l_2 = +43; end
		3015: begin l_1 = -34;
				 l_2 = -43; end
		15420: begin l_1 = -35;
				 l_2 = +37; end
		2199: begin l_1 = -35;
				 l_2 = -36; end
		8081: begin l_1 = +35;
				 l_2 = +37; end
		9538: begin l_1 = -35;
				 l_2 = -37; end
		11022: begin l_1 = +35;
				 l_2 = +38; end
		16877: begin l_1 = +35;
				 l_2 = -38; end
		742: begin l_1 = -35;
				 l_2 = +38; end
		6597: begin l_1 = -35;
				 l_2 = -38; end
		16904: begin l_1 = +35;
				 l_2 = +39; end
		10995: begin l_1 = +35;
				 l_2 = -39; end
		6624: begin l_1 = -35;
				 l_2 = +39; end
		715: begin l_1 = -35;
				 l_2 = -39; end
		11049: begin l_1 = +35;
				 l_2 = +40; end
		16850: begin l_1 = +35;
				 l_2 = -40; end
		769: begin l_1 = -35;
				 l_2 = +40; end
		6570: begin l_1 = -35;
				 l_2 = -40; end
		16958: begin l_1 = +35;
				 l_2 = +41; end
		10941: begin l_1 = +35;
				 l_2 = -41; end
		6678: begin l_1 = -35;
				 l_2 = +41; end
		661: begin l_1 = -35;
				 l_2 = -41; end
		11157: begin l_1 = +35;
				 l_2 = +42; end
		16742: begin l_1 = +35;
				 l_2 = -42; end
		877: begin l_1 = -35;
				 l_2 = +42; end
		6462: begin l_1 = -35;
				 l_2 = -42; end
		17174: begin l_1 = +35;
				 l_2 = +43; end
		10725: begin l_1 = +35;
				 l_2 = -43; end
		6894: begin l_1 = -35;
				 l_2 = +43; end
		445: begin l_1 = -35;
				 l_2 = -43; end
		13221: begin l_1 = -36;
				 l_2 = +38; end
		4398: begin l_1 = -36;
				 l_2 = -37; end
		16162: begin l_1 = +36;
				 l_2 = +38; end
		1457: begin l_1 = -36;
				 l_2 = -38; end
		4425: begin l_1 = +36;
				 l_2 = +39; end
		16135: begin l_1 = +36;
				 l_2 = -39; end
		1484: begin l_1 = -36;
				 l_2 = +39; end
		13194: begin l_1 = -36;
				 l_2 = -39; end
		16189: begin l_1 = +36;
				 l_2 = +40; end
		4371: begin l_1 = +36;
				 l_2 = -40; end
		13248: begin l_1 = -36;
				 l_2 = +40; end
		1430: begin l_1 = -36;
				 l_2 = -40; end
		4479: begin l_1 = +36;
				 l_2 = +41; end
		16081: begin l_1 = +36;
				 l_2 = -41; end
		1538: begin l_1 = -36;
				 l_2 = +41; end
		13140: begin l_1 = -36;
				 l_2 = -41; end
		16297: begin l_1 = +36;
				 l_2 = +42; end
		4263: begin l_1 = +36;
				 l_2 = -42; end
		13356: begin l_1 = -36;
				 l_2 = +42; end
		1322: begin l_1 = -36;
				 l_2 = -42; end
		4695: begin l_1 = +36;
				 l_2 = +43; end
		15865: begin l_1 = +36;
				 l_2 = -43; end
		1754: begin l_1 = -36;
				 l_2 = +43; end
		12924: begin l_1 = -36;
				 l_2 = -43; end
		8823: begin l_1 = -37;
				 l_2 = +39; end
		8796: begin l_1 = -37;
				 l_2 = -38; end
		14705: begin l_1 = +37;
				 l_2 = +39; end
		2914: begin l_1 = -37;
				 l_2 = -39; end
		8850: begin l_1 = +37;
				 l_2 = +40; end
		14651: begin l_1 = +37;
				 l_2 = -40; end
		2968: begin l_1 = -37;
				 l_2 = +40; end
		8769: begin l_1 = -37;
				 l_2 = -40; end
		14759: begin l_1 = +37;
				 l_2 = +41; end
		8742: begin l_1 = +37;
				 l_2 = -41; end
		8877: begin l_1 = -37;
				 l_2 = +41; end
		2860: begin l_1 = -37;
				 l_2 = -41; end
		8958: begin l_1 = +37;
				 l_2 = +42; end
		14543: begin l_1 = +37;
				 l_2 = -42; end
		3076: begin l_1 = -37;
				 l_2 = +42; end
		8661: begin l_1 = -37;
				 l_2 = -42; end
		14975: begin l_1 = +37;
				 l_2 = +43; end
		8526: begin l_1 = +37;
				 l_2 = -43; end
		9093: begin l_1 = -37;
				 l_2 = +43; end
		2644: begin l_1 = -37;
				 l_2 = -43; end
		27: begin l_1 = -38;
				 l_2 = +40; end
		17592: begin l_1 = -38;
				 l_2 = -39; end
		11791: begin l_1 = +38;
				 l_2 = +40; end
		5828: begin l_1 = -38;
				 l_2 = -40; end
		81: begin l_1 = +38;
				 l_2 = +41; end
		11683: begin l_1 = +38;
				 l_2 = -41; end
		5936: begin l_1 = -38;
				 l_2 = +41; end
		17538: begin l_1 = -38;
				 l_2 = -41; end
		11899: begin l_1 = +38;
				 l_2 = +42; end
		17484: begin l_1 = +38;
				 l_2 = -42; end
		135: begin l_1 = -38;
				 l_2 = +42; end
		5720: begin l_1 = -38;
				 l_2 = -42; end
		297: begin l_1 = +38;
				 l_2 = +43; end
		11467: begin l_1 = +38;
				 l_2 = -43; end
		6152: begin l_1 = -38;
				 l_2 = +43; end
		17322: begin l_1 = -38;
				 l_2 = -43; end
		54: begin l_1 = -39;
				 l_2 = +41; end
		17565: begin l_1 = -39;
				 l_2 = -40; end
		5963: begin l_1 = +39;
				 l_2 = +41; end
		11656: begin l_1 = -39;
				 l_2 = -41; end
		162: begin l_1 = +39;
				 l_2 = +42; end
		5747: begin l_1 = +39;
				 l_2 = -42; end
		11872: begin l_1 = -39;
				 l_2 = +42; end
		17457: begin l_1 = -39;
				 l_2 = -42; end
		6179: begin l_1 = +39;
				 l_2 = +43; end
		17349: begin l_1 = +39;
				 l_2 = -43; end
		270: begin l_1 = -39;
				 l_2 = +43; end
		11440: begin l_1 = -39;
				 l_2 = -43; end
		108: begin l_1 = -40;
				 l_2 = +42; end
		17511: begin l_1 = -40;
				 l_2 = -41; end
		11926: begin l_1 = +40;
				 l_2 = +42; end
		5693: begin l_1 = -40;
				 l_2 = -42; end
		324: begin l_1 = +40;
				 l_2 = +43; end
		11494: begin l_1 = +40;
				 l_2 = -43; end
		6125: begin l_1 = -40;
				 l_2 = +43; end
		17295: begin l_1 = -40;
				 l_2 = -43; end
		216: begin l_1 = -41;
				 l_2 = +43; end
		17403: begin l_1 = -41;
				 l_2 = -42; end
		6233: begin l_1 = +41;
				 l_2 = +43; end
		11386: begin l_1 = -41;
				 l_2 = -43; end
		432: begin l_1 = +42;
				 l_2 = +43; end
		17187: begin l_1 = -42;
				 l_2 = -43; end
		default: begin l_1 = 0;
					   l_2 = 0; end
	endcase
end

endmodule

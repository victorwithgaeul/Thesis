// Product (AN) Code SEC l-LUT
// SEC_lLUT20bits.v
// Received single error location l, output remainder r.
module SEC_lLUT20bits(l, r);
input	signed	[6:0]	l;
output	reg	[12:0]	r;
always@(*) begin
	case(l)
		1: r = 1;
		-1: r = 6310;
		2: r = 2;
		-2: r = 6309;
		3: r = 4;
		-3: r = 6307;
		4: r = 8;
		-4: r = 6303;
		5: r = 16;
		-5: r = 6295;
		6: r = 32;
		-6: r = 6279;
		7: r = 64;
		-7: r = 6247;
		8: r = 128;
		-8: r = 6183;
		9: r = 256;
		-9: r = 6055;
		10: r = 512;
		-10: r = 5799;
		11: r = 1024;
		-11: r = 5287;
		12: r = 2048;
		-12: r = 4263;
		13: r = 4096;
		-13: r = 2215;
		14: r = 1881;
		-14: r = 4430;
		15: r = 3762;
		-15: r = 2549;
		16: r = 1213;
		-16: r = 5098;
		17: r = 2426;
		-17: r = 3885;
		18: r = 4852;
		-18: r = 1459;
		19: r = 3393;
		-19: r = 2918;
		20: r = 475;
		-20: r = 5836;
		21: r = 950;
		-21: r = 5361;
		22: r = 1900;
		-22: r = 4411;
		23: r = 3800;
		-23: r = 2511;
		24: r = 1289;
		-24: r = 5022;
		25: r = 2578;
		-25: r = 3733;
		26: r = 5156;
		-26: r = 1155;
		27: r = 4001;
		-27: r = 2310;
		28: r = 1691;
		-28: r = 4620;
		29: r = 3382;
		-29: r = 2929;
		30: r = 453;
		-30: r = 5858;
		31: r = 906;
		-31: r = 5405;
		32: r = 1812;
		-32: r = 4499;
		33: r = 3624;
		-33: r = 2687;
		default: r = 0;
	endcase
end

endmodule

// Product (AN) Code DEC_LUT_Decoder
// DEC_LUT_Decoder52bits.v
// Received codeword W = AN + E, E is double AWE (E = e1 + e2), +2^i or -2^i.
module DEC_LUT_Decoder52bits_clk(clk, rst_n, W, found, N);

//=========================================================================
//   PARAMETER AND LOCALPARAM FOR FSM
//   W_BITS 要考慮 OVERFLOW 問題
//   N_BITS 也要考慮 OVERFLOW 問題
//=========================================================================
parameter A = 50861 , W_BITS = 69, A_BITS = 16 , N_BITS = 53;

localparam [1:0] idle=2'b00, pre=2'b01,load=2'b10, LUT=2'b11;

reg [1:0] ps;
//==========================================
//   INPUT AND OUTPUT DECLARATION
//==========================================
input   clk, rst_n;
input 	[W_BITS-1:0]	W;
output	reg  [N_BITS-1:0] N;
output  reg  found;

reg 	[N_BITS-1:0]	Q;
reg 	[A_BITS-1:0]	R;

reg	signed	[68:0]	Delta;
always@(*) begin
	case(R)
		1: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000000001;
		50860: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111111111;
		2: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000000010;
		50859: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111111110;
		4: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000000100;
		50857: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111111100;
		8: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000001000;
		50853: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111111000;
		16: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000010000;
		50845: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111110000;
		32: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000100000;
		50829: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111100000;
		64: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000001000000;
		50797: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111000000;
		128: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000010000000;
		50733: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111110000000;
		256: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000100000000;
		50605: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111100000000;
		512: Delta = 69'sb000000000000000000000000000000000000000000000000000000000001000000000;
		50349: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111000000000;
		1024: Delta = 69'sb000000000000000000000000000000000000000000000000000000000010000000000;
		49837: Delta = 69'sb111111111111111111111111111111111111111111111111111111111110000000000;
		2048: Delta = 69'sb000000000000000000000000000000000000000000000000000000000100000000000;
		48813: Delta = 69'sb111111111111111111111111111111111111111111111111111111111100000000000;
		4096: Delta = 69'sb000000000000000000000000000000000000000000000000000000001000000000000;
		46765: Delta = 69'sb111111111111111111111111111111111111111111111111111111111000000000000;
		8192: Delta = 69'sb000000000000000000000000000000000000000000000000000000010000000000000;
		42669: Delta = 69'sb111111111111111111111111111111111111111111111111111111110000000000000;
		16384: Delta = 69'sb000000000000000000000000000000000000000000000000000000100000000000000;
		34477: Delta = 69'sb111111111111111111111111111111111111111111111111111111100000000000000;
		32768: Delta = 69'sb000000000000000000000000000000000000000000000000000001000000000000000;
		18093: Delta = 69'sb111111111111111111111111111111111111111111111111111111000000000000000;
		14675: Delta = 69'sb000000000000000000000000000000000000000000000000000010000000000000000;
		36186: Delta = 69'sb111111111111111111111111111111111111111111111111111110000000000000000;
		29350: Delta = 69'sb000000000000000000000000000000000000000000000000000100000000000000000;
		21511: Delta = 69'sb111111111111111111111111111111111111111111111111111100000000000000000;
		7839: Delta = 69'sb000000000000000000000000000000000000000000000000001000000000000000000;
		43022: Delta = 69'sb111111111111111111111111111111111111111111111111111000000000000000000;
		15678: Delta = 69'sb000000000000000000000000000000000000000000000000010000000000000000000;
		35183: Delta = 69'sb111111111111111111111111111111111111111111111111110000000000000000000;
		31356: Delta = 69'sb000000000000000000000000000000000000000000000000100000000000000000000;
		19505: Delta = 69'sb111111111111111111111111111111111111111111111111100000000000000000000;
		11851: Delta = 69'sb000000000000000000000000000000000000000000000001000000000000000000000;
		39010: Delta = 69'sb111111111111111111111111111111111111111111111111000000000000000000000;
		23702: Delta = 69'sb000000000000000000000000000000000000000000000010000000000000000000000;
		27159: Delta = 69'sb111111111111111111111111111111111111111111111110000000000000000000000;
		47404: Delta = 69'sb000000000000000000000000000000000000000000000100000000000000000000000;
		3457: Delta = 69'sb111111111111111111111111111111111111111111111100000000000000000000000;
		43947: Delta = 69'sb000000000000000000000000000000000000000000001000000000000000000000000;
		6914: Delta = 69'sb111111111111111111111111111111111111111111111000000000000000000000000;
		37033: Delta = 69'sb000000000000000000000000000000000000000000010000000000000000000000000;
		13828: Delta = 69'sb111111111111111111111111111111111111111111110000000000000000000000000;
		23205: Delta = 69'sb000000000000000000000000000000000000000000100000000000000000000000000;
		27656: Delta = 69'sb111111111111111111111111111111111111111111100000000000000000000000000;
		46410: Delta = 69'sb000000000000000000000000000000000000000001000000000000000000000000000;
		4451: Delta = 69'sb111111111111111111111111111111111111111111000000000000000000000000000;
		41959: Delta = 69'sb000000000000000000000000000000000000000010000000000000000000000000000;
		8902: Delta = 69'sb111111111111111111111111111111111111111110000000000000000000000000000;
		33057: Delta = 69'sb000000000000000000000000000000000000000100000000000000000000000000000;
		17804: Delta = 69'sb111111111111111111111111111111111111111100000000000000000000000000000;
		15253: Delta = 69'sb000000000000000000000000000000000000001000000000000000000000000000000;
		35608: Delta = 69'sb111111111111111111111111111111111111111000000000000000000000000000000;
		30506: Delta = 69'sb000000000000000000000000000000000000010000000000000000000000000000000;
		20355: Delta = 69'sb111111111111111111111111111111111111110000000000000000000000000000000;
		10151: Delta = 69'sb000000000000000000000000000000000000100000000000000000000000000000000;
		40710: Delta = 69'sb111111111111111111111111111111111111100000000000000000000000000000000;
		20302: Delta = 69'sb000000000000000000000000000000000001000000000000000000000000000000000;
		30559: Delta = 69'sb111111111111111111111111111111111111000000000000000000000000000000000;
		40604: Delta = 69'sb000000000000000000000000000000000010000000000000000000000000000000000;
		10257: Delta = 69'sb111111111111111111111111111111111110000000000000000000000000000000000;
		30347: Delta = 69'sb000000000000000000000000000000000100000000000000000000000000000000000;
		20514: Delta = 69'sb111111111111111111111111111111111100000000000000000000000000000000000;
		9833: Delta = 69'sb000000000000000000000000000000001000000000000000000000000000000000000;
		41028: Delta = 69'sb111111111111111111111111111111111000000000000000000000000000000000000;
		19666: Delta = 69'sb000000000000000000000000000000010000000000000000000000000000000000000;
		31195: Delta = 69'sb111111111111111111111111111111110000000000000000000000000000000000000;
		39332: Delta = 69'sb000000000000000000000000000000100000000000000000000000000000000000000;
		11529: Delta = 69'sb111111111111111111111111111111100000000000000000000000000000000000000;
		27803: Delta = 69'sb000000000000000000000000000001000000000000000000000000000000000000000;
		23058: Delta = 69'sb111111111111111111111111111111000000000000000000000000000000000000000;
		4745: Delta = 69'sb000000000000000000000000000010000000000000000000000000000000000000000;
		46116: Delta = 69'sb111111111111111111111111111110000000000000000000000000000000000000000;
		9490: Delta = 69'sb000000000000000000000000000100000000000000000000000000000000000000000;
		41371: Delta = 69'sb111111111111111111111111111100000000000000000000000000000000000000000;
		18980: Delta = 69'sb000000000000000000000000001000000000000000000000000000000000000000000;
		31881: Delta = 69'sb111111111111111111111111111000000000000000000000000000000000000000000;
		37960: Delta = 69'sb000000000000000000000000010000000000000000000000000000000000000000000;
		12901: Delta = 69'sb111111111111111111111111110000000000000000000000000000000000000000000;
		25059: Delta = 69'sb000000000000000000000000100000000000000000000000000000000000000000000;
		25802: Delta = 69'sb111111111111111111111111100000000000000000000000000000000000000000000;
		50118: Delta = 69'sb000000000000000000000001000000000000000000000000000000000000000000000;
		743: Delta = 69'sb111111111111111111111111000000000000000000000000000000000000000000000;
		49375: Delta = 69'sb000000000000000000000010000000000000000000000000000000000000000000000;
		1486: Delta = 69'sb111111111111111111111110000000000000000000000000000000000000000000000;
		47889: Delta = 69'sb000000000000000000000100000000000000000000000000000000000000000000000;
		2972: Delta = 69'sb111111111111111111111100000000000000000000000000000000000000000000000;
		44917: Delta = 69'sb000000000000000000001000000000000000000000000000000000000000000000000;
		5944: Delta = 69'sb111111111111111111111000000000000000000000000000000000000000000000000;
		38973: Delta = 69'sb000000000000000000010000000000000000000000000000000000000000000000000;
		11888: Delta = 69'sb111111111111111111110000000000000000000000000000000000000000000000000;
		27085: Delta = 69'sb000000000000000000100000000000000000000000000000000000000000000000000;
		23776: Delta = 69'sb111111111111111111100000000000000000000000000000000000000000000000000;
		3309: Delta = 69'sb000000000000000001000000000000000000000000000000000000000000000000000;
		47552: Delta = 69'sb111111111111111111000000000000000000000000000000000000000000000000000;
		6618: Delta = 69'sb000000000000000010000000000000000000000000000000000000000000000000000;
		44243: Delta = 69'sb111111111111111110000000000000000000000000000000000000000000000000000;
		13236: Delta = 69'sb000000000000000100000000000000000000000000000000000000000000000000000;
		37625: Delta = 69'sb111111111111111100000000000000000000000000000000000000000000000000000;
		26472: Delta = 69'sb000000000000001000000000000000000000000000000000000000000000000000000;
		24389: Delta = 69'sb111111111111111000000000000000000000000000000000000000000000000000000;
		2083: Delta = 69'sb000000000000010000000000000000000000000000000000000000000000000000000;
		48778: Delta = 69'sb111111111111110000000000000000000000000000000000000000000000000000000;
		4166: Delta = 69'sb000000000000100000000000000000000000000000000000000000000000000000000;
		46695: Delta = 69'sb111111111111100000000000000000000000000000000000000000000000000000000;
		8332: Delta = 69'sb000000000001000000000000000000000000000000000000000000000000000000000;
		42529: Delta = 69'sb111111111111000000000000000000000000000000000000000000000000000000000;
		16664: Delta = 69'sb000000000010000000000000000000000000000000000000000000000000000000000;
		34197: Delta = 69'sb111111111110000000000000000000000000000000000000000000000000000000000;
		33328: Delta = 69'sb000000000100000000000000000000000000000000000000000000000000000000000;
		17533: Delta = 69'sb111111111100000000000000000000000000000000000000000000000000000000000;
		15795: Delta = 69'sb000000001000000000000000000000000000000000000000000000000000000000000;
		35066: Delta = 69'sb111111111000000000000000000000000000000000000000000000000000000000000;
		31590: Delta = 69'sb000000010000000000000000000000000000000000000000000000000000000000000;
		19271: Delta = 69'sb111111110000000000000000000000000000000000000000000000000000000000000;
		12319: Delta = 69'sb000000100000000000000000000000000000000000000000000000000000000000000;
		38542: Delta = 69'sb111111100000000000000000000000000000000000000000000000000000000000000;
		24638: Delta = 69'sb000001000000000000000000000000000000000000000000000000000000000000000;
		26223: Delta = 69'sb111111000000000000000000000000000000000000000000000000000000000000000;
		49276: Delta = 69'sb000010000000000000000000000000000000000000000000000000000000000000000;
		1585: Delta = 69'sb111110000000000000000000000000000000000000000000000000000000000000000;
		47691: Delta = 69'sb000100000000000000000000000000000000000000000000000000000000000000000;
		3170: Delta = 69'sb111100000000000000000000000000000000000000000000000000000000000000000;
		44521: Delta = 69'sb001000000000000000000000000000000000000000000000000000000000000000000;
		6340: Delta = 69'sb111000000000000000000000000000000000000000000000000000000000000000000;
		38181: Delta = 69'sb010000000000000000000000000000000000000000000000000000000000000000000;
		12680: Delta = 69'sb110000000000000000000000000000000000000000000000000000000000000000000;
		3: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000000011;
		50858: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111111101;
		5: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000000101;
		50856: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111111011;
		9: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000001001;
		50854: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111111001;
		7: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000000111;
		50852: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111110111;
		17: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000010001;
		50846: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111110001;
		15: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000001111;
		50844: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111101111;
		33: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000100001;
		50830: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111100001;
		31: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000011111;
		50828: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111011111;
		65: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000001000001;
		50798: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111000001;
		63: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000111111;
		50796: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111110111111;
		129: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000010000001;
		50734: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111110000001;
		127: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000001111111;
		50732: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111101111111;
		257: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000100000001;
		50606: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111100000001;
		255: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000011111111;
		50604: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111011111111;
		513: Delta = 69'sb000000000000000000000000000000000000000000000000000000000001000000001;
		50350: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111000000001;
		511: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000111111111;
		50348: Delta = 69'sb111111111111111111111111111111111111111111111111111111111110111111111;
		1025: Delta = 69'sb000000000000000000000000000000000000000000000000000000000010000000001;
		49838: Delta = 69'sb111111111111111111111111111111111111111111111111111111111110000000001;
		1023: Delta = 69'sb000000000000000000000000000000000000000000000000000000000001111111111;
		49836: Delta = 69'sb111111111111111111111111111111111111111111111111111111111101111111111;
		2049: Delta = 69'sb000000000000000000000000000000000000000000000000000000000100000000001;
		48814: Delta = 69'sb111111111111111111111111111111111111111111111111111111111100000000001;
		2047: Delta = 69'sb000000000000000000000000000000000000000000000000000000000011111111111;
		48812: Delta = 69'sb111111111111111111111111111111111111111111111111111111111011111111111;
		4097: Delta = 69'sb000000000000000000000000000000000000000000000000000000001000000000001;
		46766: Delta = 69'sb111111111111111111111111111111111111111111111111111111111000000000001;
		4095: Delta = 69'sb000000000000000000000000000000000000000000000000000000000111111111111;
		46764: Delta = 69'sb111111111111111111111111111111111111111111111111111111110111111111111;
		8193: Delta = 69'sb000000000000000000000000000000000000000000000000000000010000000000001;
		42670: Delta = 69'sb111111111111111111111111111111111111111111111111111111110000000000001;
		8191: Delta = 69'sb000000000000000000000000000000000000000000000000000000001111111111111;
		42668: Delta = 69'sb111111111111111111111111111111111111111111111111111111101111111111111;
		16385: Delta = 69'sb000000000000000000000000000000000000000000000000000000100000000000001;
		34478: Delta = 69'sb111111111111111111111111111111111111111111111111111111100000000000001;
		16383: Delta = 69'sb000000000000000000000000000000000000000000000000000000011111111111111;
		34476: Delta = 69'sb111111111111111111111111111111111111111111111111111111011111111111111;
		32769: Delta = 69'sb000000000000000000000000000000000000000000000000000001000000000000001;
		18094: Delta = 69'sb111111111111111111111111111111111111111111111111111111000000000000001;
		32767: Delta = 69'sb000000000000000000000000000000000000000000000000000000111111111111111;
		18092: Delta = 69'sb111111111111111111111111111111111111111111111111111110111111111111111;
		14676: Delta = 69'sb000000000000000000000000000000000000000000000000000010000000000000001;
		36187: Delta = 69'sb111111111111111111111111111111111111111111111111111110000000000000001;
		14674: Delta = 69'sb000000000000000000000000000000000000000000000000000001111111111111111;
		36185: Delta = 69'sb111111111111111111111111111111111111111111111111111101111111111111111;
		29351: Delta = 69'sb000000000000000000000000000000000000000000000000000100000000000000001;
		21512: Delta = 69'sb111111111111111111111111111111111111111111111111111100000000000000001;
		29349: Delta = 69'sb000000000000000000000000000000000000000000000000000011111111111111111;
		21510: Delta = 69'sb111111111111111111111111111111111111111111111111111011111111111111111;
		7840: Delta = 69'sb000000000000000000000000000000000000000000000000001000000000000000001;
		43023: Delta = 69'sb111111111111111111111111111111111111111111111111111000000000000000001;
		7838: Delta = 69'sb000000000000000000000000000000000000000000000000000111111111111111111;
		43021: Delta = 69'sb111111111111111111111111111111111111111111111111110111111111111111111;
		15679: Delta = 69'sb000000000000000000000000000000000000000000000000010000000000000000001;
		35184: Delta = 69'sb111111111111111111111111111111111111111111111111110000000000000000001;
		15677: Delta = 69'sb000000000000000000000000000000000000000000000000001111111111111111111;
		35182: Delta = 69'sb111111111111111111111111111111111111111111111111101111111111111111111;
		31357: Delta = 69'sb000000000000000000000000000000000000000000000000100000000000000000001;
		19506: Delta = 69'sb111111111111111111111111111111111111111111111111100000000000000000001;
		31355: Delta = 69'sb000000000000000000000000000000000000000000000000011111111111111111111;
		19504: Delta = 69'sb111111111111111111111111111111111111111111111111011111111111111111111;
		11852: Delta = 69'sb000000000000000000000000000000000000000000000001000000000000000000001;
		39011: Delta = 69'sb111111111111111111111111111111111111111111111111000000000000000000001;
		11850: Delta = 69'sb000000000000000000000000000000000000000000000000111111111111111111111;
		39009: Delta = 69'sb111111111111111111111111111111111111111111111110111111111111111111111;
		23703: Delta = 69'sb000000000000000000000000000000000000000000000010000000000000000000001;
		27160: Delta = 69'sb111111111111111111111111111111111111111111111110000000000000000000001;
		23701: Delta = 69'sb000000000000000000000000000000000000000000000001111111111111111111111;
		27158: Delta = 69'sb111111111111111111111111111111111111111111111101111111111111111111111;
		47405: Delta = 69'sb000000000000000000000000000000000000000000000100000000000000000000001;
		3458: Delta = 69'sb111111111111111111111111111111111111111111111100000000000000000000001;
		47403: Delta = 69'sb000000000000000000000000000000000000000000000011111111111111111111111;
		3456: Delta = 69'sb111111111111111111111111111111111111111111111011111111111111111111111;
		43948: Delta = 69'sb000000000000000000000000000000000000000000001000000000000000000000001;
		6915: Delta = 69'sb111111111111111111111111111111111111111111111000000000000000000000001;
		43946: Delta = 69'sb000000000000000000000000000000000000000000000111111111111111111111111;
		6913: Delta = 69'sb111111111111111111111111111111111111111111110111111111111111111111111;
		37034: Delta = 69'sb000000000000000000000000000000000000000000010000000000000000000000001;
		13829: Delta = 69'sb111111111111111111111111111111111111111111110000000000000000000000001;
		37032: Delta = 69'sb000000000000000000000000000000000000000000001111111111111111111111111;
		13827: Delta = 69'sb111111111111111111111111111111111111111111101111111111111111111111111;
		23206: Delta = 69'sb000000000000000000000000000000000000000000100000000000000000000000001;
		27657: Delta = 69'sb111111111111111111111111111111111111111111100000000000000000000000001;
		23204: Delta = 69'sb000000000000000000000000000000000000000000011111111111111111111111111;
		27655: Delta = 69'sb111111111111111111111111111111111111111111011111111111111111111111111;
		46411: Delta = 69'sb000000000000000000000000000000000000000001000000000000000000000000001;
		4452: Delta = 69'sb111111111111111111111111111111111111111111000000000000000000000000001;
		46409: Delta = 69'sb000000000000000000000000000000000000000000111111111111111111111111111;
		4450: Delta = 69'sb111111111111111111111111111111111111111110111111111111111111111111111;
		41960: Delta = 69'sb000000000000000000000000000000000000000010000000000000000000000000001;
		8903: Delta = 69'sb111111111111111111111111111111111111111110000000000000000000000000001;
		41958: Delta = 69'sb000000000000000000000000000000000000000001111111111111111111111111111;
		8901: Delta = 69'sb111111111111111111111111111111111111111101111111111111111111111111111;
		33058: Delta = 69'sb000000000000000000000000000000000000000100000000000000000000000000001;
		17805: Delta = 69'sb111111111111111111111111111111111111111100000000000000000000000000001;
		33056: Delta = 69'sb000000000000000000000000000000000000000011111111111111111111111111111;
		17803: Delta = 69'sb111111111111111111111111111111111111111011111111111111111111111111111;
		15254: Delta = 69'sb000000000000000000000000000000000000001000000000000000000000000000001;
		35609: Delta = 69'sb111111111111111111111111111111111111111000000000000000000000000000001;
		15252: Delta = 69'sb000000000000000000000000000000000000000111111111111111111111111111111;
		35607: Delta = 69'sb111111111111111111111111111111111111110111111111111111111111111111111;
		30507: Delta = 69'sb000000000000000000000000000000000000010000000000000000000000000000001;
		20356: Delta = 69'sb111111111111111111111111111111111111110000000000000000000000000000001;
		30505: Delta = 69'sb000000000000000000000000000000000000001111111111111111111111111111111;
		20354: Delta = 69'sb111111111111111111111111111111111111101111111111111111111111111111111;
		10152: Delta = 69'sb000000000000000000000000000000000000100000000000000000000000000000001;
		40711: Delta = 69'sb111111111111111111111111111111111111100000000000000000000000000000001;
		10150: Delta = 69'sb000000000000000000000000000000000000011111111111111111111111111111111;
		40709: Delta = 69'sb111111111111111111111111111111111111011111111111111111111111111111111;
		20303: Delta = 69'sb000000000000000000000000000000000001000000000000000000000000000000001;
		30560: Delta = 69'sb111111111111111111111111111111111111000000000000000000000000000000001;
		20301: Delta = 69'sb000000000000000000000000000000000000111111111111111111111111111111111;
		30558: Delta = 69'sb111111111111111111111111111111111110111111111111111111111111111111111;
		40605: Delta = 69'sb000000000000000000000000000000000010000000000000000000000000000000001;
		10258: Delta = 69'sb111111111111111111111111111111111110000000000000000000000000000000001;
		40603: Delta = 69'sb000000000000000000000000000000000001111111111111111111111111111111111;
		10256: Delta = 69'sb111111111111111111111111111111111101111111111111111111111111111111111;
		30348: Delta = 69'sb000000000000000000000000000000000100000000000000000000000000000000001;
		20515: Delta = 69'sb111111111111111111111111111111111100000000000000000000000000000000001;
		30346: Delta = 69'sb000000000000000000000000000000000011111111111111111111111111111111111;
		20513: Delta = 69'sb111111111111111111111111111111111011111111111111111111111111111111111;
		9834: Delta = 69'sb000000000000000000000000000000001000000000000000000000000000000000001;
		41029: Delta = 69'sb111111111111111111111111111111111000000000000000000000000000000000001;
		9832: Delta = 69'sb000000000000000000000000000000000111111111111111111111111111111111111;
		41027: Delta = 69'sb111111111111111111111111111111110111111111111111111111111111111111111;
		19667: Delta = 69'sb000000000000000000000000000000010000000000000000000000000000000000001;
		31196: Delta = 69'sb111111111111111111111111111111110000000000000000000000000000000000001;
		19665: Delta = 69'sb000000000000000000000000000000001111111111111111111111111111111111111;
		31194: Delta = 69'sb111111111111111111111111111111101111111111111111111111111111111111111;
		39333: Delta = 69'sb000000000000000000000000000000100000000000000000000000000000000000001;
		11530: Delta = 69'sb111111111111111111111111111111100000000000000000000000000000000000001;
		39331: Delta = 69'sb000000000000000000000000000000011111111111111111111111111111111111111;
		11528: Delta = 69'sb111111111111111111111111111111011111111111111111111111111111111111111;
		27804: Delta = 69'sb000000000000000000000000000001000000000000000000000000000000000000001;
		23059: Delta = 69'sb111111111111111111111111111111000000000000000000000000000000000000001;
		27802: Delta = 69'sb000000000000000000000000000000111111111111111111111111111111111111111;
		23057: Delta = 69'sb111111111111111111111111111110111111111111111111111111111111111111111;
		4746: Delta = 69'sb000000000000000000000000000010000000000000000000000000000000000000001;
		46117: Delta = 69'sb111111111111111111111111111110000000000000000000000000000000000000001;
		4744: Delta = 69'sb000000000000000000000000000001111111111111111111111111111111111111111;
		46115: Delta = 69'sb111111111111111111111111111101111111111111111111111111111111111111111;
		9491: Delta = 69'sb000000000000000000000000000100000000000000000000000000000000000000001;
		41372: Delta = 69'sb111111111111111111111111111100000000000000000000000000000000000000001;
		9489: Delta = 69'sb000000000000000000000000000011111111111111111111111111111111111111111;
		41370: Delta = 69'sb111111111111111111111111111011111111111111111111111111111111111111111;
		18981: Delta = 69'sb000000000000000000000000001000000000000000000000000000000000000000001;
		31882: Delta = 69'sb111111111111111111111111111000000000000000000000000000000000000000001;
		18979: Delta = 69'sb000000000000000000000000000111111111111111111111111111111111111111111;
		31880: Delta = 69'sb111111111111111111111111110111111111111111111111111111111111111111111;
		37961: Delta = 69'sb000000000000000000000000010000000000000000000000000000000000000000001;
		12902: Delta = 69'sb111111111111111111111111110000000000000000000000000000000000000000001;
		37959: Delta = 69'sb000000000000000000000000001111111111111111111111111111111111111111111;
		12900: Delta = 69'sb111111111111111111111111101111111111111111111111111111111111111111111;
		25060: Delta = 69'sb000000000000000000000000100000000000000000000000000000000000000000001;
		25803: Delta = 69'sb111111111111111111111111100000000000000000000000000000000000000000001;
		25058: Delta = 69'sb000000000000000000000000011111111111111111111111111111111111111111111;
		25801: Delta = 69'sb111111111111111111111111011111111111111111111111111111111111111111111;
		50119: Delta = 69'sb000000000000000000000001000000000000000000000000000000000000000000001;
		744: Delta = 69'sb111111111111111111111111000000000000000000000000000000000000000000001;
		50117: Delta = 69'sb000000000000000000000000111111111111111111111111111111111111111111111;
		742: Delta = 69'sb111111111111111111111110111111111111111111111111111111111111111111111;
		49376: Delta = 69'sb000000000000000000000010000000000000000000000000000000000000000000001;
		1487: Delta = 69'sb111111111111111111111110000000000000000000000000000000000000000000001;
		49374: Delta = 69'sb000000000000000000000001111111111111111111111111111111111111111111111;
		1485: Delta = 69'sb111111111111111111111101111111111111111111111111111111111111111111111;
		47890: Delta = 69'sb000000000000000000000100000000000000000000000000000000000000000000001;
		2973: Delta = 69'sb111111111111111111111100000000000000000000000000000000000000000000001;
		47888: Delta = 69'sb000000000000000000000011111111111111111111111111111111111111111111111;
		2971: Delta = 69'sb111111111111111111111011111111111111111111111111111111111111111111111;
		44918: Delta = 69'sb000000000000000000001000000000000000000000000000000000000000000000001;
		5945: Delta = 69'sb111111111111111111111000000000000000000000000000000000000000000000001;
		44916: Delta = 69'sb000000000000000000000111111111111111111111111111111111111111111111111;
		5943: Delta = 69'sb111111111111111111110111111111111111111111111111111111111111111111111;
		38974: Delta = 69'sb000000000000000000010000000000000000000000000000000000000000000000001;
		11889: Delta = 69'sb111111111111111111110000000000000000000000000000000000000000000000001;
		38972: Delta = 69'sb000000000000000000001111111111111111111111111111111111111111111111111;
		11887: Delta = 69'sb111111111111111111101111111111111111111111111111111111111111111111111;
		27086: Delta = 69'sb000000000000000000100000000000000000000000000000000000000000000000001;
		23777: Delta = 69'sb111111111111111111100000000000000000000000000000000000000000000000001;
		27084: Delta = 69'sb000000000000000000011111111111111111111111111111111111111111111111111;
		23775: Delta = 69'sb111111111111111111011111111111111111111111111111111111111111111111111;
		3310: Delta = 69'sb000000000000000001000000000000000000000000000000000000000000000000001;
		47553: Delta = 69'sb111111111111111111000000000000000000000000000000000000000000000000001;
		3308: Delta = 69'sb000000000000000000111111111111111111111111111111111111111111111111111;
		47551: Delta = 69'sb111111111111111110111111111111111111111111111111111111111111111111111;
		6619: Delta = 69'sb000000000000000010000000000000000000000000000000000000000000000000001;
		44244: Delta = 69'sb111111111111111110000000000000000000000000000000000000000000000000001;
		6617: Delta = 69'sb000000000000000001111111111111111111111111111111111111111111111111111;
		44242: Delta = 69'sb111111111111111101111111111111111111111111111111111111111111111111111;
		13237: Delta = 69'sb000000000000000100000000000000000000000000000000000000000000000000001;
		37626: Delta = 69'sb111111111111111100000000000000000000000000000000000000000000000000001;
		13235: Delta = 69'sb000000000000000011111111111111111111111111111111111111111111111111111;
		37624: Delta = 69'sb111111111111111011111111111111111111111111111111111111111111111111111;
		26473: Delta = 69'sb000000000000001000000000000000000000000000000000000000000000000000001;
		24390: Delta = 69'sb111111111111111000000000000000000000000000000000000000000000000000001;
		26471: Delta = 69'sb000000000000000111111111111111111111111111111111111111111111111111111;
		24388: Delta = 69'sb111111111111110111111111111111111111111111111111111111111111111111111;
		2084: Delta = 69'sb000000000000010000000000000000000000000000000000000000000000000000001;
		48779: Delta = 69'sb111111111111110000000000000000000000000000000000000000000000000000001;
		2082: Delta = 69'sb000000000000001111111111111111111111111111111111111111111111111111111;
		48777: Delta = 69'sb111111111111101111111111111111111111111111111111111111111111111111111;
		4167: Delta = 69'sb000000000000100000000000000000000000000000000000000000000000000000001;
		46696: Delta = 69'sb111111111111100000000000000000000000000000000000000000000000000000001;
		4165: Delta = 69'sb000000000000011111111111111111111111111111111111111111111111111111111;
		46694: Delta = 69'sb111111111111011111111111111111111111111111111111111111111111111111111;
		8333: Delta = 69'sb000000000001000000000000000000000000000000000000000000000000000000001;
		42530: Delta = 69'sb111111111111000000000000000000000000000000000000000000000000000000001;
		8331: Delta = 69'sb000000000000111111111111111111111111111111111111111111111111111111111;
		42528: Delta = 69'sb111111111110111111111111111111111111111111111111111111111111111111111;
		16665: Delta = 69'sb000000000010000000000000000000000000000000000000000000000000000000001;
		34198: Delta = 69'sb111111111110000000000000000000000000000000000000000000000000000000001;
		16663: Delta = 69'sb000000000001111111111111111111111111111111111111111111111111111111111;
		34196: Delta = 69'sb111111111101111111111111111111111111111111111111111111111111111111111;
		33329: Delta = 69'sb000000000100000000000000000000000000000000000000000000000000000000001;
		17534: Delta = 69'sb111111111100000000000000000000000000000000000000000000000000000000001;
		33327: Delta = 69'sb000000000011111111111111111111111111111111111111111111111111111111111;
		17532: Delta = 69'sb111111111011111111111111111111111111111111111111111111111111111111111;
		15796: Delta = 69'sb000000001000000000000000000000000000000000000000000000000000000000001;
		35067: Delta = 69'sb111111111000000000000000000000000000000000000000000000000000000000001;
		15794: Delta = 69'sb000000000111111111111111111111111111111111111111111111111111111111111;
		35065: Delta = 69'sb111111110111111111111111111111111111111111111111111111111111111111111;
		31591: Delta = 69'sb000000010000000000000000000000000000000000000000000000000000000000001;
		19272: Delta = 69'sb111111110000000000000000000000000000000000000000000000000000000000001;
		31589: Delta = 69'sb000000001111111111111111111111111111111111111111111111111111111111111;
		19270: Delta = 69'sb111111101111111111111111111111111111111111111111111111111111111111111;
		12320: Delta = 69'sb000000100000000000000000000000000000000000000000000000000000000000001;
		38543: Delta = 69'sb111111100000000000000000000000000000000000000000000000000000000000001;
		12318: Delta = 69'sb000000011111111111111111111111111111111111111111111111111111111111111;
		38541: Delta = 69'sb111111011111111111111111111111111111111111111111111111111111111111111;
		24639: Delta = 69'sb000001000000000000000000000000000000000000000000000000000000000000001;
		26224: Delta = 69'sb111111000000000000000000000000000000000000000000000000000000000000001;
		24637: Delta = 69'sb000000111111111111111111111111111111111111111111111111111111111111111;
		26222: Delta = 69'sb111110111111111111111111111111111111111111111111111111111111111111111;
		49277: Delta = 69'sb000010000000000000000000000000000000000000000000000000000000000000001;
		1586: Delta = 69'sb111110000000000000000000000000000000000000000000000000000000000000001;
		49275: Delta = 69'sb000001111111111111111111111111111111111111111111111111111111111111111;
		1584: Delta = 69'sb111101111111111111111111111111111111111111111111111111111111111111111;
		47692: Delta = 69'sb000100000000000000000000000000000000000000000000000000000000000000001;
		3171: Delta = 69'sb111100000000000000000000000000000000000000000000000000000000000000001;
		47690: Delta = 69'sb000011111111111111111111111111111111111111111111111111111111111111111;
		3169: Delta = 69'sb111011111111111111111111111111111111111111111111111111111111111111111;
		44522: Delta = 69'sb001000000000000000000000000000000000000000000000000000000000000000001;
		6341: Delta = 69'sb111000000000000000000000000000000000000000000000000000000000000000001;
		44520: Delta = 69'sb000111111111111111111111111111111111111111111111111111111111111111111;
		6339: Delta = 69'sb110111111111111111111111111111111111111111111111111111111111111111111;
		38182: Delta = 69'sb010000000000000000000000000000000000000000000000000000000000000000001;
		12681: Delta = 69'sb110000000000000000000000000000000000000000000000000000000000000000001;
		38180: Delta = 69'sb001111111111111111111111111111111111111111111111111111111111111111111;
		12679: Delta = 69'sb101111111111111111111111111111111111111111111111111111111111111111111;
		6: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000000110;
		50855: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111111010;
		10: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000001010;
		50851: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111110110;
		18: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000010010;
		50847: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111110010;
		14: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000001110;
		50843: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111101110;
		34: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000100010;
		50831: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111100010;
		30: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000011110;
		50827: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111011110;
		66: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000001000010;
		50799: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111000010;
		62: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000111110;
		50795: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111110111110;
		130: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000010000010;
		50735: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111110000010;
		126: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000001111110;
		50731: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111101111110;
		258: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000100000010;
		50607: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111100000010;
		254: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000011111110;
		50603: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111011111110;
		514: Delta = 69'sb000000000000000000000000000000000000000000000000000000000001000000010;
		50351: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111000000010;
		510: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000111111110;
		50347: Delta = 69'sb111111111111111111111111111111111111111111111111111111111110111111110;
		1026: Delta = 69'sb000000000000000000000000000000000000000000000000000000000010000000010;
		49839: Delta = 69'sb111111111111111111111111111111111111111111111111111111111110000000010;
		1022: Delta = 69'sb000000000000000000000000000000000000000000000000000000000001111111110;
		49835: Delta = 69'sb111111111111111111111111111111111111111111111111111111111101111111110;
		2050: Delta = 69'sb000000000000000000000000000000000000000000000000000000000100000000010;
		48815: Delta = 69'sb111111111111111111111111111111111111111111111111111111111100000000010;
		2046: Delta = 69'sb000000000000000000000000000000000000000000000000000000000011111111110;
		48811: Delta = 69'sb111111111111111111111111111111111111111111111111111111111011111111110;
		4098: Delta = 69'sb000000000000000000000000000000000000000000000000000000001000000000010;
		46767: Delta = 69'sb111111111111111111111111111111111111111111111111111111111000000000010;
		4094: Delta = 69'sb000000000000000000000000000000000000000000000000000000000111111111110;
		46763: Delta = 69'sb111111111111111111111111111111111111111111111111111111110111111111110;
		8194: Delta = 69'sb000000000000000000000000000000000000000000000000000000010000000000010;
		42671: Delta = 69'sb111111111111111111111111111111111111111111111111111111110000000000010;
		8190: Delta = 69'sb000000000000000000000000000000000000000000000000000000001111111111110;
		42667: Delta = 69'sb111111111111111111111111111111111111111111111111111111101111111111110;
		16386: Delta = 69'sb000000000000000000000000000000000000000000000000000000100000000000010;
		34479: Delta = 69'sb111111111111111111111111111111111111111111111111111111100000000000010;
		16382: Delta = 69'sb000000000000000000000000000000000000000000000000000000011111111111110;
		34475: Delta = 69'sb111111111111111111111111111111111111111111111111111111011111111111110;
		32770: Delta = 69'sb000000000000000000000000000000000000000000000000000001000000000000010;
		18095: Delta = 69'sb111111111111111111111111111111111111111111111111111111000000000000010;
		32766: Delta = 69'sb000000000000000000000000000000000000000000000000000000111111111111110;
		18091: Delta = 69'sb111111111111111111111111111111111111111111111111111110111111111111110;
		14677: Delta = 69'sb000000000000000000000000000000000000000000000000000010000000000000010;
		36188: Delta = 69'sb111111111111111111111111111111111111111111111111111110000000000000010;
		14673: Delta = 69'sb000000000000000000000000000000000000000000000000000001111111111111110;
		36184: Delta = 69'sb111111111111111111111111111111111111111111111111111101111111111111110;
		29352: Delta = 69'sb000000000000000000000000000000000000000000000000000100000000000000010;
		21513: Delta = 69'sb111111111111111111111111111111111111111111111111111100000000000000010;
		29348: Delta = 69'sb000000000000000000000000000000000000000000000000000011111111111111110;
		21509: Delta = 69'sb111111111111111111111111111111111111111111111111111011111111111111110;
		7841: Delta = 69'sb000000000000000000000000000000000000000000000000001000000000000000010;
		43024: Delta = 69'sb111111111111111111111111111111111111111111111111111000000000000000010;
		7837: Delta = 69'sb000000000000000000000000000000000000000000000000000111111111111111110;
		43020: Delta = 69'sb111111111111111111111111111111111111111111111111110111111111111111110;
		15680: Delta = 69'sb000000000000000000000000000000000000000000000000010000000000000000010;
		35185: Delta = 69'sb111111111111111111111111111111111111111111111111110000000000000000010;
		15676: Delta = 69'sb000000000000000000000000000000000000000000000000001111111111111111110;
		35181: Delta = 69'sb111111111111111111111111111111111111111111111111101111111111111111110;
		31358: Delta = 69'sb000000000000000000000000000000000000000000000000100000000000000000010;
		19507: Delta = 69'sb111111111111111111111111111111111111111111111111100000000000000000010;
		31354: Delta = 69'sb000000000000000000000000000000000000000000000000011111111111111111110;
		19503: Delta = 69'sb111111111111111111111111111111111111111111111111011111111111111111110;
		11853: Delta = 69'sb000000000000000000000000000000000000000000000001000000000000000000010;
		39012: Delta = 69'sb111111111111111111111111111111111111111111111111000000000000000000010;
		11849: Delta = 69'sb000000000000000000000000000000000000000000000000111111111111111111110;
		39008: Delta = 69'sb111111111111111111111111111111111111111111111110111111111111111111110;
		23704: Delta = 69'sb000000000000000000000000000000000000000000000010000000000000000000010;
		27161: Delta = 69'sb111111111111111111111111111111111111111111111110000000000000000000010;
		23700: Delta = 69'sb000000000000000000000000000000000000000000000001111111111111111111110;
		27157: Delta = 69'sb111111111111111111111111111111111111111111111101111111111111111111110;
		47406: Delta = 69'sb000000000000000000000000000000000000000000000100000000000000000000010;
		3459: Delta = 69'sb111111111111111111111111111111111111111111111100000000000000000000010;
		47402: Delta = 69'sb000000000000000000000000000000000000000000000011111111111111111111110;
		3455: Delta = 69'sb111111111111111111111111111111111111111111111011111111111111111111110;
		43949: Delta = 69'sb000000000000000000000000000000000000000000001000000000000000000000010;
		6916: Delta = 69'sb111111111111111111111111111111111111111111111000000000000000000000010;
		43945: Delta = 69'sb000000000000000000000000000000000000000000000111111111111111111111110;
		6912: Delta = 69'sb111111111111111111111111111111111111111111110111111111111111111111110;
		37035: Delta = 69'sb000000000000000000000000000000000000000000010000000000000000000000010;
		13830: Delta = 69'sb111111111111111111111111111111111111111111110000000000000000000000010;
		37031: Delta = 69'sb000000000000000000000000000000000000000000001111111111111111111111110;
		13826: Delta = 69'sb111111111111111111111111111111111111111111101111111111111111111111110;
		23207: Delta = 69'sb000000000000000000000000000000000000000000100000000000000000000000010;
		27658: Delta = 69'sb111111111111111111111111111111111111111111100000000000000000000000010;
		23203: Delta = 69'sb000000000000000000000000000000000000000000011111111111111111111111110;
		27654: Delta = 69'sb111111111111111111111111111111111111111111011111111111111111111111110;
		46412: Delta = 69'sb000000000000000000000000000000000000000001000000000000000000000000010;
		4453: Delta = 69'sb111111111111111111111111111111111111111111000000000000000000000000010;
		46408: Delta = 69'sb000000000000000000000000000000000000000000111111111111111111111111110;
		4449: Delta = 69'sb111111111111111111111111111111111111111110111111111111111111111111110;
		41961: Delta = 69'sb000000000000000000000000000000000000000010000000000000000000000000010;
		8904: Delta = 69'sb111111111111111111111111111111111111111110000000000000000000000000010;
		41957: Delta = 69'sb000000000000000000000000000000000000000001111111111111111111111111110;
		8900: Delta = 69'sb111111111111111111111111111111111111111101111111111111111111111111110;
		33059: Delta = 69'sb000000000000000000000000000000000000000100000000000000000000000000010;
		17806: Delta = 69'sb111111111111111111111111111111111111111100000000000000000000000000010;
		33055: Delta = 69'sb000000000000000000000000000000000000000011111111111111111111111111110;
		17802: Delta = 69'sb111111111111111111111111111111111111111011111111111111111111111111110;
		15255: Delta = 69'sb000000000000000000000000000000000000001000000000000000000000000000010;
		35610: Delta = 69'sb111111111111111111111111111111111111111000000000000000000000000000010;
		15251: Delta = 69'sb000000000000000000000000000000000000000111111111111111111111111111110;
		35606: Delta = 69'sb111111111111111111111111111111111111110111111111111111111111111111110;
		30508: Delta = 69'sb000000000000000000000000000000000000010000000000000000000000000000010;
		20357: Delta = 69'sb111111111111111111111111111111111111110000000000000000000000000000010;
		30504: Delta = 69'sb000000000000000000000000000000000000001111111111111111111111111111110;
		20353: Delta = 69'sb111111111111111111111111111111111111101111111111111111111111111111110;
		10153: Delta = 69'sb000000000000000000000000000000000000100000000000000000000000000000010;
		40712: Delta = 69'sb111111111111111111111111111111111111100000000000000000000000000000010;
		10149: Delta = 69'sb000000000000000000000000000000000000011111111111111111111111111111110;
		40708: Delta = 69'sb111111111111111111111111111111111111011111111111111111111111111111110;
		20304: Delta = 69'sb000000000000000000000000000000000001000000000000000000000000000000010;
		30561: Delta = 69'sb111111111111111111111111111111111111000000000000000000000000000000010;
		20300: Delta = 69'sb000000000000000000000000000000000000111111111111111111111111111111110;
		30557: Delta = 69'sb111111111111111111111111111111111110111111111111111111111111111111110;
		40606: Delta = 69'sb000000000000000000000000000000000010000000000000000000000000000000010;
		10259: Delta = 69'sb111111111111111111111111111111111110000000000000000000000000000000010;
		40602: Delta = 69'sb000000000000000000000000000000000001111111111111111111111111111111110;
		10255: Delta = 69'sb111111111111111111111111111111111101111111111111111111111111111111110;
		30349: Delta = 69'sb000000000000000000000000000000000100000000000000000000000000000000010;
		20516: Delta = 69'sb111111111111111111111111111111111100000000000000000000000000000000010;
		30345: Delta = 69'sb000000000000000000000000000000000011111111111111111111111111111111110;
		20512: Delta = 69'sb111111111111111111111111111111111011111111111111111111111111111111110;
		9835: Delta = 69'sb000000000000000000000000000000001000000000000000000000000000000000010;
		41030: Delta = 69'sb111111111111111111111111111111111000000000000000000000000000000000010;
		9831: Delta = 69'sb000000000000000000000000000000000111111111111111111111111111111111110;
		41026: Delta = 69'sb111111111111111111111111111111110111111111111111111111111111111111110;
		19668: Delta = 69'sb000000000000000000000000000000010000000000000000000000000000000000010;
		31197: Delta = 69'sb111111111111111111111111111111110000000000000000000000000000000000010;
		19664: Delta = 69'sb000000000000000000000000000000001111111111111111111111111111111111110;
		31193: Delta = 69'sb111111111111111111111111111111101111111111111111111111111111111111110;
		39334: Delta = 69'sb000000000000000000000000000000100000000000000000000000000000000000010;
		11531: Delta = 69'sb111111111111111111111111111111100000000000000000000000000000000000010;
		39330: Delta = 69'sb000000000000000000000000000000011111111111111111111111111111111111110;
		11527: Delta = 69'sb111111111111111111111111111111011111111111111111111111111111111111110;
		27805: Delta = 69'sb000000000000000000000000000001000000000000000000000000000000000000010;
		23060: Delta = 69'sb111111111111111111111111111111000000000000000000000000000000000000010;
		27801: Delta = 69'sb000000000000000000000000000000111111111111111111111111111111111111110;
		23056: Delta = 69'sb111111111111111111111111111110111111111111111111111111111111111111110;
		4747: Delta = 69'sb000000000000000000000000000010000000000000000000000000000000000000010;
		46118: Delta = 69'sb111111111111111111111111111110000000000000000000000000000000000000010;
		4743: Delta = 69'sb000000000000000000000000000001111111111111111111111111111111111111110;
		46114: Delta = 69'sb111111111111111111111111111101111111111111111111111111111111111111110;
		9492: Delta = 69'sb000000000000000000000000000100000000000000000000000000000000000000010;
		41373: Delta = 69'sb111111111111111111111111111100000000000000000000000000000000000000010;
		9488: Delta = 69'sb000000000000000000000000000011111111111111111111111111111111111111110;
		41369: Delta = 69'sb111111111111111111111111111011111111111111111111111111111111111111110;
		18982: Delta = 69'sb000000000000000000000000001000000000000000000000000000000000000000010;
		31883: Delta = 69'sb111111111111111111111111111000000000000000000000000000000000000000010;
		18978: Delta = 69'sb000000000000000000000000000111111111111111111111111111111111111111110;
		31879: Delta = 69'sb111111111111111111111111110111111111111111111111111111111111111111110;
		37962: Delta = 69'sb000000000000000000000000010000000000000000000000000000000000000000010;
		12903: Delta = 69'sb111111111111111111111111110000000000000000000000000000000000000000010;
		37958: Delta = 69'sb000000000000000000000000001111111111111111111111111111111111111111110;
		12899: Delta = 69'sb111111111111111111111111101111111111111111111111111111111111111111110;
		25061: Delta = 69'sb000000000000000000000000100000000000000000000000000000000000000000010;
		25804: Delta = 69'sb111111111111111111111111100000000000000000000000000000000000000000010;
		25057: Delta = 69'sb000000000000000000000000011111111111111111111111111111111111111111110;
		25800: Delta = 69'sb111111111111111111111111011111111111111111111111111111111111111111110;
		50120: Delta = 69'sb000000000000000000000001000000000000000000000000000000000000000000010;
		745: Delta = 69'sb111111111111111111111111000000000000000000000000000000000000000000010;
		50116: Delta = 69'sb000000000000000000000000111111111111111111111111111111111111111111110;
		741: Delta = 69'sb111111111111111111111110111111111111111111111111111111111111111111110;
		49377: Delta = 69'sb000000000000000000000010000000000000000000000000000000000000000000010;
		1488: Delta = 69'sb111111111111111111111110000000000000000000000000000000000000000000010;
		49373: Delta = 69'sb000000000000000000000001111111111111111111111111111111111111111111110;
		1484: Delta = 69'sb111111111111111111111101111111111111111111111111111111111111111111110;
		47891: Delta = 69'sb000000000000000000000100000000000000000000000000000000000000000000010;
		2974: Delta = 69'sb111111111111111111111100000000000000000000000000000000000000000000010;
		47887: Delta = 69'sb000000000000000000000011111111111111111111111111111111111111111111110;
		2970: Delta = 69'sb111111111111111111111011111111111111111111111111111111111111111111110;
		44919: Delta = 69'sb000000000000000000001000000000000000000000000000000000000000000000010;
		5946: Delta = 69'sb111111111111111111111000000000000000000000000000000000000000000000010;
		44915: Delta = 69'sb000000000000000000000111111111111111111111111111111111111111111111110;
		5942: Delta = 69'sb111111111111111111110111111111111111111111111111111111111111111111110;
		38975: Delta = 69'sb000000000000000000010000000000000000000000000000000000000000000000010;
		11890: Delta = 69'sb111111111111111111110000000000000000000000000000000000000000000000010;
		38971: Delta = 69'sb000000000000000000001111111111111111111111111111111111111111111111110;
		11886: Delta = 69'sb111111111111111111101111111111111111111111111111111111111111111111110;
		27087: Delta = 69'sb000000000000000000100000000000000000000000000000000000000000000000010;
		23778: Delta = 69'sb111111111111111111100000000000000000000000000000000000000000000000010;
		27083: Delta = 69'sb000000000000000000011111111111111111111111111111111111111111111111110;
		23774: Delta = 69'sb111111111111111111011111111111111111111111111111111111111111111111110;
		3311: Delta = 69'sb000000000000000001000000000000000000000000000000000000000000000000010;
		47554: Delta = 69'sb111111111111111111000000000000000000000000000000000000000000000000010;
		3307: Delta = 69'sb000000000000000000111111111111111111111111111111111111111111111111110;
		47550: Delta = 69'sb111111111111111110111111111111111111111111111111111111111111111111110;
		6620: Delta = 69'sb000000000000000010000000000000000000000000000000000000000000000000010;
		44245: Delta = 69'sb111111111111111110000000000000000000000000000000000000000000000000010;
		6616: Delta = 69'sb000000000000000001111111111111111111111111111111111111111111111111110;
		44241: Delta = 69'sb111111111111111101111111111111111111111111111111111111111111111111110;
		13238: Delta = 69'sb000000000000000100000000000000000000000000000000000000000000000000010;
		37627: Delta = 69'sb111111111111111100000000000000000000000000000000000000000000000000010;
		13234: Delta = 69'sb000000000000000011111111111111111111111111111111111111111111111111110;
		37623: Delta = 69'sb111111111111111011111111111111111111111111111111111111111111111111110;
		26474: Delta = 69'sb000000000000001000000000000000000000000000000000000000000000000000010;
		24391: Delta = 69'sb111111111111111000000000000000000000000000000000000000000000000000010;
		26470: Delta = 69'sb000000000000000111111111111111111111111111111111111111111111111111110;
		24387: Delta = 69'sb111111111111110111111111111111111111111111111111111111111111111111110;
		2085: Delta = 69'sb000000000000010000000000000000000000000000000000000000000000000000010;
		48780: Delta = 69'sb111111111111110000000000000000000000000000000000000000000000000000010;
		2081: Delta = 69'sb000000000000001111111111111111111111111111111111111111111111111111110;
		48776: Delta = 69'sb111111111111101111111111111111111111111111111111111111111111111111110;
		4168: Delta = 69'sb000000000000100000000000000000000000000000000000000000000000000000010;
		46697: Delta = 69'sb111111111111100000000000000000000000000000000000000000000000000000010;
		4164: Delta = 69'sb000000000000011111111111111111111111111111111111111111111111111111110;
		46693: Delta = 69'sb111111111111011111111111111111111111111111111111111111111111111111110;
		8334: Delta = 69'sb000000000001000000000000000000000000000000000000000000000000000000010;
		42531: Delta = 69'sb111111111111000000000000000000000000000000000000000000000000000000010;
		8330: Delta = 69'sb000000000000111111111111111111111111111111111111111111111111111111110;
		42527: Delta = 69'sb111111111110111111111111111111111111111111111111111111111111111111110;
		16666: Delta = 69'sb000000000010000000000000000000000000000000000000000000000000000000010;
		34199: Delta = 69'sb111111111110000000000000000000000000000000000000000000000000000000010;
		16662: Delta = 69'sb000000000001111111111111111111111111111111111111111111111111111111110;
		34195: Delta = 69'sb111111111101111111111111111111111111111111111111111111111111111111110;
		33330: Delta = 69'sb000000000100000000000000000000000000000000000000000000000000000000010;
		17535: Delta = 69'sb111111111100000000000000000000000000000000000000000000000000000000010;
		33326: Delta = 69'sb000000000011111111111111111111111111111111111111111111111111111111110;
		17531: Delta = 69'sb111111111011111111111111111111111111111111111111111111111111111111110;
		15797: Delta = 69'sb000000001000000000000000000000000000000000000000000000000000000000010;
		35068: Delta = 69'sb111111111000000000000000000000000000000000000000000000000000000000010;
		15793: Delta = 69'sb000000000111111111111111111111111111111111111111111111111111111111110;
		35064: Delta = 69'sb111111110111111111111111111111111111111111111111111111111111111111110;
		31592: Delta = 69'sb000000010000000000000000000000000000000000000000000000000000000000010;
		19273: Delta = 69'sb111111110000000000000000000000000000000000000000000000000000000000010;
		31588: Delta = 69'sb000000001111111111111111111111111111111111111111111111111111111111110;
		19269: Delta = 69'sb111111101111111111111111111111111111111111111111111111111111111111110;
		12321: Delta = 69'sb000000100000000000000000000000000000000000000000000000000000000000010;
		38544: Delta = 69'sb111111100000000000000000000000000000000000000000000000000000000000010;
		12317: Delta = 69'sb000000011111111111111111111111111111111111111111111111111111111111110;
		38540: Delta = 69'sb111111011111111111111111111111111111111111111111111111111111111111110;
		24640: Delta = 69'sb000001000000000000000000000000000000000000000000000000000000000000010;
		26225: Delta = 69'sb111111000000000000000000000000000000000000000000000000000000000000010;
		24636: Delta = 69'sb000000111111111111111111111111111111111111111111111111111111111111110;
		26221: Delta = 69'sb111110111111111111111111111111111111111111111111111111111111111111110;
		49278: Delta = 69'sb000010000000000000000000000000000000000000000000000000000000000000010;
		1587: Delta = 69'sb111110000000000000000000000000000000000000000000000000000000000000010;
		49274: Delta = 69'sb000001111111111111111111111111111111111111111111111111111111111111110;
		1583: Delta = 69'sb111101111111111111111111111111111111111111111111111111111111111111110;
		47693: Delta = 69'sb000100000000000000000000000000000000000000000000000000000000000000010;
		3172: Delta = 69'sb111100000000000000000000000000000000000000000000000000000000000000010;
		47689: Delta = 69'sb000011111111111111111111111111111111111111111111111111111111111111110;
		3168: Delta = 69'sb111011111111111111111111111111111111111111111111111111111111111111110;
		44523: Delta = 69'sb001000000000000000000000000000000000000000000000000000000000000000010;
		6342: Delta = 69'sb111000000000000000000000000000000000000000000000000000000000000000010;
		44519: Delta = 69'sb000111111111111111111111111111111111111111111111111111111111111111110;
		6338: Delta = 69'sb110111111111111111111111111111111111111111111111111111111111111111110;
		38183: Delta = 69'sb010000000000000000000000000000000000000000000000000000000000000000010;
		12682: Delta = 69'sb110000000000000000000000000000000000000000000000000000000000000000010;
		38179: Delta = 69'sb001111111111111111111111111111111111111111111111111111111111111111110;
		12678: Delta = 69'sb101111111111111111111111111111111111111111111111111111111111111111110;
		12: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000001100;
		50849: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111110100;
		20: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000010100;
		50841: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111101100;
		36: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000100100;
		50833: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111100100;
		28: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000011100;
		50825: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111011100;
		68: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000001000100;
		50801: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111000100;
		60: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000111100;
		50793: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111110111100;
		132: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000010000100;
		50737: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111110000100;
		124: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000001111100;
		50729: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111101111100;
		260: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000100000100;
		50609: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111100000100;
		252: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000011111100;
		50601: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111011111100;
		516: Delta = 69'sb000000000000000000000000000000000000000000000000000000000001000000100;
		50353: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111000000100;
		508: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000111111100;
		50345: Delta = 69'sb111111111111111111111111111111111111111111111111111111111110111111100;
		1028: Delta = 69'sb000000000000000000000000000000000000000000000000000000000010000000100;
		49841: Delta = 69'sb111111111111111111111111111111111111111111111111111111111110000000100;
		1020: Delta = 69'sb000000000000000000000000000000000000000000000000000000000001111111100;
		49833: Delta = 69'sb111111111111111111111111111111111111111111111111111111111101111111100;
		2052: Delta = 69'sb000000000000000000000000000000000000000000000000000000000100000000100;
		48817: Delta = 69'sb111111111111111111111111111111111111111111111111111111111100000000100;
		2044: Delta = 69'sb000000000000000000000000000000000000000000000000000000000011111111100;
		48809: Delta = 69'sb111111111111111111111111111111111111111111111111111111111011111111100;
		4100: Delta = 69'sb000000000000000000000000000000000000000000000000000000001000000000100;
		46769: Delta = 69'sb111111111111111111111111111111111111111111111111111111111000000000100;
		4092: Delta = 69'sb000000000000000000000000000000000000000000000000000000000111111111100;
		46761: Delta = 69'sb111111111111111111111111111111111111111111111111111111110111111111100;
		8196: Delta = 69'sb000000000000000000000000000000000000000000000000000000010000000000100;
		42673: Delta = 69'sb111111111111111111111111111111111111111111111111111111110000000000100;
		8188: Delta = 69'sb000000000000000000000000000000000000000000000000000000001111111111100;
		42665: Delta = 69'sb111111111111111111111111111111111111111111111111111111101111111111100;
		16388: Delta = 69'sb000000000000000000000000000000000000000000000000000000100000000000100;
		34481: Delta = 69'sb111111111111111111111111111111111111111111111111111111100000000000100;
		16380: Delta = 69'sb000000000000000000000000000000000000000000000000000000011111111111100;
		34473: Delta = 69'sb111111111111111111111111111111111111111111111111111111011111111111100;
		32772: Delta = 69'sb000000000000000000000000000000000000000000000000000001000000000000100;
		18097: Delta = 69'sb111111111111111111111111111111111111111111111111111111000000000000100;
		32764: Delta = 69'sb000000000000000000000000000000000000000000000000000000111111111111100;
		18089: Delta = 69'sb111111111111111111111111111111111111111111111111111110111111111111100;
		14679: Delta = 69'sb000000000000000000000000000000000000000000000000000010000000000000100;
		36190: Delta = 69'sb111111111111111111111111111111111111111111111111111110000000000000100;
		14671: Delta = 69'sb000000000000000000000000000000000000000000000000000001111111111111100;
		36182: Delta = 69'sb111111111111111111111111111111111111111111111111111101111111111111100;
		29354: Delta = 69'sb000000000000000000000000000000000000000000000000000100000000000000100;
		21515: Delta = 69'sb111111111111111111111111111111111111111111111111111100000000000000100;
		29346: Delta = 69'sb000000000000000000000000000000000000000000000000000011111111111111100;
		21507: Delta = 69'sb111111111111111111111111111111111111111111111111111011111111111111100;
		7843: Delta = 69'sb000000000000000000000000000000000000000000000000001000000000000000100;
		43026: Delta = 69'sb111111111111111111111111111111111111111111111111111000000000000000100;
		7835: Delta = 69'sb000000000000000000000000000000000000000000000000000111111111111111100;
		43018: Delta = 69'sb111111111111111111111111111111111111111111111111110111111111111111100;
		15682: Delta = 69'sb000000000000000000000000000000000000000000000000010000000000000000100;
		35187: Delta = 69'sb111111111111111111111111111111111111111111111111110000000000000000100;
		15674: Delta = 69'sb000000000000000000000000000000000000000000000000001111111111111111100;
		35179: Delta = 69'sb111111111111111111111111111111111111111111111111101111111111111111100;
		31360: Delta = 69'sb000000000000000000000000000000000000000000000000100000000000000000100;
		19509: Delta = 69'sb111111111111111111111111111111111111111111111111100000000000000000100;
		31352: Delta = 69'sb000000000000000000000000000000000000000000000000011111111111111111100;
		19501: Delta = 69'sb111111111111111111111111111111111111111111111111011111111111111111100;
		11855: Delta = 69'sb000000000000000000000000000000000000000000000001000000000000000000100;
		39014: Delta = 69'sb111111111111111111111111111111111111111111111111000000000000000000100;
		11847: Delta = 69'sb000000000000000000000000000000000000000000000000111111111111111111100;
		39006: Delta = 69'sb111111111111111111111111111111111111111111111110111111111111111111100;
		23706: Delta = 69'sb000000000000000000000000000000000000000000000010000000000000000000100;
		27163: Delta = 69'sb111111111111111111111111111111111111111111111110000000000000000000100;
		23698: Delta = 69'sb000000000000000000000000000000000000000000000001111111111111111111100;
		27155: Delta = 69'sb111111111111111111111111111111111111111111111101111111111111111111100;
		47408: Delta = 69'sb000000000000000000000000000000000000000000000100000000000000000000100;
		3461: Delta = 69'sb111111111111111111111111111111111111111111111100000000000000000000100;
		47400: Delta = 69'sb000000000000000000000000000000000000000000000011111111111111111111100;
		3453: Delta = 69'sb111111111111111111111111111111111111111111111011111111111111111111100;
		43951: Delta = 69'sb000000000000000000000000000000000000000000001000000000000000000000100;
		6918: Delta = 69'sb111111111111111111111111111111111111111111111000000000000000000000100;
		43943: Delta = 69'sb000000000000000000000000000000000000000000000111111111111111111111100;
		6910: Delta = 69'sb111111111111111111111111111111111111111111110111111111111111111111100;
		37037: Delta = 69'sb000000000000000000000000000000000000000000010000000000000000000000100;
		13832: Delta = 69'sb111111111111111111111111111111111111111111110000000000000000000000100;
		37029: Delta = 69'sb000000000000000000000000000000000000000000001111111111111111111111100;
		13824: Delta = 69'sb111111111111111111111111111111111111111111101111111111111111111111100;
		23209: Delta = 69'sb000000000000000000000000000000000000000000100000000000000000000000100;
		27660: Delta = 69'sb111111111111111111111111111111111111111111100000000000000000000000100;
		23201: Delta = 69'sb000000000000000000000000000000000000000000011111111111111111111111100;
		27652: Delta = 69'sb111111111111111111111111111111111111111111011111111111111111111111100;
		46414: Delta = 69'sb000000000000000000000000000000000000000001000000000000000000000000100;
		4455: Delta = 69'sb111111111111111111111111111111111111111111000000000000000000000000100;
		46406: Delta = 69'sb000000000000000000000000000000000000000000111111111111111111111111100;
		4447: Delta = 69'sb111111111111111111111111111111111111111110111111111111111111111111100;
		41963: Delta = 69'sb000000000000000000000000000000000000000010000000000000000000000000100;
		8906: Delta = 69'sb111111111111111111111111111111111111111110000000000000000000000000100;
		41955: Delta = 69'sb000000000000000000000000000000000000000001111111111111111111111111100;
		8898: Delta = 69'sb111111111111111111111111111111111111111101111111111111111111111111100;
		33061: Delta = 69'sb000000000000000000000000000000000000000100000000000000000000000000100;
		17808: Delta = 69'sb111111111111111111111111111111111111111100000000000000000000000000100;
		33053: Delta = 69'sb000000000000000000000000000000000000000011111111111111111111111111100;
		17800: Delta = 69'sb111111111111111111111111111111111111111011111111111111111111111111100;
		15257: Delta = 69'sb000000000000000000000000000000000000001000000000000000000000000000100;
		35612: Delta = 69'sb111111111111111111111111111111111111111000000000000000000000000000100;
		15249: Delta = 69'sb000000000000000000000000000000000000000111111111111111111111111111100;
		35604: Delta = 69'sb111111111111111111111111111111111111110111111111111111111111111111100;
		30510: Delta = 69'sb000000000000000000000000000000000000010000000000000000000000000000100;
		20359: Delta = 69'sb111111111111111111111111111111111111110000000000000000000000000000100;
		30502: Delta = 69'sb000000000000000000000000000000000000001111111111111111111111111111100;
		20351: Delta = 69'sb111111111111111111111111111111111111101111111111111111111111111111100;
		10155: Delta = 69'sb000000000000000000000000000000000000100000000000000000000000000000100;
		40714: Delta = 69'sb111111111111111111111111111111111111100000000000000000000000000000100;
		10147: Delta = 69'sb000000000000000000000000000000000000011111111111111111111111111111100;
		40706: Delta = 69'sb111111111111111111111111111111111111011111111111111111111111111111100;
		20306: Delta = 69'sb000000000000000000000000000000000001000000000000000000000000000000100;
		30563: Delta = 69'sb111111111111111111111111111111111111000000000000000000000000000000100;
		20298: Delta = 69'sb000000000000000000000000000000000000111111111111111111111111111111100;
		30555: Delta = 69'sb111111111111111111111111111111111110111111111111111111111111111111100;
		40608: Delta = 69'sb000000000000000000000000000000000010000000000000000000000000000000100;
		10261: Delta = 69'sb111111111111111111111111111111111110000000000000000000000000000000100;
		40600: Delta = 69'sb000000000000000000000000000000000001111111111111111111111111111111100;
		10253: Delta = 69'sb111111111111111111111111111111111101111111111111111111111111111111100;
		30351: Delta = 69'sb000000000000000000000000000000000100000000000000000000000000000000100;
		20518: Delta = 69'sb111111111111111111111111111111111100000000000000000000000000000000100;
		30343: Delta = 69'sb000000000000000000000000000000000011111111111111111111111111111111100;
		20510: Delta = 69'sb111111111111111111111111111111111011111111111111111111111111111111100;
		9837: Delta = 69'sb000000000000000000000000000000001000000000000000000000000000000000100;
		41032: Delta = 69'sb111111111111111111111111111111111000000000000000000000000000000000100;
		9829: Delta = 69'sb000000000000000000000000000000000111111111111111111111111111111111100;
		41024: Delta = 69'sb111111111111111111111111111111110111111111111111111111111111111111100;
		19670: Delta = 69'sb000000000000000000000000000000010000000000000000000000000000000000100;
		31199: Delta = 69'sb111111111111111111111111111111110000000000000000000000000000000000100;
		19662: Delta = 69'sb000000000000000000000000000000001111111111111111111111111111111111100;
		31191: Delta = 69'sb111111111111111111111111111111101111111111111111111111111111111111100;
		39336: Delta = 69'sb000000000000000000000000000000100000000000000000000000000000000000100;
		11533: Delta = 69'sb111111111111111111111111111111100000000000000000000000000000000000100;
		39328: Delta = 69'sb000000000000000000000000000000011111111111111111111111111111111111100;
		11525: Delta = 69'sb111111111111111111111111111111011111111111111111111111111111111111100;
		27807: Delta = 69'sb000000000000000000000000000001000000000000000000000000000000000000100;
		23062: Delta = 69'sb111111111111111111111111111111000000000000000000000000000000000000100;
		27799: Delta = 69'sb000000000000000000000000000000111111111111111111111111111111111111100;
		23054: Delta = 69'sb111111111111111111111111111110111111111111111111111111111111111111100;
		4749: Delta = 69'sb000000000000000000000000000010000000000000000000000000000000000000100;
		46120: Delta = 69'sb111111111111111111111111111110000000000000000000000000000000000000100;
		4741: Delta = 69'sb000000000000000000000000000001111111111111111111111111111111111111100;
		46112: Delta = 69'sb111111111111111111111111111101111111111111111111111111111111111111100;
		9494: Delta = 69'sb000000000000000000000000000100000000000000000000000000000000000000100;
		41375: Delta = 69'sb111111111111111111111111111100000000000000000000000000000000000000100;
		9486: Delta = 69'sb000000000000000000000000000011111111111111111111111111111111111111100;
		41367: Delta = 69'sb111111111111111111111111111011111111111111111111111111111111111111100;
		18984: Delta = 69'sb000000000000000000000000001000000000000000000000000000000000000000100;
		31885: Delta = 69'sb111111111111111111111111111000000000000000000000000000000000000000100;
		18976: Delta = 69'sb000000000000000000000000000111111111111111111111111111111111111111100;
		31877: Delta = 69'sb111111111111111111111111110111111111111111111111111111111111111111100;
		37964: Delta = 69'sb000000000000000000000000010000000000000000000000000000000000000000100;
		12905: Delta = 69'sb111111111111111111111111110000000000000000000000000000000000000000100;
		37956: Delta = 69'sb000000000000000000000000001111111111111111111111111111111111111111100;
		12897: Delta = 69'sb111111111111111111111111101111111111111111111111111111111111111111100;
		25063: Delta = 69'sb000000000000000000000000100000000000000000000000000000000000000000100;
		25806: Delta = 69'sb111111111111111111111111100000000000000000000000000000000000000000100;
		25055: Delta = 69'sb000000000000000000000000011111111111111111111111111111111111111111100;
		25798: Delta = 69'sb111111111111111111111111011111111111111111111111111111111111111111100;
		50122: Delta = 69'sb000000000000000000000001000000000000000000000000000000000000000000100;
		747: Delta = 69'sb111111111111111111111111000000000000000000000000000000000000000000100;
		50114: Delta = 69'sb000000000000000000000000111111111111111111111111111111111111111111100;
		739: Delta = 69'sb111111111111111111111110111111111111111111111111111111111111111111100;
		49379: Delta = 69'sb000000000000000000000010000000000000000000000000000000000000000000100;
		1490: Delta = 69'sb111111111111111111111110000000000000000000000000000000000000000000100;
		49371: Delta = 69'sb000000000000000000000001111111111111111111111111111111111111111111100;
		1482: Delta = 69'sb111111111111111111111101111111111111111111111111111111111111111111100;
		47893: Delta = 69'sb000000000000000000000100000000000000000000000000000000000000000000100;
		2976: Delta = 69'sb111111111111111111111100000000000000000000000000000000000000000000100;
		47885: Delta = 69'sb000000000000000000000011111111111111111111111111111111111111111111100;
		2968: Delta = 69'sb111111111111111111111011111111111111111111111111111111111111111111100;
		44921: Delta = 69'sb000000000000000000001000000000000000000000000000000000000000000000100;
		5948: Delta = 69'sb111111111111111111111000000000000000000000000000000000000000000000100;
		44913: Delta = 69'sb000000000000000000000111111111111111111111111111111111111111111111100;
		5940: Delta = 69'sb111111111111111111110111111111111111111111111111111111111111111111100;
		38977: Delta = 69'sb000000000000000000010000000000000000000000000000000000000000000000100;
		11892: Delta = 69'sb111111111111111111110000000000000000000000000000000000000000000000100;
		38969: Delta = 69'sb000000000000000000001111111111111111111111111111111111111111111111100;
		11884: Delta = 69'sb111111111111111111101111111111111111111111111111111111111111111111100;
		27089: Delta = 69'sb000000000000000000100000000000000000000000000000000000000000000000100;
		23780: Delta = 69'sb111111111111111111100000000000000000000000000000000000000000000000100;
		27081: Delta = 69'sb000000000000000000011111111111111111111111111111111111111111111111100;
		23772: Delta = 69'sb111111111111111111011111111111111111111111111111111111111111111111100;
		3313: Delta = 69'sb000000000000000001000000000000000000000000000000000000000000000000100;
		47556: Delta = 69'sb111111111111111111000000000000000000000000000000000000000000000000100;
		3305: Delta = 69'sb000000000000000000111111111111111111111111111111111111111111111111100;
		47548: Delta = 69'sb111111111111111110111111111111111111111111111111111111111111111111100;
		6622: Delta = 69'sb000000000000000010000000000000000000000000000000000000000000000000100;
		44247: Delta = 69'sb111111111111111110000000000000000000000000000000000000000000000000100;
		6614: Delta = 69'sb000000000000000001111111111111111111111111111111111111111111111111100;
		44239: Delta = 69'sb111111111111111101111111111111111111111111111111111111111111111111100;
		13240: Delta = 69'sb000000000000000100000000000000000000000000000000000000000000000000100;
		37629: Delta = 69'sb111111111111111100000000000000000000000000000000000000000000000000100;
		13232: Delta = 69'sb000000000000000011111111111111111111111111111111111111111111111111100;
		37621: Delta = 69'sb111111111111111011111111111111111111111111111111111111111111111111100;
		26476: Delta = 69'sb000000000000001000000000000000000000000000000000000000000000000000100;
		24393: Delta = 69'sb111111111111111000000000000000000000000000000000000000000000000000100;
		26468: Delta = 69'sb000000000000000111111111111111111111111111111111111111111111111111100;
		24385: Delta = 69'sb111111111111110111111111111111111111111111111111111111111111111111100;
		2087: Delta = 69'sb000000000000010000000000000000000000000000000000000000000000000000100;
		48782: Delta = 69'sb111111111111110000000000000000000000000000000000000000000000000000100;
		2079: Delta = 69'sb000000000000001111111111111111111111111111111111111111111111111111100;
		48774: Delta = 69'sb111111111111101111111111111111111111111111111111111111111111111111100;
		4170: Delta = 69'sb000000000000100000000000000000000000000000000000000000000000000000100;
		46699: Delta = 69'sb111111111111100000000000000000000000000000000000000000000000000000100;
		4162: Delta = 69'sb000000000000011111111111111111111111111111111111111111111111111111100;
		46691: Delta = 69'sb111111111111011111111111111111111111111111111111111111111111111111100;
		8336: Delta = 69'sb000000000001000000000000000000000000000000000000000000000000000000100;
		42533: Delta = 69'sb111111111111000000000000000000000000000000000000000000000000000000100;
		8328: Delta = 69'sb000000000000111111111111111111111111111111111111111111111111111111100;
		42525: Delta = 69'sb111111111110111111111111111111111111111111111111111111111111111111100;
		16668: Delta = 69'sb000000000010000000000000000000000000000000000000000000000000000000100;
		34201: Delta = 69'sb111111111110000000000000000000000000000000000000000000000000000000100;
		16660: Delta = 69'sb000000000001111111111111111111111111111111111111111111111111111111100;
		34193: Delta = 69'sb111111111101111111111111111111111111111111111111111111111111111111100;
		33332: Delta = 69'sb000000000100000000000000000000000000000000000000000000000000000000100;
		17537: Delta = 69'sb111111111100000000000000000000000000000000000000000000000000000000100;
		33324: Delta = 69'sb000000000011111111111111111111111111111111111111111111111111111111100;
		17529: Delta = 69'sb111111111011111111111111111111111111111111111111111111111111111111100;
		15799: Delta = 69'sb000000001000000000000000000000000000000000000000000000000000000000100;
		35070: Delta = 69'sb111111111000000000000000000000000000000000000000000000000000000000100;
		15791: Delta = 69'sb000000000111111111111111111111111111111111111111111111111111111111100;
		35062: Delta = 69'sb111111110111111111111111111111111111111111111111111111111111111111100;
		31594: Delta = 69'sb000000010000000000000000000000000000000000000000000000000000000000100;
		19275: Delta = 69'sb111111110000000000000000000000000000000000000000000000000000000000100;
		31586: Delta = 69'sb000000001111111111111111111111111111111111111111111111111111111111100;
		19267: Delta = 69'sb111111101111111111111111111111111111111111111111111111111111111111100;
		12323: Delta = 69'sb000000100000000000000000000000000000000000000000000000000000000000100;
		38546: Delta = 69'sb111111100000000000000000000000000000000000000000000000000000000000100;
		12315: Delta = 69'sb000000011111111111111111111111111111111111111111111111111111111111100;
		38538: Delta = 69'sb111111011111111111111111111111111111111111111111111111111111111111100;
		24642: Delta = 69'sb000001000000000000000000000000000000000000000000000000000000000000100;
		26227: Delta = 69'sb111111000000000000000000000000000000000000000000000000000000000000100;
		24634: Delta = 69'sb000000111111111111111111111111111111111111111111111111111111111111100;
		26219: Delta = 69'sb111110111111111111111111111111111111111111111111111111111111111111100;
		49280: Delta = 69'sb000010000000000000000000000000000000000000000000000000000000000000100;
		1589: Delta = 69'sb111110000000000000000000000000000000000000000000000000000000000000100;
		49272: Delta = 69'sb000001111111111111111111111111111111111111111111111111111111111111100;
		1581: Delta = 69'sb111101111111111111111111111111111111111111111111111111111111111111100;
		47695: Delta = 69'sb000100000000000000000000000000000000000000000000000000000000000000100;
		3174: Delta = 69'sb111100000000000000000000000000000000000000000000000000000000000000100;
		47687: Delta = 69'sb000011111111111111111111111111111111111111111111111111111111111111100;
		3166: Delta = 69'sb111011111111111111111111111111111111111111111111111111111111111111100;
		44525: Delta = 69'sb001000000000000000000000000000000000000000000000000000000000000000100;
		6344: Delta = 69'sb111000000000000000000000000000000000000000000000000000000000000000100;
		44517: Delta = 69'sb000111111111111111111111111111111111111111111111111111111111111111100;
		6336: Delta = 69'sb110111111111111111111111111111111111111111111111111111111111111111100;
		38185: Delta = 69'sb010000000000000000000000000000000000000000000000000000000000000000100;
		12684: Delta = 69'sb110000000000000000000000000000000000000000000000000000000000000000100;
		38177: Delta = 69'sb001111111111111111111111111111111111111111111111111111111111111111100;
		12676: Delta = 69'sb101111111111111111111111111111111111111111111111111111111111111111100;
		24: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000011000;
		50837: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111101000;
		40: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000101000;
		50821: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111011000;
		72: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000001001000;
		50805: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111001000;
		56: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000111000;
		50789: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111110111000;
		136: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000010001000;
		50741: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111110001000;
		120: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000001111000;
		50725: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111101111000;
		264: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000100001000;
		50613: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111100001000;
		248: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000011111000;
		50597: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111011111000;
		520: Delta = 69'sb000000000000000000000000000000000000000000000000000000000001000001000;
		50357: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111000001000;
		504: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000111111000;
		50341: Delta = 69'sb111111111111111111111111111111111111111111111111111111111110111111000;
		1032: Delta = 69'sb000000000000000000000000000000000000000000000000000000000010000001000;
		49845: Delta = 69'sb111111111111111111111111111111111111111111111111111111111110000001000;
		1016: Delta = 69'sb000000000000000000000000000000000000000000000000000000000001111111000;
		49829: Delta = 69'sb111111111111111111111111111111111111111111111111111111111101111111000;
		2056: Delta = 69'sb000000000000000000000000000000000000000000000000000000000100000001000;
		48821: Delta = 69'sb111111111111111111111111111111111111111111111111111111111100000001000;
		2040: Delta = 69'sb000000000000000000000000000000000000000000000000000000000011111111000;
		48805: Delta = 69'sb111111111111111111111111111111111111111111111111111111111011111111000;
		4104: Delta = 69'sb000000000000000000000000000000000000000000000000000000001000000001000;
		46773: Delta = 69'sb111111111111111111111111111111111111111111111111111111111000000001000;
		4088: Delta = 69'sb000000000000000000000000000000000000000000000000000000000111111111000;
		46757: Delta = 69'sb111111111111111111111111111111111111111111111111111111110111111111000;
		8200: Delta = 69'sb000000000000000000000000000000000000000000000000000000010000000001000;
		42677: Delta = 69'sb111111111111111111111111111111111111111111111111111111110000000001000;
		8184: Delta = 69'sb000000000000000000000000000000000000000000000000000000001111111111000;
		42661: Delta = 69'sb111111111111111111111111111111111111111111111111111111101111111111000;
		16392: Delta = 69'sb000000000000000000000000000000000000000000000000000000100000000001000;
		34485: Delta = 69'sb111111111111111111111111111111111111111111111111111111100000000001000;
		16376: Delta = 69'sb000000000000000000000000000000000000000000000000000000011111111111000;
		34469: Delta = 69'sb111111111111111111111111111111111111111111111111111111011111111111000;
		32776: Delta = 69'sb000000000000000000000000000000000000000000000000000001000000000001000;
		18101: Delta = 69'sb111111111111111111111111111111111111111111111111111111000000000001000;
		32760: Delta = 69'sb000000000000000000000000000000000000000000000000000000111111111111000;
		18085: Delta = 69'sb111111111111111111111111111111111111111111111111111110111111111111000;
		14683: Delta = 69'sb000000000000000000000000000000000000000000000000000010000000000001000;
		36194: Delta = 69'sb111111111111111111111111111111111111111111111111111110000000000001000;
		14667: Delta = 69'sb000000000000000000000000000000000000000000000000000001111111111111000;
		36178: Delta = 69'sb111111111111111111111111111111111111111111111111111101111111111111000;
		29358: Delta = 69'sb000000000000000000000000000000000000000000000000000100000000000001000;
		21519: Delta = 69'sb111111111111111111111111111111111111111111111111111100000000000001000;
		29342: Delta = 69'sb000000000000000000000000000000000000000000000000000011111111111111000;
		21503: Delta = 69'sb111111111111111111111111111111111111111111111111111011111111111111000;
		7847: Delta = 69'sb000000000000000000000000000000000000000000000000001000000000000001000;
		43030: Delta = 69'sb111111111111111111111111111111111111111111111111111000000000000001000;
		7831: Delta = 69'sb000000000000000000000000000000000000000000000000000111111111111111000;
		43014: Delta = 69'sb111111111111111111111111111111111111111111111111110111111111111111000;
		15686: Delta = 69'sb000000000000000000000000000000000000000000000000010000000000000001000;
		35191: Delta = 69'sb111111111111111111111111111111111111111111111111110000000000000001000;
		15670: Delta = 69'sb000000000000000000000000000000000000000000000000001111111111111111000;
		35175: Delta = 69'sb111111111111111111111111111111111111111111111111101111111111111111000;
		31364: Delta = 69'sb000000000000000000000000000000000000000000000000100000000000000001000;
		19513: Delta = 69'sb111111111111111111111111111111111111111111111111100000000000000001000;
		31348: Delta = 69'sb000000000000000000000000000000000000000000000000011111111111111111000;
		19497: Delta = 69'sb111111111111111111111111111111111111111111111111011111111111111111000;
		11859: Delta = 69'sb000000000000000000000000000000000000000000000001000000000000000001000;
		39018: Delta = 69'sb111111111111111111111111111111111111111111111111000000000000000001000;
		11843: Delta = 69'sb000000000000000000000000000000000000000000000000111111111111111111000;
		39002: Delta = 69'sb111111111111111111111111111111111111111111111110111111111111111111000;
		23710: Delta = 69'sb000000000000000000000000000000000000000000000010000000000000000001000;
		27167: Delta = 69'sb111111111111111111111111111111111111111111111110000000000000000001000;
		23694: Delta = 69'sb000000000000000000000000000000000000000000000001111111111111111111000;
		27151: Delta = 69'sb111111111111111111111111111111111111111111111101111111111111111111000;
		47412: Delta = 69'sb000000000000000000000000000000000000000000000100000000000000000001000;
		3465: Delta = 69'sb111111111111111111111111111111111111111111111100000000000000000001000;
		47396: Delta = 69'sb000000000000000000000000000000000000000000000011111111111111111111000;
		3449: Delta = 69'sb111111111111111111111111111111111111111111111011111111111111111111000;
		43955: Delta = 69'sb000000000000000000000000000000000000000000001000000000000000000001000;
		6922: Delta = 69'sb111111111111111111111111111111111111111111111000000000000000000001000;
		43939: Delta = 69'sb000000000000000000000000000000000000000000000111111111111111111111000;
		6906: Delta = 69'sb111111111111111111111111111111111111111111110111111111111111111111000;
		37041: Delta = 69'sb000000000000000000000000000000000000000000010000000000000000000001000;
		13836: Delta = 69'sb111111111111111111111111111111111111111111110000000000000000000001000;
		37025: Delta = 69'sb000000000000000000000000000000000000000000001111111111111111111111000;
		13820: Delta = 69'sb111111111111111111111111111111111111111111101111111111111111111111000;
		23213: Delta = 69'sb000000000000000000000000000000000000000000100000000000000000000001000;
		27664: Delta = 69'sb111111111111111111111111111111111111111111100000000000000000000001000;
		23197: Delta = 69'sb000000000000000000000000000000000000000000011111111111111111111111000;
		27648: Delta = 69'sb111111111111111111111111111111111111111111011111111111111111111111000;
		46418: Delta = 69'sb000000000000000000000000000000000000000001000000000000000000000001000;
		4459: Delta = 69'sb111111111111111111111111111111111111111111000000000000000000000001000;
		46402: Delta = 69'sb000000000000000000000000000000000000000000111111111111111111111111000;
		4443: Delta = 69'sb111111111111111111111111111111111111111110111111111111111111111111000;
		41967: Delta = 69'sb000000000000000000000000000000000000000010000000000000000000000001000;
		8910: Delta = 69'sb111111111111111111111111111111111111111110000000000000000000000001000;
		41951: Delta = 69'sb000000000000000000000000000000000000000001111111111111111111111111000;
		8894: Delta = 69'sb111111111111111111111111111111111111111101111111111111111111111111000;
		33065: Delta = 69'sb000000000000000000000000000000000000000100000000000000000000000001000;
		17812: Delta = 69'sb111111111111111111111111111111111111111100000000000000000000000001000;
		33049: Delta = 69'sb000000000000000000000000000000000000000011111111111111111111111111000;
		17796: Delta = 69'sb111111111111111111111111111111111111111011111111111111111111111111000;
		15261: Delta = 69'sb000000000000000000000000000000000000001000000000000000000000000001000;
		35616: Delta = 69'sb111111111111111111111111111111111111111000000000000000000000000001000;
		15245: Delta = 69'sb000000000000000000000000000000000000000111111111111111111111111111000;
		35600: Delta = 69'sb111111111111111111111111111111111111110111111111111111111111111111000;
		30514: Delta = 69'sb000000000000000000000000000000000000010000000000000000000000000001000;
		20363: Delta = 69'sb111111111111111111111111111111111111110000000000000000000000000001000;
		30498: Delta = 69'sb000000000000000000000000000000000000001111111111111111111111111111000;
		20347: Delta = 69'sb111111111111111111111111111111111111101111111111111111111111111111000;
		10159: Delta = 69'sb000000000000000000000000000000000000100000000000000000000000000001000;
		40718: Delta = 69'sb111111111111111111111111111111111111100000000000000000000000000001000;
		10143: Delta = 69'sb000000000000000000000000000000000000011111111111111111111111111111000;
		40702: Delta = 69'sb111111111111111111111111111111111111011111111111111111111111111111000;
		20310: Delta = 69'sb000000000000000000000000000000000001000000000000000000000000000001000;
		30567: Delta = 69'sb111111111111111111111111111111111111000000000000000000000000000001000;
		20294: Delta = 69'sb000000000000000000000000000000000000111111111111111111111111111111000;
		30551: Delta = 69'sb111111111111111111111111111111111110111111111111111111111111111111000;
		40612: Delta = 69'sb000000000000000000000000000000000010000000000000000000000000000001000;
		10265: Delta = 69'sb111111111111111111111111111111111110000000000000000000000000000001000;
		40596: Delta = 69'sb000000000000000000000000000000000001111111111111111111111111111111000;
		10249: Delta = 69'sb111111111111111111111111111111111101111111111111111111111111111111000;
		30355: Delta = 69'sb000000000000000000000000000000000100000000000000000000000000000001000;
		20522: Delta = 69'sb111111111111111111111111111111111100000000000000000000000000000001000;
		30339: Delta = 69'sb000000000000000000000000000000000011111111111111111111111111111111000;
		20506: Delta = 69'sb111111111111111111111111111111111011111111111111111111111111111111000;
		9841: Delta = 69'sb000000000000000000000000000000001000000000000000000000000000000001000;
		41036: Delta = 69'sb111111111111111111111111111111111000000000000000000000000000000001000;
		9825: Delta = 69'sb000000000000000000000000000000000111111111111111111111111111111111000;
		41020: Delta = 69'sb111111111111111111111111111111110111111111111111111111111111111111000;
		19674: Delta = 69'sb000000000000000000000000000000010000000000000000000000000000000001000;
		31203: Delta = 69'sb111111111111111111111111111111110000000000000000000000000000000001000;
		19658: Delta = 69'sb000000000000000000000000000000001111111111111111111111111111111111000;
		31187: Delta = 69'sb111111111111111111111111111111101111111111111111111111111111111111000;
		39340: Delta = 69'sb000000000000000000000000000000100000000000000000000000000000000001000;
		11537: Delta = 69'sb111111111111111111111111111111100000000000000000000000000000000001000;
		39324: Delta = 69'sb000000000000000000000000000000011111111111111111111111111111111111000;
		11521: Delta = 69'sb111111111111111111111111111111011111111111111111111111111111111111000;
		27811: Delta = 69'sb000000000000000000000000000001000000000000000000000000000000000001000;
		23066: Delta = 69'sb111111111111111111111111111111000000000000000000000000000000000001000;
		27795: Delta = 69'sb000000000000000000000000000000111111111111111111111111111111111111000;
		23050: Delta = 69'sb111111111111111111111111111110111111111111111111111111111111111111000;
		4753: Delta = 69'sb000000000000000000000000000010000000000000000000000000000000000001000;
		46124: Delta = 69'sb111111111111111111111111111110000000000000000000000000000000000001000;
		4737: Delta = 69'sb000000000000000000000000000001111111111111111111111111111111111111000;
		46108: Delta = 69'sb111111111111111111111111111101111111111111111111111111111111111111000;
		9498: Delta = 69'sb000000000000000000000000000100000000000000000000000000000000000001000;
		41379: Delta = 69'sb111111111111111111111111111100000000000000000000000000000000000001000;
		9482: Delta = 69'sb000000000000000000000000000011111111111111111111111111111111111111000;
		41363: Delta = 69'sb111111111111111111111111111011111111111111111111111111111111111111000;
		18988: Delta = 69'sb000000000000000000000000001000000000000000000000000000000000000001000;
		31889: Delta = 69'sb111111111111111111111111111000000000000000000000000000000000000001000;
		18972: Delta = 69'sb000000000000000000000000000111111111111111111111111111111111111111000;
		31873: Delta = 69'sb111111111111111111111111110111111111111111111111111111111111111111000;
		37968: Delta = 69'sb000000000000000000000000010000000000000000000000000000000000000001000;
		12909: Delta = 69'sb111111111111111111111111110000000000000000000000000000000000000001000;
		37952: Delta = 69'sb000000000000000000000000001111111111111111111111111111111111111111000;
		12893: Delta = 69'sb111111111111111111111111101111111111111111111111111111111111111111000;
		25067: Delta = 69'sb000000000000000000000000100000000000000000000000000000000000000001000;
		25810: Delta = 69'sb111111111111111111111111100000000000000000000000000000000000000001000;
		25051: Delta = 69'sb000000000000000000000000011111111111111111111111111111111111111111000;
		25794: Delta = 69'sb111111111111111111111111011111111111111111111111111111111111111111000;
		50126: Delta = 69'sb000000000000000000000001000000000000000000000000000000000000000001000;
		751: Delta = 69'sb111111111111111111111111000000000000000000000000000000000000000001000;
		50110: Delta = 69'sb000000000000000000000000111111111111111111111111111111111111111111000;
		735: Delta = 69'sb111111111111111111111110111111111111111111111111111111111111111111000;
		49383: Delta = 69'sb000000000000000000000010000000000000000000000000000000000000000001000;
		1494: Delta = 69'sb111111111111111111111110000000000000000000000000000000000000000001000;
		49367: Delta = 69'sb000000000000000000000001111111111111111111111111111111111111111111000;
		1478: Delta = 69'sb111111111111111111111101111111111111111111111111111111111111111111000;
		47897: Delta = 69'sb000000000000000000000100000000000000000000000000000000000000000001000;
		2980: Delta = 69'sb111111111111111111111100000000000000000000000000000000000000000001000;
		47881: Delta = 69'sb000000000000000000000011111111111111111111111111111111111111111111000;
		2964: Delta = 69'sb111111111111111111111011111111111111111111111111111111111111111111000;
		44925: Delta = 69'sb000000000000000000001000000000000000000000000000000000000000000001000;
		5952: Delta = 69'sb111111111111111111111000000000000000000000000000000000000000000001000;
		44909: Delta = 69'sb000000000000000000000111111111111111111111111111111111111111111111000;
		5936: Delta = 69'sb111111111111111111110111111111111111111111111111111111111111111111000;
		38981: Delta = 69'sb000000000000000000010000000000000000000000000000000000000000000001000;
		11896: Delta = 69'sb111111111111111111110000000000000000000000000000000000000000000001000;
		38965: Delta = 69'sb000000000000000000001111111111111111111111111111111111111111111111000;
		11880: Delta = 69'sb111111111111111111101111111111111111111111111111111111111111111111000;
		27093: Delta = 69'sb000000000000000000100000000000000000000000000000000000000000000001000;
		23784: Delta = 69'sb111111111111111111100000000000000000000000000000000000000000000001000;
		27077: Delta = 69'sb000000000000000000011111111111111111111111111111111111111111111111000;
		23768: Delta = 69'sb111111111111111111011111111111111111111111111111111111111111111111000;
		3317: Delta = 69'sb000000000000000001000000000000000000000000000000000000000000000001000;
		47560: Delta = 69'sb111111111111111111000000000000000000000000000000000000000000000001000;
		3301: Delta = 69'sb000000000000000000111111111111111111111111111111111111111111111111000;
		47544: Delta = 69'sb111111111111111110111111111111111111111111111111111111111111111111000;
		6626: Delta = 69'sb000000000000000010000000000000000000000000000000000000000000000001000;
		44251: Delta = 69'sb111111111111111110000000000000000000000000000000000000000000000001000;
		6610: Delta = 69'sb000000000000000001111111111111111111111111111111111111111111111111000;
		44235: Delta = 69'sb111111111111111101111111111111111111111111111111111111111111111111000;
		13244: Delta = 69'sb000000000000000100000000000000000000000000000000000000000000000001000;
		37633: Delta = 69'sb111111111111111100000000000000000000000000000000000000000000000001000;
		13228: Delta = 69'sb000000000000000011111111111111111111111111111111111111111111111111000;
		37617: Delta = 69'sb111111111111111011111111111111111111111111111111111111111111111111000;
		26480: Delta = 69'sb000000000000001000000000000000000000000000000000000000000000000001000;
		24397: Delta = 69'sb111111111111111000000000000000000000000000000000000000000000000001000;
		26464: Delta = 69'sb000000000000000111111111111111111111111111111111111111111111111111000;
		24381: Delta = 69'sb111111111111110111111111111111111111111111111111111111111111111111000;
		2091: Delta = 69'sb000000000000010000000000000000000000000000000000000000000000000001000;
		48786: Delta = 69'sb111111111111110000000000000000000000000000000000000000000000000001000;
		2075: Delta = 69'sb000000000000001111111111111111111111111111111111111111111111111111000;
		48770: Delta = 69'sb111111111111101111111111111111111111111111111111111111111111111111000;
		4174: Delta = 69'sb000000000000100000000000000000000000000000000000000000000000000001000;
		46703: Delta = 69'sb111111111111100000000000000000000000000000000000000000000000000001000;
		4158: Delta = 69'sb000000000000011111111111111111111111111111111111111111111111111111000;
		46687: Delta = 69'sb111111111111011111111111111111111111111111111111111111111111111111000;
		8340: Delta = 69'sb000000000001000000000000000000000000000000000000000000000000000001000;
		42537: Delta = 69'sb111111111111000000000000000000000000000000000000000000000000000001000;
		8324: Delta = 69'sb000000000000111111111111111111111111111111111111111111111111111111000;
		42521: Delta = 69'sb111111111110111111111111111111111111111111111111111111111111111111000;
		16672: Delta = 69'sb000000000010000000000000000000000000000000000000000000000000000001000;
		34205: Delta = 69'sb111111111110000000000000000000000000000000000000000000000000000001000;
		16656: Delta = 69'sb000000000001111111111111111111111111111111111111111111111111111111000;
		34189: Delta = 69'sb111111111101111111111111111111111111111111111111111111111111111111000;
		33336: Delta = 69'sb000000000100000000000000000000000000000000000000000000000000000001000;
		17541: Delta = 69'sb111111111100000000000000000000000000000000000000000000000000000001000;
		33320: Delta = 69'sb000000000011111111111111111111111111111111111111111111111111111111000;
		17525: Delta = 69'sb111111111011111111111111111111111111111111111111111111111111111111000;
		15803: Delta = 69'sb000000001000000000000000000000000000000000000000000000000000000001000;
		35074: Delta = 69'sb111111111000000000000000000000000000000000000000000000000000000001000;
		15787: Delta = 69'sb000000000111111111111111111111111111111111111111111111111111111111000;
		35058: Delta = 69'sb111111110111111111111111111111111111111111111111111111111111111111000;
		31598: Delta = 69'sb000000010000000000000000000000000000000000000000000000000000000001000;
		19279: Delta = 69'sb111111110000000000000000000000000000000000000000000000000000000001000;
		31582: Delta = 69'sb000000001111111111111111111111111111111111111111111111111111111111000;
		19263: Delta = 69'sb111111101111111111111111111111111111111111111111111111111111111111000;
		12327: Delta = 69'sb000000100000000000000000000000000000000000000000000000000000000001000;
		38550: Delta = 69'sb111111100000000000000000000000000000000000000000000000000000000001000;
		12311: Delta = 69'sb000000011111111111111111111111111111111111111111111111111111111111000;
		38534: Delta = 69'sb111111011111111111111111111111111111111111111111111111111111111111000;
		24646: Delta = 69'sb000001000000000000000000000000000000000000000000000000000000000001000;
		26231: Delta = 69'sb111111000000000000000000000000000000000000000000000000000000000001000;
		24630: Delta = 69'sb000000111111111111111111111111111111111111111111111111111111111111000;
		26215: Delta = 69'sb111110111111111111111111111111111111111111111111111111111111111111000;
		49284: Delta = 69'sb000010000000000000000000000000000000000000000000000000000000000001000;
		1593: Delta = 69'sb111110000000000000000000000000000000000000000000000000000000000001000;
		49268: Delta = 69'sb000001111111111111111111111111111111111111111111111111111111111111000;
		1577: Delta = 69'sb111101111111111111111111111111111111111111111111111111111111111111000;
		47699: Delta = 69'sb000100000000000000000000000000000000000000000000000000000000000001000;
		3178: Delta = 69'sb111100000000000000000000000000000000000000000000000000000000000001000;
		47683: Delta = 69'sb000011111111111111111111111111111111111111111111111111111111111111000;
		3162: Delta = 69'sb111011111111111111111111111111111111111111111111111111111111111111000;
		44529: Delta = 69'sb001000000000000000000000000000000000000000000000000000000000000001000;
		6348: Delta = 69'sb111000000000000000000000000000000000000000000000000000000000000001000;
		44513: Delta = 69'sb000111111111111111111111111111111111111111111111111111111111111111000;
		6332: Delta = 69'sb110111111111111111111111111111111111111111111111111111111111111111000;
		38189: Delta = 69'sb010000000000000000000000000000000000000000000000000000000000000001000;
		12688: Delta = 69'sb110000000000000000000000000000000000000000000000000000000000000001000;
		38173: Delta = 69'sb001111111111111111111111111111111111111111111111111111111111111111000;
		12672: Delta = 69'sb101111111111111111111111111111111111111111111111111111111111111111000;
		48: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000000110000;
		50813: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111111010000;
		80: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000001010000;
		50781: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111110110000;
		144: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000010010000;
		50749: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111110010000;
		112: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000001110000;
		50717: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111101110000;
		272: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000100010000;
		50621: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111100010000;
		240: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000011110000;
		50589: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111011110000;
		528: Delta = 69'sb000000000000000000000000000000000000000000000000000000000001000010000;
		50365: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111000010000;
		496: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000111110000;
		50333: Delta = 69'sb111111111111111111111111111111111111111111111111111111111110111110000;
		1040: Delta = 69'sb000000000000000000000000000000000000000000000000000000000010000010000;
		49853: Delta = 69'sb111111111111111111111111111111111111111111111111111111111110000010000;
		1008: Delta = 69'sb000000000000000000000000000000000000000000000000000000000001111110000;
		49821: Delta = 69'sb111111111111111111111111111111111111111111111111111111111101111110000;
		2064: Delta = 69'sb000000000000000000000000000000000000000000000000000000000100000010000;
		48829: Delta = 69'sb111111111111111111111111111111111111111111111111111111111100000010000;
		2032: Delta = 69'sb000000000000000000000000000000000000000000000000000000000011111110000;
		48797: Delta = 69'sb111111111111111111111111111111111111111111111111111111111011111110000;
		4112: Delta = 69'sb000000000000000000000000000000000000000000000000000000001000000010000;
		46781: Delta = 69'sb111111111111111111111111111111111111111111111111111111111000000010000;
		4080: Delta = 69'sb000000000000000000000000000000000000000000000000000000000111111110000;
		46749: Delta = 69'sb111111111111111111111111111111111111111111111111111111110111111110000;
		8208: Delta = 69'sb000000000000000000000000000000000000000000000000000000010000000010000;
		42685: Delta = 69'sb111111111111111111111111111111111111111111111111111111110000000010000;
		8176: Delta = 69'sb000000000000000000000000000000000000000000000000000000001111111110000;
		42653: Delta = 69'sb111111111111111111111111111111111111111111111111111111101111111110000;
		16400: Delta = 69'sb000000000000000000000000000000000000000000000000000000100000000010000;
		34493: Delta = 69'sb111111111111111111111111111111111111111111111111111111100000000010000;
		16368: Delta = 69'sb000000000000000000000000000000000000000000000000000000011111111110000;
		34461: Delta = 69'sb111111111111111111111111111111111111111111111111111111011111111110000;
		32784: Delta = 69'sb000000000000000000000000000000000000000000000000000001000000000010000;
		18109: Delta = 69'sb111111111111111111111111111111111111111111111111111111000000000010000;
		32752: Delta = 69'sb000000000000000000000000000000000000000000000000000000111111111110000;
		18077: Delta = 69'sb111111111111111111111111111111111111111111111111111110111111111110000;
		14691: Delta = 69'sb000000000000000000000000000000000000000000000000000010000000000010000;
		36202: Delta = 69'sb111111111111111111111111111111111111111111111111111110000000000010000;
		14659: Delta = 69'sb000000000000000000000000000000000000000000000000000001111111111110000;
		36170: Delta = 69'sb111111111111111111111111111111111111111111111111111101111111111110000;
		29366: Delta = 69'sb000000000000000000000000000000000000000000000000000100000000000010000;
		21527: Delta = 69'sb111111111111111111111111111111111111111111111111111100000000000010000;
		29334: Delta = 69'sb000000000000000000000000000000000000000000000000000011111111111110000;
		21495: Delta = 69'sb111111111111111111111111111111111111111111111111111011111111111110000;
		7855: Delta = 69'sb000000000000000000000000000000000000000000000000001000000000000010000;
		43038: Delta = 69'sb111111111111111111111111111111111111111111111111111000000000000010000;
		7823: Delta = 69'sb000000000000000000000000000000000000000000000000000111111111111110000;
		43006: Delta = 69'sb111111111111111111111111111111111111111111111111110111111111111110000;
		15694: Delta = 69'sb000000000000000000000000000000000000000000000000010000000000000010000;
		35199: Delta = 69'sb111111111111111111111111111111111111111111111111110000000000000010000;
		15662: Delta = 69'sb000000000000000000000000000000000000000000000000001111111111111110000;
		35167: Delta = 69'sb111111111111111111111111111111111111111111111111101111111111111110000;
		31372: Delta = 69'sb000000000000000000000000000000000000000000000000100000000000000010000;
		19521: Delta = 69'sb111111111111111111111111111111111111111111111111100000000000000010000;
		31340: Delta = 69'sb000000000000000000000000000000000000000000000000011111111111111110000;
		19489: Delta = 69'sb111111111111111111111111111111111111111111111111011111111111111110000;
		11867: Delta = 69'sb000000000000000000000000000000000000000000000001000000000000000010000;
		39026: Delta = 69'sb111111111111111111111111111111111111111111111111000000000000000010000;
		11835: Delta = 69'sb000000000000000000000000000000000000000000000000111111111111111110000;
		38994: Delta = 69'sb111111111111111111111111111111111111111111111110111111111111111110000;
		23718: Delta = 69'sb000000000000000000000000000000000000000000000010000000000000000010000;
		27175: Delta = 69'sb111111111111111111111111111111111111111111111110000000000000000010000;
		23686: Delta = 69'sb000000000000000000000000000000000000000000000001111111111111111110000;
		27143: Delta = 69'sb111111111111111111111111111111111111111111111101111111111111111110000;
		47420: Delta = 69'sb000000000000000000000000000000000000000000000100000000000000000010000;
		3473: Delta = 69'sb111111111111111111111111111111111111111111111100000000000000000010000;
		47388: Delta = 69'sb000000000000000000000000000000000000000000000011111111111111111110000;
		3441: Delta = 69'sb111111111111111111111111111111111111111111111011111111111111111110000;
		43963: Delta = 69'sb000000000000000000000000000000000000000000001000000000000000000010000;
		6930: Delta = 69'sb111111111111111111111111111111111111111111111000000000000000000010000;
		43931: Delta = 69'sb000000000000000000000000000000000000000000000111111111111111111110000;
		6898: Delta = 69'sb111111111111111111111111111111111111111111110111111111111111111110000;
		37049: Delta = 69'sb000000000000000000000000000000000000000000010000000000000000000010000;
		13844: Delta = 69'sb111111111111111111111111111111111111111111110000000000000000000010000;
		37017: Delta = 69'sb000000000000000000000000000000000000000000001111111111111111111110000;
		13812: Delta = 69'sb111111111111111111111111111111111111111111101111111111111111111110000;
		23221: Delta = 69'sb000000000000000000000000000000000000000000100000000000000000000010000;
		27672: Delta = 69'sb111111111111111111111111111111111111111111100000000000000000000010000;
		23189: Delta = 69'sb000000000000000000000000000000000000000000011111111111111111111110000;
		27640: Delta = 69'sb111111111111111111111111111111111111111111011111111111111111111110000;
		46426: Delta = 69'sb000000000000000000000000000000000000000001000000000000000000000010000;
		4467: Delta = 69'sb111111111111111111111111111111111111111111000000000000000000000010000;
		46394: Delta = 69'sb000000000000000000000000000000000000000000111111111111111111111110000;
		4435: Delta = 69'sb111111111111111111111111111111111111111110111111111111111111111110000;
		41975: Delta = 69'sb000000000000000000000000000000000000000010000000000000000000000010000;
		8918: Delta = 69'sb111111111111111111111111111111111111111110000000000000000000000010000;
		41943: Delta = 69'sb000000000000000000000000000000000000000001111111111111111111111110000;
		8886: Delta = 69'sb111111111111111111111111111111111111111101111111111111111111111110000;
		33073: Delta = 69'sb000000000000000000000000000000000000000100000000000000000000000010000;
		17820: Delta = 69'sb111111111111111111111111111111111111111100000000000000000000000010000;
		33041: Delta = 69'sb000000000000000000000000000000000000000011111111111111111111111110000;
		17788: Delta = 69'sb111111111111111111111111111111111111111011111111111111111111111110000;
		15269: Delta = 69'sb000000000000000000000000000000000000001000000000000000000000000010000;
		35624: Delta = 69'sb111111111111111111111111111111111111111000000000000000000000000010000;
		15237: Delta = 69'sb000000000000000000000000000000000000000111111111111111111111111110000;
		35592: Delta = 69'sb111111111111111111111111111111111111110111111111111111111111111110000;
		30522: Delta = 69'sb000000000000000000000000000000000000010000000000000000000000000010000;
		20371: Delta = 69'sb111111111111111111111111111111111111110000000000000000000000000010000;
		30490: Delta = 69'sb000000000000000000000000000000000000001111111111111111111111111110000;
		20339: Delta = 69'sb111111111111111111111111111111111111101111111111111111111111111110000;
		10167: Delta = 69'sb000000000000000000000000000000000000100000000000000000000000000010000;
		40726: Delta = 69'sb111111111111111111111111111111111111100000000000000000000000000010000;
		10135: Delta = 69'sb000000000000000000000000000000000000011111111111111111111111111110000;
		40694: Delta = 69'sb111111111111111111111111111111111111011111111111111111111111111110000;
		20318: Delta = 69'sb000000000000000000000000000000000001000000000000000000000000000010000;
		30575: Delta = 69'sb111111111111111111111111111111111111000000000000000000000000000010000;
		20286: Delta = 69'sb000000000000000000000000000000000000111111111111111111111111111110000;
		30543: Delta = 69'sb111111111111111111111111111111111110111111111111111111111111111110000;
		40620: Delta = 69'sb000000000000000000000000000000000010000000000000000000000000000010000;
		10273: Delta = 69'sb111111111111111111111111111111111110000000000000000000000000000010000;
		40588: Delta = 69'sb000000000000000000000000000000000001111111111111111111111111111110000;
		10241: Delta = 69'sb111111111111111111111111111111111101111111111111111111111111111110000;
		30363: Delta = 69'sb000000000000000000000000000000000100000000000000000000000000000010000;
		20530: Delta = 69'sb111111111111111111111111111111111100000000000000000000000000000010000;
		30331: Delta = 69'sb000000000000000000000000000000000011111111111111111111111111111110000;
		20498: Delta = 69'sb111111111111111111111111111111111011111111111111111111111111111110000;
		9849: Delta = 69'sb000000000000000000000000000000001000000000000000000000000000000010000;
		41044: Delta = 69'sb111111111111111111111111111111111000000000000000000000000000000010000;
		9817: Delta = 69'sb000000000000000000000000000000000111111111111111111111111111111110000;
		41012: Delta = 69'sb111111111111111111111111111111110111111111111111111111111111111110000;
		19682: Delta = 69'sb000000000000000000000000000000010000000000000000000000000000000010000;
		31211: Delta = 69'sb111111111111111111111111111111110000000000000000000000000000000010000;
		19650: Delta = 69'sb000000000000000000000000000000001111111111111111111111111111111110000;
		31179: Delta = 69'sb111111111111111111111111111111101111111111111111111111111111111110000;
		39348: Delta = 69'sb000000000000000000000000000000100000000000000000000000000000000010000;
		11545: Delta = 69'sb111111111111111111111111111111100000000000000000000000000000000010000;
		39316: Delta = 69'sb000000000000000000000000000000011111111111111111111111111111111110000;
		11513: Delta = 69'sb111111111111111111111111111111011111111111111111111111111111111110000;
		27819: Delta = 69'sb000000000000000000000000000001000000000000000000000000000000000010000;
		23074: Delta = 69'sb111111111111111111111111111111000000000000000000000000000000000010000;
		27787: Delta = 69'sb000000000000000000000000000000111111111111111111111111111111111110000;
		23042: Delta = 69'sb111111111111111111111111111110111111111111111111111111111111111110000;
		4761: Delta = 69'sb000000000000000000000000000010000000000000000000000000000000000010000;
		46132: Delta = 69'sb111111111111111111111111111110000000000000000000000000000000000010000;
		4729: Delta = 69'sb000000000000000000000000000001111111111111111111111111111111111110000;
		46100: Delta = 69'sb111111111111111111111111111101111111111111111111111111111111111110000;
		9506: Delta = 69'sb000000000000000000000000000100000000000000000000000000000000000010000;
		41387: Delta = 69'sb111111111111111111111111111100000000000000000000000000000000000010000;
		9474: Delta = 69'sb000000000000000000000000000011111111111111111111111111111111111110000;
		41355: Delta = 69'sb111111111111111111111111111011111111111111111111111111111111111110000;
		18996: Delta = 69'sb000000000000000000000000001000000000000000000000000000000000000010000;
		31897: Delta = 69'sb111111111111111111111111111000000000000000000000000000000000000010000;
		18964: Delta = 69'sb000000000000000000000000000111111111111111111111111111111111111110000;
		31865: Delta = 69'sb111111111111111111111111110111111111111111111111111111111111111110000;
		37976: Delta = 69'sb000000000000000000000000010000000000000000000000000000000000000010000;
		12917: Delta = 69'sb111111111111111111111111110000000000000000000000000000000000000010000;
		37944: Delta = 69'sb000000000000000000000000001111111111111111111111111111111111111110000;
		12885: Delta = 69'sb111111111111111111111111101111111111111111111111111111111111111110000;
		25075: Delta = 69'sb000000000000000000000000100000000000000000000000000000000000000010000;
		25818: Delta = 69'sb111111111111111111111111100000000000000000000000000000000000000010000;
		25043: Delta = 69'sb000000000000000000000000011111111111111111111111111111111111111110000;
		25786: Delta = 69'sb111111111111111111111111011111111111111111111111111111111111111110000;
		50134: Delta = 69'sb000000000000000000000001000000000000000000000000000000000000000010000;
		759: Delta = 69'sb111111111111111111111111000000000000000000000000000000000000000010000;
		50102: Delta = 69'sb000000000000000000000000111111111111111111111111111111111111111110000;
		727: Delta = 69'sb111111111111111111111110111111111111111111111111111111111111111110000;
		49391: Delta = 69'sb000000000000000000000010000000000000000000000000000000000000000010000;
		1502: Delta = 69'sb111111111111111111111110000000000000000000000000000000000000000010000;
		49359: Delta = 69'sb000000000000000000000001111111111111111111111111111111111111111110000;
		1470: Delta = 69'sb111111111111111111111101111111111111111111111111111111111111111110000;
		47905: Delta = 69'sb000000000000000000000100000000000000000000000000000000000000000010000;
		2988: Delta = 69'sb111111111111111111111100000000000000000000000000000000000000000010000;
		47873: Delta = 69'sb000000000000000000000011111111111111111111111111111111111111111110000;
		2956: Delta = 69'sb111111111111111111111011111111111111111111111111111111111111111110000;
		44933: Delta = 69'sb000000000000000000001000000000000000000000000000000000000000000010000;
		5960: Delta = 69'sb111111111111111111111000000000000000000000000000000000000000000010000;
		44901: Delta = 69'sb000000000000000000000111111111111111111111111111111111111111111110000;
		5928: Delta = 69'sb111111111111111111110111111111111111111111111111111111111111111110000;
		38989: Delta = 69'sb000000000000000000010000000000000000000000000000000000000000000010000;
		11904: Delta = 69'sb111111111111111111110000000000000000000000000000000000000000000010000;
		38957: Delta = 69'sb000000000000000000001111111111111111111111111111111111111111111110000;
		11872: Delta = 69'sb111111111111111111101111111111111111111111111111111111111111111110000;
		27101: Delta = 69'sb000000000000000000100000000000000000000000000000000000000000000010000;
		23792: Delta = 69'sb111111111111111111100000000000000000000000000000000000000000000010000;
		27069: Delta = 69'sb000000000000000000011111111111111111111111111111111111111111111110000;
		23760: Delta = 69'sb111111111111111111011111111111111111111111111111111111111111111110000;
		3325: Delta = 69'sb000000000000000001000000000000000000000000000000000000000000000010000;
		47568: Delta = 69'sb111111111111111111000000000000000000000000000000000000000000000010000;
		3293: Delta = 69'sb000000000000000000111111111111111111111111111111111111111111111110000;
		47536: Delta = 69'sb111111111111111110111111111111111111111111111111111111111111111110000;
		6634: Delta = 69'sb000000000000000010000000000000000000000000000000000000000000000010000;
		44259: Delta = 69'sb111111111111111110000000000000000000000000000000000000000000000010000;
		6602: Delta = 69'sb000000000000000001111111111111111111111111111111111111111111111110000;
		44227: Delta = 69'sb111111111111111101111111111111111111111111111111111111111111111110000;
		13252: Delta = 69'sb000000000000000100000000000000000000000000000000000000000000000010000;
		37641: Delta = 69'sb111111111111111100000000000000000000000000000000000000000000000010000;
		13220: Delta = 69'sb000000000000000011111111111111111111111111111111111111111111111110000;
		37609: Delta = 69'sb111111111111111011111111111111111111111111111111111111111111111110000;
		26488: Delta = 69'sb000000000000001000000000000000000000000000000000000000000000000010000;
		24405: Delta = 69'sb111111111111111000000000000000000000000000000000000000000000000010000;
		26456: Delta = 69'sb000000000000000111111111111111111111111111111111111111111111111110000;
		24373: Delta = 69'sb111111111111110111111111111111111111111111111111111111111111111110000;
		2099: Delta = 69'sb000000000000010000000000000000000000000000000000000000000000000010000;
		48794: Delta = 69'sb111111111111110000000000000000000000000000000000000000000000000010000;
		2067: Delta = 69'sb000000000000001111111111111111111111111111111111111111111111111110000;
		48762: Delta = 69'sb111111111111101111111111111111111111111111111111111111111111111110000;
		4182: Delta = 69'sb000000000000100000000000000000000000000000000000000000000000000010000;
		46711: Delta = 69'sb111111111111100000000000000000000000000000000000000000000000000010000;
		4150: Delta = 69'sb000000000000011111111111111111111111111111111111111111111111111110000;
		46679: Delta = 69'sb111111111111011111111111111111111111111111111111111111111111111110000;
		8348: Delta = 69'sb000000000001000000000000000000000000000000000000000000000000000010000;
		42545: Delta = 69'sb111111111111000000000000000000000000000000000000000000000000000010000;
		8316: Delta = 69'sb000000000000111111111111111111111111111111111111111111111111111110000;
		42513: Delta = 69'sb111111111110111111111111111111111111111111111111111111111111111110000;
		16680: Delta = 69'sb000000000010000000000000000000000000000000000000000000000000000010000;
		34213: Delta = 69'sb111111111110000000000000000000000000000000000000000000000000000010000;
		16648: Delta = 69'sb000000000001111111111111111111111111111111111111111111111111111110000;
		34181: Delta = 69'sb111111111101111111111111111111111111111111111111111111111111111110000;
		33344: Delta = 69'sb000000000100000000000000000000000000000000000000000000000000000010000;
		17549: Delta = 69'sb111111111100000000000000000000000000000000000000000000000000000010000;
		33312: Delta = 69'sb000000000011111111111111111111111111111111111111111111111111111110000;
		17517: Delta = 69'sb111111111011111111111111111111111111111111111111111111111111111110000;
		15811: Delta = 69'sb000000001000000000000000000000000000000000000000000000000000000010000;
		35082: Delta = 69'sb111111111000000000000000000000000000000000000000000000000000000010000;
		15779: Delta = 69'sb000000000111111111111111111111111111111111111111111111111111111110000;
		35050: Delta = 69'sb111111110111111111111111111111111111111111111111111111111111111110000;
		31606: Delta = 69'sb000000010000000000000000000000000000000000000000000000000000000010000;
		19287: Delta = 69'sb111111110000000000000000000000000000000000000000000000000000000010000;
		31574: Delta = 69'sb000000001111111111111111111111111111111111111111111111111111111110000;
		19255: Delta = 69'sb111111101111111111111111111111111111111111111111111111111111111110000;
		12335: Delta = 69'sb000000100000000000000000000000000000000000000000000000000000000010000;
		38558: Delta = 69'sb111111100000000000000000000000000000000000000000000000000000000010000;
		12303: Delta = 69'sb000000011111111111111111111111111111111111111111111111111111111110000;
		38526: Delta = 69'sb111111011111111111111111111111111111111111111111111111111111111110000;
		24654: Delta = 69'sb000001000000000000000000000000000000000000000000000000000000000010000;
		26239: Delta = 69'sb111111000000000000000000000000000000000000000000000000000000000010000;
		24622: Delta = 69'sb000000111111111111111111111111111111111111111111111111111111111110000;
		26207: Delta = 69'sb111110111111111111111111111111111111111111111111111111111111111110000;
		49292: Delta = 69'sb000010000000000000000000000000000000000000000000000000000000000010000;
		1601: Delta = 69'sb111110000000000000000000000000000000000000000000000000000000000010000;
		49260: Delta = 69'sb000001111111111111111111111111111111111111111111111111111111111110000;
		1569: Delta = 69'sb111101111111111111111111111111111111111111111111111111111111111110000;
		47707: Delta = 69'sb000100000000000000000000000000000000000000000000000000000000000010000;
		3186: Delta = 69'sb111100000000000000000000000000000000000000000000000000000000000010000;
		47675: Delta = 69'sb000011111111111111111111111111111111111111111111111111111111111110000;
		3154: Delta = 69'sb111011111111111111111111111111111111111111111111111111111111111110000;
		44537: Delta = 69'sb001000000000000000000000000000000000000000000000000000000000000010000;
		6356: Delta = 69'sb111000000000000000000000000000000000000000000000000000000000000010000;
		44505: Delta = 69'sb000111111111111111111111111111111111111111111111111111111111111110000;
		6324: Delta = 69'sb110111111111111111111111111111111111111111111111111111111111111110000;
		38197: Delta = 69'sb010000000000000000000000000000000000000000000000000000000000000010000;
		12696: Delta = 69'sb110000000000000000000000000000000000000000000000000000000000000010000;
		38165: Delta = 69'sb001111111111111111111111111111111111111111111111111111111111111110000;
		12664: Delta = 69'sb101111111111111111111111111111111111111111111111111111111111111110000;
		96: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000001100000;
		50765: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111110100000;
		160: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000010100000;
		50701: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111101100000;
		288: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000100100000;
		50637: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111100100000;
		224: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000011100000;
		50573: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111011100000;
		544: Delta = 69'sb000000000000000000000000000000000000000000000000000000000001000100000;
		50381: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111000100000;
		480: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000111100000;
		50317: Delta = 69'sb111111111111111111111111111111111111111111111111111111111110111100000;
		1056: Delta = 69'sb000000000000000000000000000000000000000000000000000000000010000100000;
		49869: Delta = 69'sb111111111111111111111111111111111111111111111111111111111110000100000;
		992: Delta = 69'sb000000000000000000000000000000000000000000000000000000000001111100000;
		49805: Delta = 69'sb111111111111111111111111111111111111111111111111111111111101111100000;
		2080: Delta = 69'sb000000000000000000000000000000000000000000000000000000000100000100000;
		48845: Delta = 69'sb111111111111111111111111111111111111111111111111111111111100000100000;
		2016: Delta = 69'sb000000000000000000000000000000000000000000000000000000000011111100000;
		48781: Delta = 69'sb111111111111111111111111111111111111111111111111111111111011111100000;
		4128: Delta = 69'sb000000000000000000000000000000000000000000000000000000001000000100000;
		46797: Delta = 69'sb111111111111111111111111111111111111111111111111111111111000000100000;
		4064: Delta = 69'sb000000000000000000000000000000000000000000000000000000000111111100000;
		46733: Delta = 69'sb111111111111111111111111111111111111111111111111111111110111111100000;
		8224: Delta = 69'sb000000000000000000000000000000000000000000000000000000010000000100000;
		42701: Delta = 69'sb111111111111111111111111111111111111111111111111111111110000000100000;
		8160: Delta = 69'sb000000000000000000000000000000000000000000000000000000001111111100000;
		42637: Delta = 69'sb111111111111111111111111111111111111111111111111111111101111111100000;
		16416: Delta = 69'sb000000000000000000000000000000000000000000000000000000100000000100000;
		34509: Delta = 69'sb111111111111111111111111111111111111111111111111111111100000000100000;
		16352: Delta = 69'sb000000000000000000000000000000000000000000000000000000011111111100000;
		34445: Delta = 69'sb111111111111111111111111111111111111111111111111111111011111111100000;
		32800: Delta = 69'sb000000000000000000000000000000000000000000000000000001000000000100000;
		18125: Delta = 69'sb111111111111111111111111111111111111111111111111111111000000000100000;
		32736: Delta = 69'sb000000000000000000000000000000000000000000000000000000111111111100000;
		18061: Delta = 69'sb111111111111111111111111111111111111111111111111111110111111111100000;
		14707: Delta = 69'sb000000000000000000000000000000000000000000000000000010000000000100000;
		36218: Delta = 69'sb111111111111111111111111111111111111111111111111111110000000000100000;
		14643: Delta = 69'sb000000000000000000000000000000000000000000000000000001111111111100000;
		36154: Delta = 69'sb111111111111111111111111111111111111111111111111111101111111111100000;
		29382: Delta = 69'sb000000000000000000000000000000000000000000000000000100000000000100000;
		21543: Delta = 69'sb111111111111111111111111111111111111111111111111111100000000000100000;
		29318: Delta = 69'sb000000000000000000000000000000000000000000000000000011111111111100000;
		21479: Delta = 69'sb111111111111111111111111111111111111111111111111111011111111111100000;
		7871: Delta = 69'sb000000000000000000000000000000000000000000000000001000000000000100000;
		43054: Delta = 69'sb111111111111111111111111111111111111111111111111111000000000000100000;
		7807: Delta = 69'sb000000000000000000000000000000000000000000000000000111111111111100000;
		42990: Delta = 69'sb111111111111111111111111111111111111111111111111110111111111111100000;
		15710: Delta = 69'sb000000000000000000000000000000000000000000000000010000000000000100000;
		35215: Delta = 69'sb111111111111111111111111111111111111111111111111110000000000000100000;
		15646: Delta = 69'sb000000000000000000000000000000000000000000000000001111111111111100000;
		35151: Delta = 69'sb111111111111111111111111111111111111111111111111101111111111111100000;
		31388: Delta = 69'sb000000000000000000000000000000000000000000000000100000000000000100000;
		19537: Delta = 69'sb111111111111111111111111111111111111111111111111100000000000000100000;
		31324: Delta = 69'sb000000000000000000000000000000000000000000000000011111111111111100000;
		19473: Delta = 69'sb111111111111111111111111111111111111111111111111011111111111111100000;
		11883: Delta = 69'sb000000000000000000000000000000000000000000000001000000000000000100000;
		39042: Delta = 69'sb111111111111111111111111111111111111111111111111000000000000000100000;
		11819: Delta = 69'sb000000000000000000000000000000000000000000000000111111111111111100000;
		38978: Delta = 69'sb111111111111111111111111111111111111111111111110111111111111111100000;
		23734: Delta = 69'sb000000000000000000000000000000000000000000000010000000000000000100000;
		27191: Delta = 69'sb111111111111111111111111111111111111111111111110000000000000000100000;
		23670: Delta = 69'sb000000000000000000000000000000000000000000000001111111111111111100000;
		27127: Delta = 69'sb111111111111111111111111111111111111111111111101111111111111111100000;
		47436: Delta = 69'sb000000000000000000000000000000000000000000000100000000000000000100000;
		3489: Delta = 69'sb111111111111111111111111111111111111111111111100000000000000000100000;
		47372: Delta = 69'sb000000000000000000000000000000000000000000000011111111111111111100000;
		3425: Delta = 69'sb111111111111111111111111111111111111111111111011111111111111111100000;
		43979: Delta = 69'sb000000000000000000000000000000000000000000001000000000000000000100000;
		6946: Delta = 69'sb111111111111111111111111111111111111111111111000000000000000000100000;
		43915: Delta = 69'sb000000000000000000000000000000000000000000000111111111111111111100000;
		6882: Delta = 69'sb111111111111111111111111111111111111111111110111111111111111111100000;
		37065: Delta = 69'sb000000000000000000000000000000000000000000010000000000000000000100000;
		13860: Delta = 69'sb111111111111111111111111111111111111111111110000000000000000000100000;
		37001: Delta = 69'sb000000000000000000000000000000000000000000001111111111111111111100000;
		13796: Delta = 69'sb111111111111111111111111111111111111111111101111111111111111111100000;
		23237: Delta = 69'sb000000000000000000000000000000000000000000100000000000000000000100000;
		27688: Delta = 69'sb111111111111111111111111111111111111111111100000000000000000000100000;
		23173: Delta = 69'sb000000000000000000000000000000000000000000011111111111111111111100000;
		27624: Delta = 69'sb111111111111111111111111111111111111111111011111111111111111111100000;
		46442: Delta = 69'sb000000000000000000000000000000000000000001000000000000000000000100000;
		4483: Delta = 69'sb111111111111111111111111111111111111111111000000000000000000000100000;
		46378: Delta = 69'sb000000000000000000000000000000000000000000111111111111111111111100000;
		4419: Delta = 69'sb111111111111111111111111111111111111111110111111111111111111111100000;
		41991: Delta = 69'sb000000000000000000000000000000000000000010000000000000000000000100000;
		8934: Delta = 69'sb111111111111111111111111111111111111111110000000000000000000000100000;
		41927: Delta = 69'sb000000000000000000000000000000000000000001111111111111111111111100000;
		8870: Delta = 69'sb111111111111111111111111111111111111111101111111111111111111111100000;
		33089: Delta = 69'sb000000000000000000000000000000000000000100000000000000000000000100000;
		17836: Delta = 69'sb111111111111111111111111111111111111111100000000000000000000000100000;
		33025: Delta = 69'sb000000000000000000000000000000000000000011111111111111111111111100000;
		17772: Delta = 69'sb111111111111111111111111111111111111111011111111111111111111111100000;
		15285: Delta = 69'sb000000000000000000000000000000000000001000000000000000000000000100000;
		35640: Delta = 69'sb111111111111111111111111111111111111111000000000000000000000000100000;
		15221: Delta = 69'sb000000000000000000000000000000000000000111111111111111111111111100000;
		35576: Delta = 69'sb111111111111111111111111111111111111110111111111111111111111111100000;
		30538: Delta = 69'sb000000000000000000000000000000000000010000000000000000000000000100000;
		20387: Delta = 69'sb111111111111111111111111111111111111110000000000000000000000000100000;
		30474: Delta = 69'sb000000000000000000000000000000000000001111111111111111111111111100000;
		20323: Delta = 69'sb111111111111111111111111111111111111101111111111111111111111111100000;
		10183: Delta = 69'sb000000000000000000000000000000000000100000000000000000000000000100000;
		40742: Delta = 69'sb111111111111111111111111111111111111100000000000000000000000000100000;
		10119: Delta = 69'sb000000000000000000000000000000000000011111111111111111111111111100000;
		40678: Delta = 69'sb111111111111111111111111111111111111011111111111111111111111111100000;
		20334: Delta = 69'sb000000000000000000000000000000000001000000000000000000000000000100000;
		30591: Delta = 69'sb111111111111111111111111111111111111000000000000000000000000000100000;
		20270: Delta = 69'sb000000000000000000000000000000000000111111111111111111111111111100000;
		30527: Delta = 69'sb111111111111111111111111111111111110111111111111111111111111111100000;
		40636: Delta = 69'sb000000000000000000000000000000000010000000000000000000000000000100000;
		10289: Delta = 69'sb111111111111111111111111111111111110000000000000000000000000000100000;
		40572: Delta = 69'sb000000000000000000000000000000000001111111111111111111111111111100000;
		10225: Delta = 69'sb111111111111111111111111111111111101111111111111111111111111111100000;
		30379: Delta = 69'sb000000000000000000000000000000000100000000000000000000000000000100000;
		20546: Delta = 69'sb111111111111111111111111111111111100000000000000000000000000000100000;
		30315: Delta = 69'sb000000000000000000000000000000000011111111111111111111111111111100000;
		20482: Delta = 69'sb111111111111111111111111111111111011111111111111111111111111111100000;
		9865: Delta = 69'sb000000000000000000000000000000001000000000000000000000000000000100000;
		41060: Delta = 69'sb111111111111111111111111111111111000000000000000000000000000000100000;
		9801: Delta = 69'sb000000000000000000000000000000000111111111111111111111111111111100000;
		40996: Delta = 69'sb111111111111111111111111111111110111111111111111111111111111111100000;
		19698: Delta = 69'sb000000000000000000000000000000010000000000000000000000000000000100000;
		31227: Delta = 69'sb111111111111111111111111111111110000000000000000000000000000000100000;
		19634: Delta = 69'sb000000000000000000000000000000001111111111111111111111111111111100000;
		31163: Delta = 69'sb111111111111111111111111111111101111111111111111111111111111111100000;
		39364: Delta = 69'sb000000000000000000000000000000100000000000000000000000000000000100000;
		11561: Delta = 69'sb111111111111111111111111111111100000000000000000000000000000000100000;
		39300: Delta = 69'sb000000000000000000000000000000011111111111111111111111111111111100000;
		11497: Delta = 69'sb111111111111111111111111111111011111111111111111111111111111111100000;
		27835: Delta = 69'sb000000000000000000000000000001000000000000000000000000000000000100000;
		23090: Delta = 69'sb111111111111111111111111111111000000000000000000000000000000000100000;
		27771: Delta = 69'sb000000000000000000000000000000111111111111111111111111111111111100000;
		23026: Delta = 69'sb111111111111111111111111111110111111111111111111111111111111111100000;
		4777: Delta = 69'sb000000000000000000000000000010000000000000000000000000000000000100000;
		46148: Delta = 69'sb111111111111111111111111111110000000000000000000000000000000000100000;
		4713: Delta = 69'sb000000000000000000000000000001111111111111111111111111111111111100000;
		46084: Delta = 69'sb111111111111111111111111111101111111111111111111111111111111111100000;
		9522: Delta = 69'sb000000000000000000000000000100000000000000000000000000000000000100000;
		41403: Delta = 69'sb111111111111111111111111111100000000000000000000000000000000000100000;
		9458: Delta = 69'sb000000000000000000000000000011111111111111111111111111111111111100000;
		41339: Delta = 69'sb111111111111111111111111111011111111111111111111111111111111111100000;
		19012: Delta = 69'sb000000000000000000000000001000000000000000000000000000000000000100000;
		31913: Delta = 69'sb111111111111111111111111111000000000000000000000000000000000000100000;
		18948: Delta = 69'sb000000000000000000000000000111111111111111111111111111111111111100000;
		31849: Delta = 69'sb111111111111111111111111110111111111111111111111111111111111111100000;
		37992: Delta = 69'sb000000000000000000000000010000000000000000000000000000000000000100000;
		12933: Delta = 69'sb111111111111111111111111110000000000000000000000000000000000000100000;
		37928: Delta = 69'sb000000000000000000000000001111111111111111111111111111111111111100000;
		12869: Delta = 69'sb111111111111111111111111101111111111111111111111111111111111111100000;
		25091: Delta = 69'sb000000000000000000000000100000000000000000000000000000000000000100000;
		25834: Delta = 69'sb111111111111111111111111100000000000000000000000000000000000000100000;
		25027: Delta = 69'sb000000000000000000000000011111111111111111111111111111111111111100000;
		25770: Delta = 69'sb111111111111111111111111011111111111111111111111111111111111111100000;
		50150: Delta = 69'sb000000000000000000000001000000000000000000000000000000000000000100000;
		775: Delta = 69'sb111111111111111111111111000000000000000000000000000000000000000100000;
		50086: Delta = 69'sb000000000000000000000000111111111111111111111111111111111111111100000;
		711: Delta = 69'sb111111111111111111111110111111111111111111111111111111111111111100000;
		49407: Delta = 69'sb000000000000000000000010000000000000000000000000000000000000000100000;
		1518: Delta = 69'sb111111111111111111111110000000000000000000000000000000000000000100000;
		49343: Delta = 69'sb000000000000000000000001111111111111111111111111111111111111111100000;
		1454: Delta = 69'sb111111111111111111111101111111111111111111111111111111111111111100000;
		47921: Delta = 69'sb000000000000000000000100000000000000000000000000000000000000000100000;
		3004: Delta = 69'sb111111111111111111111100000000000000000000000000000000000000000100000;
		47857: Delta = 69'sb000000000000000000000011111111111111111111111111111111111111111100000;
		2940: Delta = 69'sb111111111111111111111011111111111111111111111111111111111111111100000;
		44949: Delta = 69'sb000000000000000000001000000000000000000000000000000000000000000100000;
		5976: Delta = 69'sb111111111111111111111000000000000000000000000000000000000000000100000;
		44885: Delta = 69'sb000000000000000000000111111111111111111111111111111111111111111100000;
		5912: Delta = 69'sb111111111111111111110111111111111111111111111111111111111111111100000;
		39005: Delta = 69'sb000000000000000000010000000000000000000000000000000000000000000100000;
		11920: Delta = 69'sb111111111111111111110000000000000000000000000000000000000000000100000;
		38941: Delta = 69'sb000000000000000000001111111111111111111111111111111111111111111100000;
		11856: Delta = 69'sb111111111111111111101111111111111111111111111111111111111111111100000;
		27117: Delta = 69'sb000000000000000000100000000000000000000000000000000000000000000100000;
		23808: Delta = 69'sb111111111111111111100000000000000000000000000000000000000000000100000;
		27053: Delta = 69'sb000000000000000000011111111111111111111111111111111111111111111100000;
		23744: Delta = 69'sb111111111111111111011111111111111111111111111111111111111111111100000;
		3341: Delta = 69'sb000000000000000001000000000000000000000000000000000000000000000100000;
		47584: Delta = 69'sb111111111111111111000000000000000000000000000000000000000000000100000;
		3277: Delta = 69'sb000000000000000000111111111111111111111111111111111111111111111100000;
		47520: Delta = 69'sb111111111111111110111111111111111111111111111111111111111111111100000;
		6650: Delta = 69'sb000000000000000010000000000000000000000000000000000000000000000100000;
		44275: Delta = 69'sb111111111111111110000000000000000000000000000000000000000000000100000;
		6586: Delta = 69'sb000000000000000001111111111111111111111111111111111111111111111100000;
		44211: Delta = 69'sb111111111111111101111111111111111111111111111111111111111111111100000;
		13268: Delta = 69'sb000000000000000100000000000000000000000000000000000000000000000100000;
		37657: Delta = 69'sb111111111111111100000000000000000000000000000000000000000000000100000;
		13204: Delta = 69'sb000000000000000011111111111111111111111111111111111111111111111100000;
		37593: Delta = 69'sb111111111111111011111111111111111111111111111111111111111111111100000;
		26504: Delta = 69'sb000000000000001000000000000000000000000000000000000000000000000100000;
		24421: Delta = 69'sb111111111111111000000000000000000000000000000000000000000000000100000;
		26440: Delta = 69'sb000000000000000111111111111111111111111111111111111111111111111100000;
		24357: Delta = 69'sb111111111111110111111111111111111111111111111111111111111111111100000;
		2115: Delta = 69'sb000000000000010000000000000000000000000000000000000000000000000100000;
		48810: Delta = 69'sb111111111111110000000000000000000000000000000000000000000000000100000;
		2051: Delta = 69'sb000000000000001111111111111111111111111111111111111111111111111100000;
		48746: Delta = 69'sb111111111111101111111111111111111111111111111111111111111111111100000;
		4198: Delta = 69'sb000000000000100000000000000000000000000000000000000000000000000100000;
		46727: Delta = 69'sb111111111111100000000000000000000000000000000000000000000000000100000;
		4134: Delta = 69'sb000000000000011111111111111111111111111111111111111111111111111100000;
		46663: Delta = 69'sb111111111111011111111111111111111111111111111111111111111111111100000;
		8364: Delta = 69'sb000000000001000000000000000000000000000000000000000000000000000100000;
		42561: Delta = 69'sb111111111111000000000000000000000000000000000000000000000000000100000;
		8300: Delta = 69'sb000000000000111111111111111111111111111111111111111111111111111100000;
		42497: Delta = 69'sb111111111110111111111111111111111111111111111111111111111111111100000;
		16696: Delta = 69'sb000000000010000000000000000000000000000000000000000000000000000100000;
		34229: Delta = 69'sb111111111110000000000000000000000000000000000000000000000000000100000;
		16632: Delta = 69'sb000000000001111111111111111111111111111111111111111111111111111100000;
		34165: Delta = 69'sb111111111101111111111111111111111111111111111111111111111111111100000;
		33360: Delta = 69'sb000000000100000000000000000000000000000000000000000000000000000100000;
		17565: Delta = 69'sb111111111100000000000000000000000000000000000000000000000000000100000;
		33296: Delta = 69'sb000000000011111111111111111111111111111111111111111111111111111100000;
		17501: Delta = 69'sb111111111011111111111111111111111111111111111111111111111111111100000;
		15827: Delta = 69'sb000000001000000000000000000000000000000000000000000000000000000100000;
		35098: Delta = 69'sb111111111000000000000000000000000000000000000000000000000000000100000;
		15763: Delta = 69'sb000000000111111111111111111111111111111111111111111111111111111100000;
		35034: Delta = 69'sb111111110111111111111111111111111111111111111111111111111111111100000;
		31622: Delta = 69'sb000000010000000000000000000000000000000000000000000000000000000100000;
		19303: Delta = 69'sb111111110000000000000000000000000000000000000000000000000000000100000;
		31558: Delta = 69'sb000000001111111111111111111111111111111111111111111111111111111100000;
		19239: Delta = 69'sb111111101111111111111111111111111111111111111111111111111111111100000;
		12351: Delta = 69'sb000000100000000000000000000000000000000000000000000000000000000100000;
		38574: Delta = 69'sb111111100000000000000000000000000000000000000000000000000000000100000;
		12287: Delta = 69'sb000000011111111111111111111111111111111111111111111111111111111100000;
		38510: Delta = 69'sb111111011111111111111111111111111111111111111111111111111111111100000;
		24670: Delta = 69'sb000001000000000000000000000000000000000000000000000000000000000100000;
		26255: Delta = 69'sb111111000000000000000000000000000000000000000000000000000000000100000;
		24606: Delta = 69'sb000000111111111111111111111111111111111111111111111111111111111100000;
		26191: Delta = 69'sb111110111111111111111111111111111111111111111111111111111111111100000;
		49308: Delta = 69'sb000010000000000000000000000000000000000000000000000000000000000100000;
		1617: Delta = 69'sb111110000000000000000000000000000000000000000000000000000000000100000;
		49244: Delta = 69'sb000001111111111111111111111111111111111111111111111111111111111100000;
		1553: Delta = 69'sb111101111111111111111111111111111111111111111111111111111111111100000;
		47723: Delta = 69'sb000100000000000000000000000000000000000000000000000000000000000100000;
		3202: Delta = 69'sb111100000000000000000000000000000000000000000000000000000000000100000;
		47659: Delta = 69'sb000011111111111111111111111111111111111111111111111111111111111100000;
		3138: Delta = 69'sb111011111111111111111111111111111111111111111111111111111111111100000;
		44553: Delta = 69'sb001000000000000000000000000000000000000000000000000000000000000100000;
		6372: Delta = 69'sb111000000000000000000000000000000000000000000000000000000000000100000;
		44489: Delta = 69'sb000111111111111111111111111111111111111111111111111111111111111100000;
		6308: Delta = 69'sb110111111111111111111111111111111111111111111111111111111111111100000;
		38213: Delta = 69'sb010000000000000000000000000000000000000000000000000000000000000100000;
		12712: Delta = 69'sb110000000000000000000000000000000000000000000000000000000000000100000;
		38149: Delta = 69'sb001111111111111111111111111111111111111111111111111111111111111100000;
		12648: Delta = 69'sb101111111111111111111111111111111111111111111111111111111111111100000;
		192: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000011000000;
		50669: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111101000000;
		320: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000101000000;
		50541: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111011000000;
		576: Delta = 69'sb000000000000000000000000000000000000000000000000000000000001001000000;
		50413: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111001000000;
		448: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000111000000;
		50285: Delta = 69'sb111111111111111111111111111111111111111111111111111111111110111000000;
		1088: Delta = 69'sb000000000000000000000000000000000000000000000000000000000010001000000;
		49901: Delta = 69'sb111111111111111111111111111111111111111111111111111111111110001000000;
		960: Delta = 69'sb000000000000000000000000000000000000000000000000000000000001111000000;
		49773: Delta = 69'sb111111111111111111111111111111111111111111111111111111111101111000000;
		2112: Delta = 69'sb000000000000000000000000000000000000000000000000000000000100001000000;
		48877: Delta = 69'sb111111111111111111111111111111111111111111111111111111111100001000000;
		1984: Delta = 69'sb000000000000000000000000000000000000000000000000000000000011111000000;
		48749: Delta = 69'sb111111111111111111111111111111111111111111111111111111111011111000000;
		4160: Delta = 69'sb000000000000000000000000000000000000000000000000000000001000001000000;
		46829: Delta = 69'sb111111111111111111111111111111111111111111111111111111111000001000000;
		4032: Delta = 69'sb000000000000000000000000000000000000000000000000000000000111111000000;
		46701: Delta = 69'sb111111111111111111111111111111111111111111111111111111110111111000000;
		8256: Delta = 69'sb000000000000000000000000000000000000000000000000000000010000001000000;
		42733: Delta = 69'sb111111111111111111111111111111111111111111111111111111110000001000000;
		8128: Delta = 69'sb000000000000000000000000000000000000000000000000000000001111111000000;
		42605: Delta = 69'sb111111111111111111111111111111111111111111111111111111101111111000000;
		16448: Delta = 69'sb000000000000000000000000000000000000000000000000000000100000001000000;
		34541: Delta = 69'sb111111111111111111111111111111111111111111111111111111100000001000000;
		16320: Delta = 69'sb000000000000000000000000000000000000000000000000000000011111111000000;
		34413: Delta = 69'sb111111111111111111111111111111111111111111111111111111011111111000000;
		32832: Delta = 69'sb000000000000000000000000000000000000000000000000000001000000001000000;
		18157: Delta = 69'sb111111111111111111111111111111111111111111111111111111000000001000000;
		32704: Delta = 69'sb000000000000000000000000000000000000000000000000000000111111111000000;
		18029: Delta = 69'sb111111111111111111111111111111111111111111111111111110111111111000000;
		14739: Delta = 69'sb000000000000000000000000000000000000000000000000000010000000001000000;
		36250: Delta = 69'sb111111111111111111111111111111111111111111111111111110000000001000000;
		14611: Delta = 69'sb000000000000000000000000000000000000000000000000000001111111111000000;
		36122: Delta = 69'sb111111111111111111111111111111111111111111111111111101111111111000000;
		29414: Delta = 69'sb000000000000000000000000000000000000000000000000000100000000001000000;
		21575: Delta = 69'sb111111111111111111111111111111111111111111111111111100000000001000000;
		29286: Delta = 69'sb000000000000000000000000000000000000000000000000000011111111111000000;
		21447: Delta = 69'sb111111111111111111111111111111111111111111111111111011111111111000000;
		7903: Delta = 69'sb000000000000000000000000000000000000000000000000001000000000001000000;
		43086: Delta = 69'sb111111111111111111111111111111111111111111111111111000000000001000000;
		7775: Delta = 69'sb000000000000000000000000000000000000000000000000000111111111111000000;
		42958: Delta = 69'sb111111111111111111111111111111111111111111111111110111111111111000000;
		15742: Delta = 69'sb000000000000000000000000000000000000000000000000010000000000001000000;
		35247: Delta = 69'sb111111111111111111111111111111111111111111111111110000000000001000000;
		15614: Delta = 69'sb000000000000000000000000000000000000000000000000001111111111111000000;
		35119: Delta = 69'sb111111111111111111111111111111111111111111111111101111111111111000000;
		31420: Delta = 69'sb000000000000000000000000000000000000000000000000100000000000001000000;
		19569: Delta = 69'sb111111111111111111111111111111111111111111111111100000000000001000000;
		31292: Delta = 69'sb000000000000000000000000000000000000000000000000011111111111111000000;
		19441: Delta = 69'sb111111111111111111111111111111111111111111111111011111111111111000000;
		11915: Delta = 69'sb000000000000000000000000000000000000000000000001000000000000001000000;
		39074: Delta = 69'sb111111111111111111111111111111111111111111111111000000000000001000000;
		11787: Delta = 69'sb000000000000000000000000000000000000000000000000111111111111111000000;
		38946: Delta = 69'sb111111111111111111111111111111111111111111111110111111111111111000000;
		23766: Delta = 69'sb000000000000000000000000000000000000000000000010000000000000001000000;
		27223: Delta = 69'sb111111111111111111111111111111111111111111111110000000000000001000000;
		23638: Delta = 69'sb000000000000000000000000000000000000000000000001111111111111111000000;
		27095: Delta = 69'sb111111111111111111111111111111111111111111111101111111111111111000000;
		47468: Delta = 69'sb000000000000000000000000000000000000000000000100000000000000001000000;
		3521: Delta = 69'sb111111111111111111111111111111111111111111111100000000000000001000000;
		47340: Delta = 69'sb000000000000000000000000000000000000000000000011111111111111111000000;
		3393: Delta = 69'sb111111111111111111111111111111111111111111111011111111111111111000000;
		44011: Delta = 69'sb000000000000000000000000000000000000000000001000000000000000001000000;
		6978: Delta = 69'sb111111111111111111111111111111111111111111111000000000000000001000000;
		43883: Delta = 69'sb000000000000000000000000000000000000000000000111111111111111111000000;
		6850: Delta = 69'sb111111111111111111111111111111111111111111110111111111111111111000000;
		37097: Delta = 69'sb000000000000000000000000000000000000000000010000000000000000001000000;
		13892: Delta = 69'sb111111111111111111111111111111111111111111110000000000000000001000000;
		36969: Delta = 69'sb000000000000000000000000000000000000000000001111111111111111111000000;
		13764: Delta = 69'sb111111111111111111111111111111111111111111101111111111111111111000000;
		23269: Delta = 69'sb000000000000000000000000000000000000000000100000000000000000001000000;
		27720: Delta = 69'sb111111111111111111111111111111111111111111100000000000000000001000000;
		23141: Delta = 69'sb000000000000000000000000000000000000000000011111111111111111111000000;
		27592: Delta = 69'sb111111111111111111111111111111111111111111011111111111111111111000000;
		46474: Delta = 69'sb000000000000000000000000000000000000000001000000000000000000001000000;
		4515: Delta = 69'sb111111111111111111111111111111111111111111000000000000000000001000000;
		46346: Delta = 69'sb000000000000000000000000000000000000000000111111111111111111111000000;
		4387: Delta = 69'sb111111111111111111111111111111111111111110111111111111111111111000000;
		42023: Delta = 69'sb000000000000000000000000000000000000000010000000000000000000001000000;
		8966: Delta = 69'sb111111111111111111111111111111111111111110000000000000000000001000000;
		41895: Delta = 69'sb000000000000000000000000000000000000000001111111111111111111111000000;
		8838: Delta = 69'sb111111111111111111111111111111111111111101111111111111111111111000000;
		33121: Delta = 69'sb000000000000000000000000000000000000000100000000000000000000001000000;
		17868: Delta = 69'sb111111111111111111111111111111111111111100000000000000000000001000000;
		32993: Delta = 69'sb000000000000000000000000000000000000000011111111111111111111111000000;
		17740: Delta = 69'sb111111111111111111111111111111111111111011111111111111111111111000000;
		15317: Delta = 69'sb000000000000000000000000000000000000001000000000000000000000001000000;
		35672: Delta = 69'sb111111111111111111111111111111111111111000000000000000000000001000000;
		15189: Delta = 69'sb000000000000000000000000000000000000000111111111111111111111111000000;
		35544: Delta = 69'sb111111111111111111111111111111111111110111111111111111111111111000000;
		30570: Delta = 69'sb000000000000000000000000000000000000010000000000000000000000001000000;
		20419: Delta = 69'sb111111111111111111111111111111111111110000000000000000000000001000000;
		30442: Delta = 69'sb000000000000000000000000000000000000001111111111111111111111111000000;
		20291: Delta = 69'sb111111111111111111111111111111111111101111111111111111111111111000000;
		10215: Delta = 69'sb000000000000000000000000000000000000100000000000000000000000001000000;
		40774: Delta = 69'sb111111111111111111111111111111111111100000000000000000000000001000000;
		10087: Delta = 69'sb000000000000000000000000000000000000011111111111111111111111111000000;
		40646: Delta = 69'sb111111111111111111111111111111111111011111111111111111111111111000000;
		20366: Delta = 69'sb000000000000000000000000000000000001000000000000000000000000001000000;
		30623: Delta = 69'sb111111111111111111111111111111111111000000000000000000000000001000000;
		20238: Delta = 69'sb000000000000000000000000000000000000111111111111111111111111111000000;
		30495: Delta = 69'sb111111111111111111111111111111111110111111111111111111111111111000000;
		40668: Delta = 69'sb000000000000000000000000000000000010000000000000000000000000001000000;
		10321: Delta = 69'sb111111111111111111111111111111111110000000000000000000000000001000000;
		40540: Delta = 69'sb000000000000000000000000000000000001111111111111111111111111111000000;
		10193: Delta = 69'sb111111111111111111111111111111111101111111111111111111111111111000000;
		30411: Delta = 69'sb000000000000000000000000000000000100000000000000000000000000001000000;
		20578: Delta = 69'sb111111111111111111111111111111111100000000000000000000000000001000000;
		30283: Delta = 69'sb000000000000000000000000000000000011111111111111111111111111111000000;
		20450: Delta = 69'sb111111111111111111111111111111111011111111111111111111111111111000000;
		9897: Delta = 69'sb000000000000000000000000000000001000000000000000000000000000001000000;
		41092: Delta = 69'sb111111111111111111111111111111111000000000000000000000000000001000000;
		9769: Delta = 69'sb000000000000000000000000000000000111111111111111111111111111111000000;
		40964: Delta = 69'sb111111111111111111111111111111110111111111111111111111111111111000000;
		19730: Delta = 69'sb000000000000000000000000000000010000000000000000000000000000001000000;
		31259: Delta = 69'sb111111111111111111111111111111110000000000000000000000000000001000000;
		19602: Delta = 69'sb000000000000000000000000000000001111111111111111111111111111111000000;
		31131: Delta = 69'sb111111111111111111111111111111101111111111111111111111111111111000000;
		39396: Delta = 69'sb000000000000000000000000000000100000000000000000000000000000001000000;
		11593: Delta = 69'sb111111111111111111111111111111100000000000000000000000000000001000000;
		39268: Delta = 69'sb000000000000000000000000000000011111111111111111111111111111111000000;
		11465: Delta = 69'sb111111111111111111111111111111011111111111111111111111111111111000000;
		27867: Delta = 69'sb000000000000000000000000000001000000000000000000000000000000001000000;
		23122: Delta = 69'sb111111111111111111111111111111000000000000000000000000000000001000000;
		27739: Delta = 69'sb000000000000000000000000000000111111111111111111111111111111111000000;
		22994: Delta = 69'sb111111111111111111111111111110111111111111111111111111111111111000000;
		4809: Delta = 69'sb000000000000000000000000000010000000000000000000000000000000001000000;
		46180: Delta = 69'sb111111111111111111111111111110000000000000000000000000000000001000000;
		4681: Delta = 69'sb000000000000000000000000000001111111111111111111111111111111111000000;
		46052: Delta = 69'sb111111111111111111111111111101111111111111111111111111111111111000000;
		9554: Delta = 69'sb000000000000000000000000000100000000000000000000000000000000001000000;
		41435: Delta = 69'sb111111111111111111111111111100000000000000000000000000000000001000000;
		9426: Delta = 69'sb000000000000000000000000000011111111111111111111111111111111111000000;
		41307: Delta = 69'sb111111111111111111111111111011111111111111111111111111111111111000000;
		19044: Delta = 69'sb000000000000000000000000001000000000000000000000000000000000001000000;
		31945: Delta = 69'sb111111111111111111111111111000000000000000000000000000000000001000000;
		18916: Delta = 69'sb000000000000000000000000000111111111111111111111111111111111111000000;
		31817: Delta = 69'sb111111111111111111111111110111111111111111111111111111111111111000000;
		38024: Delta = 69'sb000000000000000000000000010000000000000000000000000000000000001000000;
		12965: Delta = 69'sb111111111111111111111111110000000000000000000000000000000000001000000;
		37896: Delta = 69'sb000000000000000000000000001111111111111111111111111111111111111000000;
		12837: Delta = 69'sb111111111111111111111111101111111111111111111111111111111111111000000;
		25123: Delta = 69'sb000000000000000000000000100000000000000000000000000000000000001000000;
		25866: Delta = 69'sb111111111111111111111111100000000000000000000000000000000000001000000;
		24995: Delta = 69'sb000000000000000000000000011111111111111111111111111111111111111000000;
		25738: Delta = 69'sb111111111111111111111111011111111111111111111111111111111111111000000;
		50182: Delta = 69'sb000000000000000000000001000000000000000000000000000000000000001000000;
		807: Delta = 69'sb111111111111111111111111000000000000000000000000000000000000001000000;
		50054: Delta = 69'sb000000000000000000000000111111111111111111111111111111111111111000000;
		679: Delta = 69'sb111111111111111111111110111111111111111111111111111111111111111000000;
		49439: Delta = 69'sb000000000000000000000010000000000000000000000000000000000000001000000;
		1550: Delta = 69'sb111111111111111111111110000000000000000000000000000000000000001000000;
		49311: Delta = 69'sb000000000000000000000001111111111111111111111111111111111111111000000;
		1422: Delta = 69'sb111111111111111111111101111111111111111111111111111111111111111000000;
		47953: Delta = 69'sb000000000000000000000100000000000000000000000000000000000000001000000;
		3036: Delta = 69'sb111111111111111111111100000000000000000000000000000000000000001000000;
		47825: Delta = 69'sb000000000000000000000011111111111111111111111111111111111111111000000;
		2908: Delta = 69'sb111111111111111111111011111111111111111111111111111111111111111000000;
		44981: Delta = 69'sb000000000000000000001000000000000000000000000000000000000000001000000;
		6008: Delta = 69'sb111111111111111111111000000000000000000000000000000000000000001000000;
		44853: Delta = 69'sb000000000000000000000111111111111111111111111111111111111111111000000;
		5880: Delta = 69'sb111111111111111111110111111111111111111111111111111111111111111000000;
		39037: Delta = 69'sb000000000000000000010000000000000000000000000000000000000000001000000;
		11952: Delta = 69'sb111111111111111111110000000000000000000000000000000000000000001000000;
		38909: Delta = 69'sb000000000000000000001111111111111111111111111111111111111111111000000;
		11824: Delta = 69'sb111111111111111111101111111111111111111111111111111111111111111000000;
		27149: Delta = 69'sb000000000000000000100000000000000000000000000000000000000000001000000;
		23840: Delta = 69'sb111111111111111111100000000000000000000000000000000000000000001000000;
		27021: Delta = 69'sb000000000000000000011111111111111111111111111111111111111111111000000;
		23712: Delta = 69'sb111111111111111111011111111111111111111111111111111111111111111000000;
		3373: Delta = 69'sb000000000000000001000000000000000000000000000000000000000000001000000;
		47616: Delta = 69'sb111111111111111111000000000000000000000000000000000000000000001000000;
		3245: Delta = 69'sb000000000000000000111111111111111111111111111111111111111111111000000;
		47488: Delta = 69'sb111111111111111110111111111111111111111111111111111111111111111000000;
		6682: Delta = 69'sb000000000000000010000000000000000000000000000000000000000000001000000;
		44307: Delta = 69'sb111111111111111110000000000000000000000000000000000000000000001000000;
		6554: Delta = 69'sb000000000000000001111111111111111111111111111111111111111111111000000;
		44179: Delta = 69'sb111111111111111101111111111111111111111111111111111111111111111000000;
		13300: Delta = 69'sb000000000000000100000000000000000000000000000000000000000000001000000;
		37689: Delta = 69'sb111111111111111100000000000000000000000000000000000000000000001000000;
		13172: Delta = 69'sb000000000000000011111111111111111111111111111111111111111111111000000;
		37561: Delta = 69'sb111111111111111011111111111111111111111111111111111111111111111000000;
		26536: Delta = 69'sb000000000000001000000000000000000000000000000000000000000000001000000;
		24453: Delta = 69'sb111111111111111000000000000000000000000000000000000000000000001000000;
		26408: Delta = 69'sb000000000000000111111111111111111111111111111111111111111111111000000;
		24325: Delta = 69'sb111111111111110111111111111111111111111111111111111111111111111000000;
		2147: Delta = 69'sb000000000000010000000000000000000000000000000000000000000000001000000;
		48842: Delta = 69'sb111111111111110000000000000000000000000000000000000000000000001000000;
		2019: Delta = 69'sb000000000000001111111111111111111111111111111111111111111111111000000;
		48714: Delta = 69'sb111111111111101111111111111111111111111111111111111111111111111000000;
		4230: Delta = 69'sb000000000000100000000000000000000000000000000000000000000000001000000;
		46759: Delta = 69'sb111111111111100000000000000000000000000000000000000000000000001000000;
		4102: Delta = 69'sb000000000000011111111111111111111111111111111111111111111111111000000;
		46631: Delta = 69'sb111111111111011111111111111111111111111111111111111111111111111000000;
		8396: Delta = 69'sb000000000001000000000000000000000000000000000000000000000000001000000;
		42593: Delta = 69'sb111111111111000000000000000000000000000000000000000000000000001000000;
		8268: Delta = 69'sb000000000000111111111111111111111111111111111111111111111111111000000;
		42465: Delta = 69'sb111111111110111111111111111111111111111111111111111111111111111000000;
		16728: Delta = 69'sb000000000010000000000000000000000000000000000000000000000000001000000;
		34261: Delta = 69'sb111111111110000000000000000000000000000000000000000000000000001000000;
		16600: Delta = 69'sb000000000001111111111111111111111111111111111111111111111111111000000;
		34133: Delta = 69'sb111111111101111111111111111111111111111111111111111111111111111000000;
		33392: Delta = 69'sb000000000100000000000000000000000000000000000000000000000000001000000;
		17597: Delta = 69'sb111111111100000000000000000000000000000000000000000000000000001000000;
		33264: Delta = 69'sb000000000011111111111111111111111111111111111111111111111111111000000;
		17469: Delta = 69'sb111111111011111111111111111111111111111111111111111111111111111000000;
		15859: Delta = 69'sb000000001000000000000000000000000000000000000000000000000000001000000;
		35130: Delta = 69'sb111111111000000000000000000000000000000000000000000000000000001000000;
		15731: Delta = 69'sb000000000111111111111111111111111111111111111111111111111111111000000;
		35002: Delta = 69'sb111111110111111111111111111111111111111111111111111111111111111000000;
		31654: Delta = 69'sb000000010000000000000000000000000000000000000000000000000000001000000;
		19335: Delta = 69'sb111111110000000000000000000000000000000000000000000000000000001000000;
		31526: Delta = 69'sb000000001111111111111111111111111111111111111111111111111111111000000;
		19207: Delta = 69'sb111111101111111111111111111111111111111111111111111111111111111000000;
		12383: Delta = 69'sb000000100000000000000000000000000000000000000000000000000000001000000;
		38606: Delta = 69'sb111111100000000000000000000000000000000000000000000000000000001000000;
		12255: Delta = 69'sb000000011111111111111111111111111111111111111111111111111111111000000;
		38478: Delta = 69'sb111111011111111111111111111111111111111111111111111111111111111000000;
		24702: Delta = 69'sb000001000000000000000000000000000000000000000000000000000000001000000;
		26287: Delta = 69'sb111111000000000000000000000000000000000000000000000000000000001000000;
		24574: Delta = 69'sb000000111111111111111111111111111111111111111111111111111111111000000;
		26159: Delta = 69'sb111110111111111111111111111111111111111111111111111111111111111000000;
		49340: Delta = 69'sb000010000000000000000000000000000000000000000000000000000000001000000;
		1649: Delta = 69'sb111110000000000000000000000000000000000000000000000000000000001000000;
		49212: Delta = 69'sb000001111111111111111111111111111111111111111111111111111111111000000;
		1521: Delta = 69'sb111101111111111111111111111111111111111111111111111111111111111000000;
		47755: Delta = 69'sb000100000000000000000000000000000000000000000000000000000000001000000;
		3234: Delta = 69'sb111100000000000000000000000000000000000000000000000000000000001000000;
		47627: Delta = 69'sb000011111111111111111111111111111111111111111111111111111111111000000;
		3106: Delta = 69'sb111011111111111111111111111111111111111111111111111111111111111000000;
		44585: Delta = 69'sb001000000000000000000000000000000000000000000000000000000000001000000;
		6404: Delta = 69'sb111000000000000000000000000000000000000000000000000000000000001000000;
		44457: Delta = 69'sb000111111111111111111111111111111111111111111111111111111111111000000;
		6276: Delta = 69'sb110111111111111111111111111111111111111111111111111111111111111000000;
		38245: Delta = 69'sb010000000000000000000000000000000000000000000000000000000000001000000;
		12744: Delta = 69'sb110000000000000000000000000000000000000000000000000000000000001000000;
		38117: Delta = 69'sb001111111111111111111111111111111111111111111111111111111111111000000;
		12616: Delta = 69'sb101111111111111111111111111111111111111111111111111111111111111000000;
		384: Delta = 69'sb000000000000000000000000000000000000000000000000000000000000110000000;
		50477: Delta = 69'sb111111111111111111111111111111111111111111111111111111111111010000000;
		640: Delta = 69'sb000000000000000000000000000000000000000000000000000000000001010000000;
		50221: Delta = 69'sb111111111111111111111111111111111111111111111111111111111110110000000;
		1152: Delta = 69'sb000000000000000000000000000000000000000000000000000000000010010000000;
		49965: Delta = 69'sb111111111111111111111111111111111111111111111111111111111110010000000;
		896: Delta = 69'sb000000000000000000000000000000000000000000000000000000000001110000000;
		49709: Delta = 69'sb111111111111111111111111111111111111111111111111111111111101110000000;
		2176: Delta = 69'sb000000000000000000000000000000000000000000000000000000000100010000000;
		48941: Delta = 69'sb111111111111111111111111111111111111111111111111111111111100010000000;
		1920: Delta = 69'sb000000000000000000000000000000000000000000000000000000000011110000000;
		48685: Delta = 69'sb111111111111111111111111111111111111111111111111111111111011110000000;
		4224: Delta = 69'sb000000000000000000000000000000000000000000000000000000001000010000000;
		46893: Delta = 69'sb111111111111111111111111111111111111111111111111111111111000010000000;
		3968: Delta = 69'sb000000000000000000000000000000000000000000000000000000000111110000000;
		46637: Delta = 69'sb111111111111111111111111111111111111111111111111111111110111110000000;
		8320: Delta = 69'sb000000000000000000000000000000000000000000000000000000010000010000000;
		42797: Delta = 69'sb111111111111111111111111111111111111111111111111111111110000010000000;
		8064: Delta = 69'sb000000000000000000000000000000000000000000000000000000001111110000000;
		42541: Delta = 69'sb111111111111111111111111111111111111111111111111111111101111110000000;
		16512: Delta = 69'sb000000000000000000000000000000000000000000000000000000100000010000000;
		34605: Delta = 69'sb111111111111111111111111111111111111111111111111111111100000010000000;
		16256: Delta = 69'sb000000000000000000000000000000000000000000000000000000011111110000000;
		34349: Delta = 69'sb111111111111111111111111111111111111111111111111111111011111110000000;
		32896: Delta = 69'sb000000000000000000000000000000000000000000000000000001000000010000000;
		18221: Delta = 69'sb111111111111111111111111111111111111111111111111111111000000010000000;
		32640: Delta = 69'sb000000000000000000000000000000000000000000000000000000111111110000000;
		17965: Delta = 69'sb111111111111111111111111111111111111111111111111111110111111110000000;
		14803: Delta = 69'sb000000000000000000000000000000000000000000000000000010000000010000000;
		36314: Delta = 69'sb111111111111111111111111111111111111111111111111111110000000010000000;
		14547: Delta = 69'sb000000000000000000000000000000000000000000000000000001111111110000000;
		36058: Delta = 69'sb111111111111111111111111111111111111111111111111111101111111110000000;
		29478: Delta = 69'sb000000000000000000000000000000000000000000000000000100000000010000000;
		21639: Delta = 69'sb111111111111111111111111111111111111111111111111111100000000010000000;
		29222: Delta = 69'sb000000000000000000000000000000000000000000000000000011111111110000000;
		21383: Delta = 69'sb111111111111111111111111111111111111111111111111111011111111110000000;
		7967: Delta = 69'sb000000000000000000000000000000000000000000000000001000000000010000000;
		43150: Delta = 69'sb111111111111111111111111111111111111111111111111111000000000010000000;
		7711: Delta = 69'sb000000000000000000000000000000000000000000000000000111111111110000000;
		42894: Delta = 69'sb111111111111111111111111111111111111111111111111110111111111110000000;
		15806: Delta = 69'sb000000000000000000000000000000000000000000000000010000000000010000000;
		35311: Delta = 69'sb111111111111111111111111111111111111111111111111110000000000010000000;
		15550: Delta = 69'sb000000000000000000000000000000000000000000000000001111111111110000000;
		35055: Delta = 69'sb111111111111111111111111111111111111111111111111101111111111110000000;
		31484: Delta = 69'sb000000000000000000000000000000000000000000000000100000000000010000000;
		19633: Delta = 69'sb111111111111111111111111111111111111111111111111100000000000010000000;
		31228: Delta = 69'sb000000000000000000000000000000000000000000000000011111111111110000000;
		19377: Delta = 69'sb111111111111111111111111111111111111111111111111011111111111110000000;
		11979: Delta = 69'sb000000000000000000000000000000000000000000000001000000000000010000000;
		39138: Delta = 69'sb111111111111111111111111111111111111111111111111000000000000010000000;
		11723: Delta = 69'sb000000000000000000000000000000000000000000000000111111111111110000000;
		38882: Delta = 69'sb111111111111111111111111111111111111111111111110111111111111110000000;
		23830: Delta = 69'sb000000000000000000000000000000000000000000000010000000000000010000000;
		27287: Delta = 69'sb111111111111111111111111111111111111111111111110000000000000010000000;
		23574: Delta = 69'sb000000000000000000000000000000000000000000000001111111111111110000000;
		27031: Delta = 69'sb111111111111111111111111111111111111111111111101111111111111110000000;
		47532: Delta = 69'sb000000000000000000000000000000000000000000000100000000000000010000000;
		3585: Delta = 69'sb111111111111111111111111111111111111111111111100000000000000010000000;
		47276: Delta = 69'sb000000000000000000000000000000000000000000000011111111111111110000000;
		3329: Delta = 69'sb111111111111111111111111111111111111111111111011111111111111110000000;
		44075: Delta = 69'sb000000000000000000000000000000000000000000001000000000000000010000000;
		7042: Delta = 69'sb111111111111111111111111111111111111111111111000000000000000010000000;
		43819: Delta = 69'sb000000000000000000000000000000000000000000000111111111111111110000000;
		6786: Delta = 69'sb111111111111111111111111111111111111111111110111111111111111110000000;
		37161: Delta = 69'sb000000000000000000000000000000000000000000010000000000000000010000000;
		13956: Delta = 69'sb111111111111111111111111111111111111111111110000000000000000010000000;
		36905: Delta = 69'sb000000000000000000000000000000000000000000001111111111111111110000000;
		13700: Delta = 69'sb111111111111111111111111111111111111111111101111111111111111110000000;
		23333: Delta = 69'sb000000000000000000000000000000000000000000100000000000000000010000000;
		27784: Delta = 69'sb111111111111111111111111111111111111111111100000000000000000010000000;
		23077: Delta = 69'sb000000000000000000000000000000000000000000011111111111111111110000000;
		27528: Delta = 69'sb111111111111111111111111111111111111111111011111111111111111110000000;
		46538: Delta = 69'sb000000000000000000000000000000000000000001000000000000000000010000000;
		4579: Delta = 69'sb111111111111111111111111111111111111111111000000000000000000010000000;
		46282: Delta = 69'sb000000000000000000000000000000000000000000111111111111111111110000000;
		4323: Delta = 69'sb111111111111111111111111111111111111111110111111111111111111110000000;
		42087: Delta = 69'sb000000000000000000000000000000000000000010000000000000000000010000000;
		9030: Delta = 69'sb111111111111111111111111111111111111111110000000000000000000010000000;
		41831: Delta = 69'sb000000000000000000000000000000000000000001111111111111111111110000000;
		8774: Delta = 69'sb111111111111111111111111111111111111111101111111111111111111110000000;
		33185: Delta = 69'sb000000000000000000000000000000000000000100000000000000000000010000000;
		17932: Delta = 69'sb111111111111111111111111111111111111111100000000000000000000010000000;
		32929: Delta = 69'sb000000000000000000000000000000000000000011111111111111111111110000000;
		17676: Delta = 69'sb111111111111111111111111111111111111111011111111111111111111110000000;
		15381: Delta = 69'sb000000000000000000000000000000000000001000000000000000000000010000000;
		35736: Delta = 69'sb111111111111111111111111111111111111111000000000000000000000010000000;
		15125: Delta = 69'sb000000000000000000000000000000000000000111111111111111111111110000000;
		35480: Delta = 69'sb111111111111111111111111111111111111110111111111111111111111110000000;
		30634: Delta = 69'sb000000000000000000000000000000000000010000000000000000000000010000000;
		20483: Delta = 69'sb111111111111111111111111111111111111110000000000000000000000010000000;
		30378: Delta = 69'sb000000000000000000000000000000000000001111111111111111111111110000000;
		20227: Delta = 69'sb111111111111111111111111111111111111101111111111111111111111110000000;
		10279: Delta = 69'sb000000000000000000000000000000000000100000000000000000000000010000000;
		40838: Delta = 69'sb111111111111111111111111111111111111100000000000000000000000010000000;
		10023: Delta = 69'sb000000000000000000000000000000000000011111111111111111111111110000000;
		40582: Delta = 69'sb111111111111111111111111111111111111011111111111111111111111110000000;
		20430: Delta = 69'sb000000000000000000000000000000000001000000000000000000000000010000000;
		30687: Delta = 69'sb111111111111111111111111111111111111000000000000000000000000010000000;
		20174: Delta = 69'sb000000000000000000000000000000000000111111111111111111111111110000000;
		30431: Delta = 69'sb111111111111111111111111111111111110111111111111111111111111110000000;
		40732: Delta = 69'sb000000000000000000000000000000000010000000000000000000000000010000000;
		10385: Delta = 69'sb111111111111111111111111111111111110000000000000000000000000010000000;
		40476: Delta = 69'sb000000000000000000000000000000000001111111111111111111111111110000000;
		10129: Delta = 69'sb111111111111111111111111111111111101111111111111111111111111110000000;
		30475: Delta = 69'sb000000000000000000000000000000000100000000000000000000000000010000000;
		20642: Delta = 69'sb111111111111111111111111111111111100000000000000000000000000010000000;
		30219: Delta = 69'sb000000000000000000000000000000000011111111111111111111111111110000000;
		20386: Delta = 69'sb111111111111111111111111111111111011111111111111111111111111110000000;
		9961: Delta = 69'sb000000000000000000000000000000001000000000000000000000000000010000000;
		41156: Delta = 69'sb111111111111111111111111111111111000000000000000000000000000010000000;
		9705: Delta = 69'sb000000000000000000000000000000000111111111111111111111111111110000000;
		40900: Delta = 69'sb111111111111111111111111111111110111111111111111111111111111110000000;
		19794: Delta = 69'sb000000000000000000000000000000010000000000000000000000000000010000000;
		31323: Delta = 69'sb111111111111111111111111111111110000000000000000000000000000010000000;
		19538: Delta = 69'sb000000000000000000000000000000001111111111111111111111111111110000000;
		31067: Delta = 69'sb111111111111111111111111111111101111111111111111111111111111110000000;
		39460: Delta = 69'sb000000000000000000000000000000100000000000000000000000000000010000000;
		11657: Delta = 69'sb111111111111111111111111111111100000000000000000000000000000010000000;
		39204: Delta = 69'sb000000000000000000000000000000011111111111111111111111111111110000000;
		11401: Delta = 69'sb111111111111111111111111111111011111111111111111111111111111110000000;
		27931: Delta = 69'sb000000000000000000000000000001000000000000000000000000000000010000000;
		23186: Delta = 69'sb111111111111111111111111111111000000000000000000000000000000010000000;
		27675: Delta = 69'sb000000000000000000000000000000111111111111111111111111111111110000000;
		22930: Delta = 69'sb111111111111111111111111111110111111111111111111111111111111110000000;
		4873: Delta = 69'sb000000000000000000000000000010000000000000000000000000000000010000000;
		46244: Delta = 69'sb111111111111111111111111111110000000000000000000000000000000010000000;
		4617: Delta = 69'sb000000000000000000000000000001111111111111111111111111111111110000000;
		45988: Delta = 69'sb111111111111111111111111111101111111111111111111111111111111110000000;
		9618: Delta = 69'sb000000000000000000000000000100000000000000000000000000000000010000000;
		41499: Delta = 69'sb111111111111111111111111111100000000000000000000000000000000010000000;
		9362: Delta = 69'sb000000000000000000000000000011111111111111111111111111111111110000000;
		41243: Delta = 69'sb111111111111111111111111111011111111111111111111111111111111110000000;
		19108: Delta = 69'sb000000000000000000000000001000000000000000000000000000000000010000000;
		32009: Delta = 69'sb111111111111111111111111111000000000000000000000000000000000010000000;
		18852: Delta = 69'sb000000000000000000000000000111111111111111111111111111111111110000000;
		31753: Delta = 69'sb111111111111111111111111110111111111111111111111111111111111110000000;
		38088: Delta = 69'sb000000000000000000000000010000000000000000000000000000000000010000000;
		13029: Delta = 69'sb111111111111111111111111110000000000000000000000000000000000010000000;
		37832: Delta = 69'sb000000000000000000000000001111111111111111111111111111111111110000000;
		12773: Delta = 69'sb111111111111111111111111101111111111111111111111111111111111110000000;
		25187: Delta = 69'sb000000000000000000000000100000000000000000000000000000000000010000000;
		25930: Delta = 69'sb111111111111111111111111100000000000000000000000000000000000010000000;
		24931: Delta = 69'sb000000000000000000000000011111111111111111111111111111111111110000000;
		25674: Delta = 69'sb111111111111111111111111011111111111111111111111111111111111110000000;
		50246: Delta = 69'sb000000000000000000000001000000000000000000000000000000000000010000000;
		871: Delta = 69'sb111111111111111111111111000000000000000000000000000000000000010000000;
		49990: Delta = 69'sb000000000000000000000000111111111111111111111111111111111111110000000;
		615: Delta = 69'sb111111111111111111111110111111111111111111111111111111111111110000000;
		49503: Delta = 69'sb000000000000000000000010000000000000000000000000000000000000010000000;
		1614: Delta = 69'sb111111111111111111111110000000000000000000000000000000000000010000000;
		49247: Delta = 69'sb000000000000000000000001111111111111111111111111111111111111110000000;
		1358: Delta = 69'sb111111111111111111111101111111111111111111111111111111111111110000000;
		48017: Delta = 69'sb000000000000000000000100000000000000000000000000000000000000010000000;
		3100: Delta = 69'sb111111111111111111111100000000000000000000000000000000000000010000000;
		47761: Delta = 69'sb000000000000000000000011111111111111111111111111111111111111110000000;
		2844: Delta = 69'sb111111111111111111111011111111111111111111111111111111111111110000000;
		45045: Delta = 69'sb000000000000000000001000000000000000000000000000000000000000010000000;
		6072: Delta = 69'sb111111111111111111111000000000000000000000000000000000000000010000000;
		44789: Delta = 69'sb000000000000000000000111111111111111111111111111111111111111110000000;
		5816: Delta = 69'sb111111111111111111110111111111111111111111111111111111111111110000000;
		39101: Delta = 69'sb000000000000000000010000000000000000000000000000000000000000010000000;
		12016: Delta = 69'sb111111111111111111110000000000000000000000000000000000000000010000000;
		38845: Delta = 69'sb000000000000000000001111111111111111111111111111111111111111110000000;
		11760: Delta = 69'sb111111111111111111101111111111111111111111111111111111111111110000000;
		27213: Delta = 69'sb000000000000000000100000000000000000000000000000000000000000010000000;
		23904: Delta = 69'sb111111111111111111100000000000000000000000000000000000000000010000000;
		26957: Delta = 69'sb000000000000000000011111111111111111111111111111111111111111110000000;
		23648: Delta = 69'sb111111111111111111011111111111111111111111111111111111111111110000000;
		3437: Delta = 69'sb000000000000000001000000000000000000000000000000000000000000010000000;
		47680: Delta = 69'sb111111111111111111000000000000000000000000000000000000000000010000000;
		3181: Delta = 69'sb000000000000000000111111111111111111111111111111111111111111110000000;
		47424: Delta = 69'sb111111111111111110111111111111111111111111111111111111111111110000000;
		6746: Delta = 69'sb000000000000000010000000000000000000000000000000000000000000010000000;
		44371: Delta = 69'sb111111111111111110000000000000000000000000000000000000000000010000000;
		6490: Delta = 69'sb000000000000000001111111111111111111111111111111111111111111110000000;
		44115: Delta = 69'sb111111111111111101111111111111111111111111111111111111111111110000000;
		13364: Delta = 69'sb000000000000000100000000000000000000000000000000000000000000010000000;
		37753: Delta = 69'sb111111111111111100000000000000000000000000000000000000000000010000000;
		13108: Delta = 69'sb000000000000000011111111111111111111111111111111111111111111110000000;
		37497: Delta = 69'sb111111111111111011111111111111111111111111111111111111111111110000000;
		26600: Delta = 69'sb000000000000001000000000000000000000000000000000000000000000010000000;
		24517: Delta = 69'sb111111111111111000000000000000000000000000000000000000000000010000000;
		26344: Delta = 69'sb000000000000000111111111111111111111111111111111111111111111110000000;
		24261: Delta = 69'sb111111111111110111111111111111111111111111111111111111111111110000000;
		2211: Delta = 69'sb000000000000010000000000000000000000000000000000000000000000010000000;
		48906: Delta = 69'sb111111111111110000000000000000000000000000000000000000000000010000000;
		1955: Delta = 69'sb000000000000001111111111111111111111111111111111111111111111110000000;
		48650: Delta = 69'sb111111111111101111111111111111111111111111111111111111111111110000000;
		4294: Delta = 69'sb000000000000100000000000000000000000000000000000000000000000010000000;
		46823: Delta = 69'sb111111111111100000000000000000000000000000000000000000000000010000000;
		4038: Delta = 69'sb000000000000011111111111111111111111111111111111111111111111110000000;
		46567: Delta = 69'sb111111111111011111111111111111111111111111111111111111111111110000000;
		8460: Delta = 69'sb000000000001000000000000000000000000000000000000000000000000010000000;
		42657: Delta = 69'sb111111111111000000000000000000000000000000000000000000000000010000000;
		8204: Delta = 69'sb000000000000111111111111111111111111111111111111111111111111110000000;
		42401: Delta = 69'sb111111111110111111111111111111111111111111111111111111111111110000000;
		16792: Delta = 69'sb000000000010000000000000000000000000000000000000000000000000010000000;
		34325: Delta = 69'sb111111111110000000000000000000000000000000000000000000000000010000000;
		16536: Delta = 69'sb000000000001111111111111111111111111111111111111111111111111110000000;
		34069: Delta = 69'sb111111111101111111111111111111111111111111111111111111111111110000000;
		33456: Delta = 69'sb000000000100000000000000000000000000000000000000000000000000010000000;
		17661: Delta = 69'sb111111111100000000000000000000000000000000000000000000000000010000000;
		33200: Delta = 69'sb000000000011111111111111111111111111111111111111111111111111110000000;
		17405: Delta = 69'sb111111111011111111111111111111111111111111111111111111111111110000000;
		15923: Delta = 69'sb000000001000000000000000000000000000000000000000000000000000010000000;
		35194: Delta = 69'sb111111111000000000000000000000000000000000000000000000000000010000000;
		15667: Delta = 69'sb000000000111111111111111111111111111111111111111111111111111110000000;
		34938: Delta = 69'sb111111110111111111111111111111111111111111111111111111111111110000000;
		31718: Delta = 69'sb000000010000000000000000000000000000000000000000000000000000010000000;
		19399: Delta = 69'sb111111110000000000000000000000000000000000000000000000000000010000000;
		31462: Delta = 69'sb000000001111111111111111111111111111111111111111111111111111110000000;
		19143: Delta = 69'sb111111101111111111111111111111111111111111111111111111111111110000000;
		12447: Delta = 69'sb000000100000000000000000000000000000000000000000000000000000010000000;
		38670: Delta = 69'sb111111100000000000000000000000000000000000000000000000000000010000000;
		12191: Delta = 69'sb000000011111111111111111111111111111111111111111111111111111110000000;
		38414: Delta = 69'sb111111011111111111111111111111111111111111111111111111111111110000000;
		24766: Delta = 69'sb000001000000000000000000000000000000000000000000000000000000010000000;
		26351: Delta = 69'sb111111000000000000000000000000000000000000000000000000000000010000000;
		24510: Delta = 69'sb000000111111111111111111111111111111111111111111111111111111110000000;
		26095: Delta = 69'sb111110111111111111111111111111111111111111111111111111111111110000000;
		49404: Delta = 69'sb000010000000000000000000000000000000000000000000000000000000010000000;
		1713: Delta = 69'sb111110000000000000000000000000000000000000000000000000000000010000000;
		49148: Delta = 69'sb000001111111111111111111111111111111111111111111111111111111110000000;
		1457: Delta = 69'sb111101111111111111111111111111111111111111111111111111111111110000000;
		47819: Delta = 69'sb000100000000000000000000000000000000000000000000000000000000010000000;
		3298: Delta = 69'sb111100000000000000000000000000000000000000000000000000000000010000000;
		47563: Delta = 69'sb000011111111111111111111111111111111111111111111111111111111110000000;
		3042: Delta = 69'sb111011111111111111111111111111111111111111111111111111111111110000000;
		44649: Delta = 69'sb001000000000000000000000000000000000000000000000000000000000010000000;
		6468: Delta = 69'sb111000000000000000000000000000000000000000000000000000000000010000000;
		44393: Delta = 69'sb000111111111111111111111111111111111111111111111111111111111110000000;
		6212: Delta = 69'sb110111111111111111111111111111111111111111111111111111111111110000000;
		38309: Delta = 69'sb010000000000000000000000000000000000000000000000000000000000010000000;
		12808: Delta = 69'sb110000000000000000000000000000000000000000000000000000000000010000000;
		38053: Delta = 69'sb001111111111111111111111111111111111111111111111111111111111110000000;
		12552: Delta = 69'sb101111111111111111111111111111111111111111111111111111111111110000000;
		768: Delta = 69'sb000000000000000000000000000000000000000000000000000000000001100000000;
		50093: Delta = 69'sb111111111111111111111111111111111111111111111111111111111110100000000;
		1280: Delta = 69'sb000000000000000000000000000000000000000000000000000000000010100000000;
		49581: Delta = 69'sb111111111111111111111111111111111111111111111111111111111101100000000;
		2304: Delta = 69'sb000000000000000000000000000000000000000000000000000000000100100000000;
		49069: Delta = 69'sb111111111111111111111111111111111111111111111111111111111100100000000;
		1792: Delta = 69'sb000000000000000000000000000000000000000000000000000000000011100000000;
		48557: Delta = 69'sb111111111111111111111111111111111111111111111111111111111011100000000;
		4352: Delta = 69'sb000000000000000000000000000000000000000000000000000000001000100000000;
		47021: Delta = 69'sb111111111111111111111111111111111111111111111111111111111000100000000;
		3840: Delta = 69'sb000000000000000000000000000000000000000000000000000000000111100000000;
		46509: Delta = 69'sb111111111111111111111111111111111111111111111111111111110111100000000;
		8448: Delta = 69'sb000000000000000000000000000000000000000000000000000000010000100000000;
		42925: Delta = 69'sb111111111111111111111111111111111111111111111111111111110000100000000;
		7936: Delta = 69'sb000000000000000000000000000000000000000000000000000000001111100000000;
		42413: Delta = 69'sb111111111111111111111111111111111111111111111111111111101111100000000;
		16640: Delta = 69'sb000000000000000000000000000000000000000000000000000000100000100000000;
		34733: Delta = 69'sb111111111111111111111111111111111111111111111111111111100000100000000;
		16128: Delta = 69'sb000000000000000000000000000000000000000000000000000000011111100000000;
		34221: Delta = 69'sb111111111111111111111111111111111111111111111111111111011111100000000;
		33024: Delta = 69'sb000000000000000000000000000000000000000000000000000001000000100000000;
		18349: Delta = 69'sb111111111111111111111111111111111111111111111111111111000000100000000;
		32512: Delta = 69'sb000000000000000000000000000000000000000000000000000000111111100000000;
		17837: Delta = 69'sb111111111111111111111111111111111111111111111111111110111111100000000;
		14931: Delta = 69'sb000000000000000000000000000000000000000000000000000010000000100000000;
		36442: Delta = 69'sb111111111111111111111111111111111111111111111111111110000000100000000;
		14419: Delta = 69'sb000000000000000000000000000000000000000000000000000001111111100000000;
		35930: Delta = 69'sb111111111111111111111111111111111111111111111111111101111111100000000;
		29606: Delta = 69'sb000000000000000000000000000000000000000000000000000100000000100000000;
		21767: Delta = 69'sb111111111111111111111111111111111111111111111111111100000000100000000;
		29094: Delta = 69'sb000000000000000000000000000000000000000000000000000011111111100000000;
		21255: Delta = 69'sb111111111111111111111111111111111111111111111111111011111111100000000;
		8095: Delta = 69'sb000000000000000000000000000000000000000000000000001000000000100000000;
		43278: Delta = 69'sb111111111111111111111111111111111111111111111111111000000000100000000;
		7583: Delta = 69'sb000000000000000000000000000000000000000000000000000111111111100000000;
		42766: Delta = 69'sb111111111111111111111111111111111111111111111111110111111111100000000;
		15934: Delta = 69'sb000000000000000000000000000000000000000000000000010000000000100000000;
		35439: Delta = 69'sb111111111111111111111111111111111111111111111111110000000000100000000;
		15422: Delta = 69'sb000000000000000000000000000000000000000000000000001111111111100000000;
		34927: Delta = 69'sb111111111111111111111111111111111111111111111111101111111111100000000;
		31612: Delta = 69'sb000000000000000000000000000000000000000000000000100000000000100000000;
		19761: Delta = 69'sb111111111111111111111111111111111111111111111111100000000000100000000;
		31100: Delta = 69'sb000000000000000000000000000000000000000000000000011111111111100000000;
		19249: Delta = 69'sb111111111111111111111111111111111111111111111111011111111111100000000;
		12107: Delta = 69'sb000000000000000000000000000000000000000000000001000000000000100000000;
		39266: Delta = 69'sb111111111111111111111111111111111111111111111111000000000000100000000;
		11595: Delta = 69'sb000000000000000000000000000000000000000000000000111111111111100000000;
		38754: Delta = 69'sb111111111111111111111111111111111111111111111110111111111111100000000;
		23958: Delta = 69'sb000000000000000000000000000000000000000000000010000000000000100000000;
		27415: Delta = 69'sb111111111111111111111111111111111111111111111110000000000000100000000;
		23446: Delta = 69'sb000000000000000000000000000000000000000000000001111111111111100000000;
		26903: Delta = 69'sb111111111111111111111111111111111111111111111101111111111111100000000;
		47660: Delta = 69'sb000000000000000000000000000000000000000000000100000000000000100000000;
		3713: Delta = 69'sb111111111111111111111111111111111111111111111100000000000000100000000;
		47148: Delta = 69'sb000000000000000000000000000000000000000000000011111111111111100000000;
		3201: Delta = 69'sb111111111111111111111111111111111111111111111011111111111111100000000;
		44203: Delta = 69'sb000000000000000000000000000000000000000000001000000000000000100000000;
		7170: Delta = 69'sb111111111111111111111111111111111111111111111000000000000000100000000;
		43691: Delta = 69'sb000000000000000000000000000000000000000000000111111111111111100000000;
		6658: Delta = 69'sb111111111111111111111111111111111111111111110111111111111111100000000;
		37289: Delta = 69'sb000000000000000000000000000000000000000000010000000000000000100000000;
		14084: Delta = 69'sb111111111111111111111111111111111111111111110000000000000000100000000;
		36777: Delta = 69'sb000000000000000000000000000000000000000000001111111111111111100000000;
		13572: Delta = 69'sb111111111111111111111111111111111111111111101111111111111111100000000;
		23461: Delta = 69'sb000000000000000000000000000000000000000000100000000000000000100000000;
		27912: Delta = 69'sb111111111111111111111111111111111111111111100000000000000000100000000;
		22949: Delta = 69'sb000000000000000000000000000000000000000000011111111111111111100000000;
		27400: Delta = 69'sb111111111111111111111111111111111111111111011111111111111111100000000;
		46666: Delta = 69'sb000000000000000000000000000000000000000001000000000000000000100000000;
		4707: Delta = 69'sb111111111111111111111111111111111111111111000000000000000000100000000;
		46154: Delta = 69'sb000000000000000000000000000000000000000000111111111111111111100000000;
		4195: Delta = 69'sb111111111111111111111111111111111111111110111111111111111111100000000;
		42215: Delta = 69'sb000000000000000000000000000000000000000010000000000000000000100000000;
		9158: Delta = 69'sb111111111111111111111111111111111111111110000000000000000000100000000;
		41703: Delta = 69'sb000000000000000000000000000000000000000001111111111111111111100000000;
		8646: Delta = 69'sb111111111111111111111111111111111111111101111111111111111111100000000;
		33313: Delta = 69'sb000000000000000000000000000000000000000100000000000000000000100000000;
		18060: Delta = 69'sb111111111111111111111111111111111111111100000000000000000000100000000;
		32801: Delta = 69'sb000000000000000000000000000000000000000011111111111111111111100000000;
		17548: Delta = 69'sb111111111111111111111111111111111111111011111111111111111111100000000;
		15509: Delta = 69'sb000000000000000000000000000000000000001000000000000000000000100000000;
		35864: Delta = 69'sb111111111111111111111111111111111111111000000000000000000000100000000;
		14997: Delta = 69'sb000000000000000000000000000000000000000111111111111111111111100000000;
		35352: Delta = 69'sb111111111111111111111111111111111111110111111111111111111111100000000;
		30762: Delta = 69'sb000000000000000000000000000000000000010000000000000000000000100000000;
		20611: Delta = 69'sb111111111111111111111111111111111111110000000000000000000000100000000;
		30250: Delta = 69'sb000000000000000000000000000000000000001111111111111111111111100000000;
		20099: Delta = 69'sb111111111111111111111111111111111111101111111111111111111111100000000;
		10407: Delta = 69'sb000000000000000000000000000000000000100000000000000000000000100000000;
		40966: Delta = 69'sb111111111111111111111111111111111111100000000000000000000000100000000;
		9895: Delta = 69'sb000000000000000000000000000000000000011111111111111111111111100000000;
		40454: Delta = 69'sb111111111111111111111111111111111111011111111111111111111111100000000;
		20558: Delta = 69'sb000000000000000000000000000000000001000000000000000000000000100000000;
		30815: Delta = 69'sb111111111111111111111111111111111111000000000000000000000000100000000;
		20046: Delta = 69'sb000000000000000000000000000000000000111111111111111111111111100000000;
		30303: Delta = 69'sb111111111111111111111111111111111110111111111111111111111111100000000;
		40860: Delta = 69'sb000000000000000000000000000000000010000000000000000000000000100000000;
		10513: Delta = 69'sb111111111111111111111111111111111110000000000000000000000000100000000;
		40348: Delta = 69'sb000000000000000000000000000000000001111111111111111111111111100000000;
		10001: Delta = 69'sb111111111111111111111111111111111101111111111111111111111111100000000;
		30603: Delta = 69'sb000000000000000000000000000000000100000000000000000000000000100000000;
		20770: Delta = 69'sb111111111111111111111111111111111100000000000000000000000000100000000;
		30091: Delta = 69'sb000000000000000000000000000000000011111111111111111111111111100000000;
		20258: Delta = 69'sb111111111111111111111111111111111011111111111111111111111111100000000;
		10089: Delta = 69'sb000000000000000000000000000000001000000000000000000000000000100000000;
		41284: Delta = 69'sb111111111111111111111111111111111000000000000000000000000000100000000;
		9577: Delta = 69'sb000000000000000000000000000000000111111111111111111111111111100000000;
		40772: Delta = 69'sb111111111111111111111111111111110111111111111111111111111111100000000;
		19922: Delta = 69'sb000000000000000000000000000000010000000000000000000000000000100000000;
		31451: Delta = 69'sb111111111111111111111111111111110000000000000000000000000000100000000;
		19410: Delta = 69'sb000000000000000000000000000000001111111111111111111111111111100000000;
		30939: Delta = 69'sb111111111111111111111111111111101111111111111111111111111111100000000;
		39588: Delta = 69'sb000000000000000000000000000000100000000000000000000000000000100000000;
		11785: Delta = 69'sb111111111111111111111111111111100000000000000000000000000000100000000;
		39076: Delta = 69'sb000000000000000000000000000000011111111111111111111111111111100000000;
		11273: Delta = 69'sb111111111111111111111111111111011111111111111111111111111111100000000;
		28059: Delta = 69'sb000000000000000000000000000001000000000000000000000000000000100000000;
		23314: Delta = 69'sb111111111111111111111111111111000000000000000000000000000000100000000;
		27547: Delta = 69'sb000000000000000000000000000000111111111111111111111111111111100000000;
		22802: Delta = 69'sb111111111111111111111111111110111111111111111111111111111111100000000;
		5001: Delta = 69'sb000000000000000000000000000010000000000000000000000000000000100000000;
		46372: Delta = 69'sb111111111111111111111111111110000000000000000000000000000000100000000;
		4489: Delta = 69'sb000000000000000000000000000001111111111111111111111111111111100000000;
		45860: Delta = 69'sb111111111111111111111111111101111111111111111111111111111111100000000;
		9746: Delta = 69'sb000000000000000000000000000100000000000000000000000000000000100000000;
		41627: Delta = 69'sb111111111111111111111111111100000000000000000000000000000000100000000;
		9234: Delta = 69'sb000000000000000000000000000011111111111111111111111111111111100000000;
		41115: Delta = 69'sb111111111111111111111111111011111111111111111111111111111111100000000;
		19236: Delta = 69'sb000000000000000000000000001000000000000000000000000000000000100000000;
		32137: Delta = 69'sb111111111111111111111111111000000000000000000000000000000000100000000;
		18724: Delta = 69'sb000000000000000000000000000111111111111111111111111111111111100000000;
		31625: Delta = 69'sb111111111111111111111111110111111111111111111111111111111111100000000;
		38216: Delta = 69'sb000000000000000000000000010000000000000000000000000000000000100000000;
		13157: Delta = 69'sb111111111111111111111111110000000000000000000000000000000000100000000;
		37704: Delta = 69'sb000000000000000000000000001111111111111111111111111111111111100000000;
		12645: Delta = 69'sb111111111111111111111111101111111111111111111111111111111111100000000;
		25315: Delta = 69'sb000000000000000000000000100000000000000000000000000000000000100000000;
		26058: Delta = 69'sb111111111111111111111111100000000000000000000000000000000000100000000;
		24803: Delta = 69'sb000000000000000000000000011111111111111111111111111111111111100000000;
		25546: Delta = 69'sb111111111111111111111111011111111111111111111111111111111111100000000;
		50374: Delta = 69'sb000000000000000000000001000000000000000000000000000000000000100000000;
		999: Delta = 69'sb111111111111111111111111000000000000000000000000000000000000100000000;
		49862: Delta = 69'sb000000000000000000000000111111111111111111111111111111111111100000000;
		487: Delta = 69'sb111111111111111111111110111111111111111111111111111111111111100000000;
		49631: Delta = 69'sb000000000000000000000010000000000000000000000000000000000000100000000;
		1742: Delta = 69'sb111111111111111111111110000000000000000000000000000000000000100000000;
		49119: Delta = 69'sb000000000000000000000001111111111111111111111111111111111111100000000;
		1230: Delta = 69'sb111111111111111111111101111111111111111111111111111111111111100000000;
		48145: Delta = 69'sb000000000000000000000100000000000000000000000000000000000000100000000;
		3228: Delta = 69'sb111111111111111111111100000000000000000000000000000000000000100000000;
		47633: Delta = 69'sb000000000000000000000011111111111111111111111111111111111111100000000;
		2716: Delta = 69'sb111111111111111111111011111111111111111111111111111111111111100000000;
		45173: Delta = 69'sb000000000000000000001000000000000000000000000000000000000000100000000;
		6200: Delta = 69'sb111111111111111111111000000000000000000000000000000000000000100000000;
		44661: Delta = 69'sb000000000000000000000111111111111111111111111111111111111111100000000;
		5688: Delta = 69'sb111111111111111111110111111111111111111111111111111111111111100000000;
		39229: Delta = 69'sb000000000000000000010000000000000000000000000000000000000000100000000;
		12144: Delta = 69'sb111111111111111111110000000000000000000000000000000000000000100000000;
		38717: Delta = 69'sb000000000000000000001111111111111111111111111111111111111111100000000;
		11632: Delta = 69'sb111111111111111111101111111111111111111111111111111111111111100000000;
		27341: Delta = 69'sb000000000000000000100000000000000000000000000000000000000000100000000;
		24032: Delta = 69'sb111111111111111111100000000000000000000000000000000000000000100000000;
		26829: Delta = 69'sb000000000000000000011111111111111111111111111111111111111111100000000;
		23520: Delta = 69'sb111111111111111111011111111111111111111111111111111111111111100000000;
		3565: Delta = 69'sb000000000000000001000000000000000000000000000000000000000000100000000;
		47808: Delta = 69'sb111111111111111111000000000000000000000000000000000000000000100000000;
		3053: Delta = 69'sb000000000000000000111111111111111111111111111111111111111111100000000;
		47296: Delta = 69'sb111111111111111110111111111111111111111111111111111111111111100000000;
		6874: Delta = 69'sb000000000000000010000000000000000000000000000000000000000000100000000;
		44499: Delta = 69'sb111111111111111110000000000000000000000000000000000000000000100000000;
		6362: Delta = 69'sb000000000000000001111111111111111111111111111111111111111111100000000;
		43987: Delta = 69'sb111111111111111101111111111111111111111111111111111111111111100000000;
		13492: Delta = 69'sb000000000000000100000000000000000000000000000000000000000000100000000;
		37881: Delta = 69'sb111111111111111100000000000000000000000000000000000000000000100000000;
		12980: Delta = 69'sb000000000000000011111111111111111111111111111111111111111111100000000;
		37369: Delta = 69'sb111111111111111011111111111111111111111111111111111111111111100000000;
		26728: Delta = 69'sb000000000000001000000000000000000000000000000000000000000000100000000;
		24645: Delta = 69'sb111111111111111000000000000000000000000000000000000000000000100000000;
		26216: Delta = 69'sb000000000000000111111111111111111111111111111111111111111111100000000;
		24133: Delta = 69'sb111111111111110111111111111111111111111111111111111111111111100000000;
		2339: Delta = 69'sb000000000000010000000000000000000000000000000000000000000000100000000;
		49034: Delta = 69'sb111111111111110000000000000000000000000000000000000000000000100000000;
		1827: Delta = 69'sb000000000000001111111111111111111111111111111111111111111111100000000;
		48522: Delta = 69'sb111111111111101111111111111111111111111111111111111111111111100000000;
		4422: Delta = 69'sb000000000000100000000000000000000000000000000000000000000000100000000;
		46951: Delta = 69'sb111111111111100000000000000000000000000000000000000000000000100000000;
		3910: Delta = 69'sb000000000000011111111111111111111111111111111111111111111111100000000;
		46439: Delta = 69'sb111111111111011111111111111111111111111111111111111111111111100000000;
		8588: Delta = 69'sb000000000001000000000000000000000000000000000000000000000000100000000;
		42785: Delta = 69'sb111111111111000000000000000000000000000000000000000000000000100000000;
		8076: Delta = 69'sb000000000000111111111111111111111111111111111111111111111111100000000;
		42273: Delta = 69'sb111111111110111111111111111111111111111111111111111111111111100000000;
		16920: Delta = 69'sb000000000010000000000000000000000000000000000000000000000000100000000;
		34453: Delta = 69'sb111111111110000000000000000000000000000000000000000000000000100000000;
		16408: Delta = 69'sb000000000001111111111111111111111111111111111111111111111111100000000;
		33941: Delta = 69'sb111111111101111111111111111111111111111111111111111111111111100000000;
		33584: Delta = 69'sb000000000100000000000000000000000000000000000000000000000000100000000;
		17789: Delta = 69'sb111111111100000000000000000000000000000000000000000000000000100000000;
		33072: Delta = 69'sb000000000011111111111111111111111111111111111111111111111111100000000;
		17277: Delta = 69'sb111111111011111111111111111111111111111111111111111111111111100000000;
		16051: Delta = 69'sb000000001000000000000000000000000000000000000000000000000000100000000;
		35322: Delta = 69'sb111111111000000000000000000000000000000000000000000000000000100000000;
		15539: Delta = 69'sb000000000111111111111111111111111111111111111111111111111111100000000;
		34810: Delta = 69'sb111111110111111111111111111111111111111111111111111111111111100000000;
		31846: Delta = 69'sb000000010000000000000000000000000000000000000000000000000000100000000;
		19527: Delta = 69'sb111111110000000000000000000000000000000000000000000000000000100000000;
		31334: Delta = 69'sb000000001111111111111111111111111111111111111111111111111111100000000;
		19015: Delta = 69'sb111111101111111111111111111111111111111111111111111111111111100000000;
		12575: Delta = 69'sb000000100000000000000000000000000000000000000000000000000000100000000;
		38798: Delta = 69'sb111111100000000000000000000000000000000000000000000000000000100000000;
		12063: Delta = 69'sb000000011111111111111111111111111111111111111111111111111111100000000;
		38286: Delta = 69'sb111111011111111111111111111111111111111111111111111111111111100000000;
		24894: Delta = 69'sb000001000000000000000000000000000000000000000000000000000000100000000;
		26479: Delta = 69'sb111111000000000000000000000000000000000000000000000000000000100000000;
		24382: Delta = 69'sb000000111111111111111111111111111111111111111111111111111111100000000;
		25967: Delta = 69'sb111110111111111111111111111111111111111111111111111111111111100000000;
		49532: Delta = 69'sb000010000000000000000000000000000000000000000000000000000000100000000;
		1841: Delta = 69'sb111110000000000000000000000000000000000000000000000000000000100000000;
		49020: Delta = 69'sb000001111111111111111111111111111111111111111111111111111111100000000;
		1329: Delta = 69'sb111101111111111111111111111111111111111111111111111111111111100000000;
		47947: Delta = 69'sb000100000000000000000000000000000000000000000000000000000000100000000;
		3426: Delta = 69'sb111100000000000000000000000000000000000000000000000000000000100000000;
		47435: Delta = 69'sb000011111111111111111111111111111111111111111111111111111111100000000;
		2914: Delta = 69'sb111011111111111111111111111111111111111111111111111111111111100000000;
		44777: Delta = 69'sb001000000000000000000000000000000000000000000000000000000000100000000;
		6596: Delta = 69'sb111000000000000000000000000000000000000000000000000000000000100000000;
		44265: Delta = 69'sb000111111111111111111111111111111111111111111111111111111111100000000;
		6084: Delta = 69'sb110111111111111111111111111111111111111111111111111111111111100000000;
		38437: Delta = 69'sb010000000000000000000000000000000000000000000000000000000000100000000;
		12936: Delta = 69'sb110000000000000000000000000000000000000000000000000000000000100000000;
		37925: Delta = 69'sb001111111111111111111111111111111111111111111111111111111111100000000;
		12424: Delta = 69'sb101111111111111111111111111111111111111111111111111111111111100000000;
		1536: Delta = 69'sb000000000000000000000000000000000000000000000000000000000011000000000;
		49325: Delta = 69'sb111111111111111111111111111111111111111111111111111111111101000000000;
		2560: Delta = 69'sb000000000000000000000000000000000000000000000000000000000101000000000;
		48301: Delta = 69'sb111111111111111111111111111111111111111111111111111111111011000000000;
		4608: Delta = 69'sb000000000000000000000000000000000000000000000000000000001001000000000;
		47277: Delta = 69'sb111111111111111111111111111111111111111111111111111111111001000000000;
		3584: Delta = 69'sb000000000000000000000000000000000000000000000000000000000111000000000;
		46253: Delta = 69'sb111111111111111111111111111111111111111111111111111111110111000000000;
		8704: Delta = 69'sb000000000000000000000000000000000000000000000000000000010001000000000;
		43181: Delta = 69'sb111111111111111111111111111111111111111111111111111111110001000000000;
		7680: Delta = 69'sb000000000000000000000000000000000000000000000000000000001111000000000;
		42157: Delta = 69'sb111111111111111111111111111111111111111111111111111111101111000000000;
		16896: Delta = 69'sb000000000000000000000000000000000000000000000000000000100001000000000;
		34989: Delta = 69'sb111111111111111111111111111111111111111111111111111111100001000000000;
		15872: Delta = 69'sb000000000000000000000000000000000000000000000000000000011111000000000;
		33965: Delta = 69'sb111111111111111111111111111111111111111111111111111111011111000000000;
		33280: Delta = 69'sb000000000000000000000000000000000000000000000000000001000001000000000;
		18605: Delta = 69'sb111111111111111111111111111111111111111111111111111111000001000000000;
		32256: Delta = 69'sb000000000000000000000000000000000000000000000000000000111111000000000;
		17581: Delta = 69'sb111111111111111111111111111111111111111111111111111110111111000000000;
		15187: Delta = 69'sb000000000000000000000000000000000000000000000000000010000001000000000;
		36698: Delta = 69'sb111111111111111111111111111111111111111111111111111110000001000000000;
		14163: Delta = 69'sb000000000000000000000000000000000000000000000000000001111111000000000;
		35674: Delta = 69'sb111111111111111111111111111111111111111111111111111101111111000000000;
		29862: Delta = 69'sb000000000000000000000000000000000000000000000000000100000001000000000;
		22023: Delta = 69'sb111111111111111111111111111111111111111111111111111100000001000000000;
		28838: Delta = 69'sb000000000000000000000000000000000000000000000000000011111111000000000;
		20999: Delta = 69'sb111111111111111111111111111111111111111111111111111011111111000000000;
		8351: Delta = 69'sb000000000000000000000000000000000000000000000000001000000001000000000;
		43534: Delta = 69'sb111111111111111111111111111111111111111111111111111000000001000000000;
		7327: Delta = 69'sb000000000000000000000000000000000000000000000000000111111111000000000;
		42510: Delta = 69'sb111111111111111111111111111111111111111111111111110111111111000000000;
		16190: Delta = 69'sb000000000000000000000000000000000000000000000000010000000001000000000;
		35695: Delta = 69'sb111111111111111111111111111111111111111111111111110000000001000000000;
		15166: Delta = 69'sb000000000000000000000000000000000000000000000000001111111111000000000;
		34671: Delta = 69'sb111111111111111111111111111111111111111111111111101111111111000000000;
		31868: Delta = 69'sb000000000000000000000000000000000000000000000000100000000001000000000;
		20017: Delta = 69'sb111111111111111111111111111111111111111111111111100000000001000000000;
		30844: Delta = 69'sb000000000000000000000000000000000000000000000000011111111111000000000;
		18993: Delta = 69'sb111111111111111111111111111111111111111111111111011111111111000000000;
		12363: Delta = 69'sb000000000000000000000000000000000000000000000001000000000001000000000;
		39522: Delta = 69'sb111111111111111111111111111111111111111111111111000000000001000000000;
		11339: Delta = 69'sb000000000000000000000000000000000000000000000000111111111111000000000;
		38498: Delta = 69'sb111111111111111111111111111111111111111111111110111111111111000000000;
		24214: Delta = 69'sb000000000000000000000000000000000000000000000010000000000001000000000;
		27671: Delta = 69'sb111111111111111111111111111111111111111111111110000000000001000000000;
		23190: Delta = 69'sb000000000000000000000000000000000000000000000001111111111111000000000;
		26647: Delta = 69'sb111111111111111111111111111111111111111111111101111111111111000000000;
		47916: Delta = 69'sb000000000000000000000000000000000000000000000100000000000001000000000;
		3969: Delta = 69'sb111111111111111111111111111111111111111111111100000000000001000000000;
		46892: Delta = 69'sb000000000000000000000000000000000000000000000011111111111111000000000;
		2945: Delta = 69'sb111111111111111111111111111111111111111111111011111111111111000000000;
		44459: Delta = 69'sb000000000000000000000000000000000000000000001000000000000001000000000;
		7426: Delta = 69'sb111111111111111111111111111111111111111111111000000000000001000000000;
		43435: Delta = 69'sb000000000000000000000000000000000000000000000111111111111111000000000;
		6402: Delta = 69'sb111111111111111111111111111111111111111111110111111111111111000000000;
		37545: Delta = 69'sb000000000000000000000000000000000000000000010000000000000001000000000;
		14340: Delta = 69'sb111111111111111111111111111111111111111111110000000000000001000000000;
		36521: Delta = 69'sb000000000000000000000000000000000000000000001111111111111111000000000;
		13316: Delta = 69'sb111111111111111111111111111111111111111111101111111111111111000000000;
		23717: Delta = 69'sb000000000000000000000000000000000000000000100000000000000001000000000;
		28168: Delta = 69'sb111111111111111111111111111111111111111111100000000000000001000000000;
		22693: Delta = 69'sb000000000000000000000000000000000000000000011111111111111111000000000;
		27144: Delta = 69'sb111111111111111111111111111111111111111111011111111111111111000000000;
		46922: Delta = 69'sb000000000000000000000000000000000000000001000000000000000001000000000;
		4963: Delta = 69'sb111111111111111111111111111111111111111111000000000000000001000000000;
		45898: Delta = 69'sb000000000000000000000000000000000000000000111111111111111111000000000;
		3939: Delta = 69'sb111111111111111111111111111111111111111110111111111111111111000000000;
		42471: Delta = 69'sb000000000000000000000000000000000000000010000000000000000001000000000;
		9414: Delta = 69'sb111111111111111111111111111111111111111110000000000000000001000000000;
		41447: Delta = 69'sb000000000000000000000000000000000000000001111111111111111111000000000;
		8390: Delta = 69'sb111111111111111111111111111111111111111101111111111111111111000000000;
		33569: Delta = 69'sb000000000000000000000000000000000000000100000000000000000001000000000;
		18316: Delta = 69'sb111111111111111111111111111111111111111100000000000000000001000000000;
		32545: Delta = 69'sb000000000000000000000000000000000000000011111111111111111111000000000;
		17292: Delta = 69'sb111111111111111111111111111111111111111011111111111111111111000000000;
		15765: Delta = 69'sb000000000000000000000000000000000000001000000000000000000001000000000;
		36120: Delta = 69'sb111111111111111111111111111111111111111000000000000000000001000000000;
		14741: Delta = 69'sb000000000000000000000000000000000000000111111111111111111111000000000;
		35096: Delta = 69'sb111111111111111111111111111111111111110111111111111111111111000000000;
		31018: Delta = 69'sb000000000000000000000000000000000000010000000000000000000001000000000;
		20867: Delta = 69'sb111111111111111111111111111111111111110000000000000000000001000000000;
		29994: Delta = 69'sb000000000000000000000000000000000000001111111111111111111111000000000;
		19843: Delta = 69'sb111111111111111111111111111111111111101111111111111111111111000000000;
		10663: Delta = 69'sb000000000000000000000000000000000000100000000000000000000001000000000;
		41222: Delta = 69'sb111111111111111111111111111111111111100000000000000000000001000000000;
		9639: Delta = 69'sb000000000000000000000000000000000000011111111111111111111111000000000;
		40198: Delta = 69'sb111111111111111111111111111111111111011111111111111111111111000000000;
		20814: Delta = 69'sb000000000000000000000000000000000001000000000000000000000001000000000;
		31071: Delta = 69'sb111111111111111111111111111111111111000000000000000000000001000000000;
		19790: Delta = 69'sb000000000000000000000000000000000000111111111111111111111111000000000;
		30047: Delta = 69'sb111111111111111111111111111111111110111111111111111111111111000000000;
		41116: Delta = 69'sb000000000000000000000000000000000010000000000000000000000001000000000;
		10769: Delta = 69'sb111111111111111111111111111111111110000000000000000000000001000000000;
		40092: Delta = 69'sb000000000000000000000000000000000001111111111111111111111111000000000;
		9745: Delta = 69'sb111111111111111111111111111111111101111111111111111111111111000000000;
		30859: Delta = 69'sb000000000000000000000000000000000100000000000000000000000001000000000;
		21026: Delta = 69'sb111111111111111111111111111111111100000000000000000000000001000000000;
		29835: Delta = 69'sb000000000000000000000000000000000011111111111111111111111111000000000;
		20002: Delta = 69'sb111111111111111111111111111111111011111111111111111111111111000000000;
		10345: Delta = 69'sb000000000000000000000000000000001000000000000000000000000001000000000;
		41540: Delta = 69'sb111111111111111111111111111111111000000000000000000000000001000000000;
		9321: Delta = 69'sb000000000000000000000000000000000111111111111111111111111111000000000;
		40516: Delta = 69'sb111111111111111111111111111111110111111111111111111111111111000000000;
		20178: Delta = 69'sb000000000000000000000000000000010000000000000000000000000001000000000;
		31707: Delta = 69'sb111111111111111111111111111111110000000000000000000000000001000000000;
		19154: Delta = 69'sb000000000000000000000000000000001111111111111111111111111111000000000;
		30683: Delta = 69'sb111111111111111111111111111111101111111111111111111111111111000000000;
		39844: Delta = 69'sb000000000000000000000000000000100000000000000000000000000001000000000;
		12041: Delta = 69'sb111111111111111111111111111111100000000000000000000000000001000000000;
		38820: Delta = 69'sb000000000000000000000000000000011111111111111111111111111111000000000;
		11017: Delta = 69'sb111111111111111111111111111111011111111111111111111111111111000000000;
		28315: Delta = 69'sb000000000000000000000000000001000000000000000000000000000001000000000;
		23570: Delta = 69'sb111111111111111111111111111111000000000000000000000000000001000000000;
		27291: Delta = 69'sb000000000000000000000000000000111111111111111111111111111111000000000;
		22546: Delta = 69'sb111111111111111111111111111110111111111111111111111111111111000000000;
		5257: Delta = 69'sb000000000000000000000000000010000000000000000000000000000001000000000;
		46628: Delta = 69'sb111111111111111111111111111110000000000000000000000000000001000000000;
		4233: Delta = 69'sb000000000000000000000000000001111111111111111111111111111111000000000;
		45604: Delta = 69'sb111111111111111111111111111101111111111111111111111111111111000000000;
		10002: Delta = 69'sb000000000000000000000000000100000000000000000000000000000001000000000;
		41883: Delta = 69'sb111111111111111111111111111100000000000000000000000000000001000000000;
		8978: Delta = 69'sb000000000000000000000000000011111111111111111111111111111111000000000;
		40859: Delta = 69'sb111111111111111111111111111011111111111111111111111111111111000000000;
		19492: Delta = 69'sb000000000000000000000000001000000000000000000000000000000001000000000;
		32393: Delta = 69'sb111111111111111111111111111000000000000000000000000000000001000000000;
		18468: Delta = 69'sb000000000000000000000000000111111111111111111111111111111111000000000;
		31369: Delta = 69'sb111111111111111111111111110111111111111111111111111111111111000000000;
		38472: Delta = 69'sb000000000000000000000000010000000000000000000000000000000001000000000;
		13413: Delta = 69'sb111111111111111111111111110000000000000000000000000000000001000000000;
		37448: Delta = 69'sb000000000000000000000000001111111111111111111111111111111111000000000;
		12389: Delta = 69'sb111111111111111111111111101111111111111111111111111111111111000000000;
		25571: Delta = 69'sb000000000000000000000000100000000000000000000000000000000001000000000;
		26314: Delta = 69'sb111111111111111111111111100000000000000000000000000000000001000000000;
		24547: Delta = 69'sb000000000000000000000000011111111111111111111111111111111111000000000;
		25290: Delta = 69'sb111111111111111111111111011111111111111111111111111111111111000000000;
		50630: Delta = 69'sb000000000000000000000001000000000000000000000000000000000001000000000;
		1255: Delta = 69'sb111111111111111111111111000000000000000000000000000000000001000000000;
		49606: Delta = 69'sb000000000000000000000000111111111111111111111111111111111111000000000;
		231: Delta = 69'sb111111111111111111111110111111111111111111111111111111111111000000000;
		49887: Delta = 69'sb000000000000000000000010000000000000000000000000000000000001000000000;
		1998: Delta = 69'sb111111111111111111111110000000000000000000000000000000000001000000000;
		48863: Delta = 69'sb000000000000000000000001111111111111111111111111111111111111000000000;
		974: Delta = 69'sb111111111111111111111101111111111111111111111111111111111111000000000;
		48401: Delta = 69'sb000000000000000000000100000000000000000000000000000000000001000000000;
		3484: Delta = 69'sb111111111111111111111100000000000000000000000000000000000001000000000;
		47377: Delta = 69'sb000000000000000000000011111111111111111111111111111111111111000000000;
		2460: Delta = 69'sb111111111111111111111011111111111111111111111111111111111111000000000;
		45429: Delta = 69'sb000000000000000000001000000000000000000000000000000000000001000000000;
		6456: Delta = 69'sb111111111111111111111000000000000000000000000000000000000001000000000;
		44405: Delta = 69'sb000000000000000000000111111111111111111111111111111111111111000000000;
		5432: Delta = 69'sb111111111111111111110111111111111111111111111111111111111111000000000;
		39485: Delta = 69'sb000000000000000000010000000000000000000000000000000000000001000000000;
		12400: Delta = 69'sb111111111111111111110000000000000000000000000000000000000001000000000;
		38461: Delta = 69'sb000000000000000000001111111111111111111111111111111111111111000000000;
		11376: Delta = 69'sb111111111111111111101111111111111111111111111111111111111111000000000;
		27597: Delta = 69'sb000000000000000000100000000000000000000000000000000000000001000000000;
		24288: Delta = 69'sb111111111111111111100000000000000000000000000000000000000001000000000;
		26573: Delta = 69'sb000000000000000000011111111111111111111111111111111111111111000000000;
		23264: Delta = 69'sb111111111111111111011111111111111111111111111111111111111111000000000;
		3821: Delta = 69'sb000000000000000001000000000000000000000000000000000000000001000000000;
		48064: Delta = 69'sb111111111111111111000000000000000000000000000000000000000001000000000;
		2797: Delta = 69'sb000000000000000000111111111111111111111111111111111111111111000000000;
		47040: Delta = 69'sb111111111111111110111111111111111111111111111111111111111111000000000;
		7130: Delta = 69'sb000000000000000010000000000000000000000000000000000000000001000000000;
		44755: Delta = 69'sb111111111111111110000000000000000000000000000000000000000001000000000;
		6106: Delta = 69'sb000000000000000001111111111111111111111111111111111111111111000000000;
		43731: Delta = 69'sb111111111111111101111111111111111111111111111111111111111111000000000;
		13748: Delta = 69'sb000000000000000100000000000000000000000000000000000000000001000000000;
		38137: Delta = 69'sb111111111111111100000000000000000000000000000000000000000001000000000;
		12724: Delta = 69'sb000000000000000011111111111111111111111111111111111111111111000000000;
		37113: Delta = 69'sb111111111111111011111111111111111111111111111111111111111111000000000;
		26984: Delta = 69'sb000000000000001000000000000000000000000000000000000000000001000000000;
		24901: Delta = 69'sb111111111111111000000000000000000000000000000000000000000001000000000;
		25960: Delta = 69'sb000000000000000111111111111111111111111111111111111111111111000000000;
		23877: Delta = 69'sb111111111111110111111111111111111111111111111111111111111111000000000;
		2595: Delta = 69'sb000000000000010000000000000000000000000000000000000000000001000000000;
		49290: Delta = 69'sb111111111111110000000000000000000000000000000000000000000001000000000;
		1571: Delta = 69'sb000000000000001111111111111111111111111111111111111111111111000000000;
		48266: Delta = 69'sb111111111111101111111111111111111111111111111111111111111111000000000;
		4678: Delta = 69'sb000000000000100000000000000000000000000000000000000000000001000000000;
		47207: Delta = 69'sb111111111111100000000000000000000000000000000000000000000001000000000;
		3654: Delta = 69'sb000000000000011111111111111111111111111111111111111111111111000000000;
		46183: Delta = 69'sb111111111111011111111111111111111111111111111111111111111111000000000;
		8844: Delta = 69'sb000000000001000000000000000000000000000000000000000000000001000000000;
		43041: Delta = 69'sb111111111111000000000000000000000000000000000000000000000001000000000;
		7820: Delta = 69'sb000000000000111111111111111111111111111111111111111111111111000000000;
		42017: Delta = 69'sb111111111110111111111111111111111111111111111111111111111111000000000;
		17176: Delta = 69'sb000000000010000000000000000000000000000000000000000000000001000000000;
		34709: Delta = 69'sb111111111110000000000000000000000000000000000000000000000001000000000;
		16152: Delta = 69'sb000000000001111111111111111111111111111111111111111111111111000000000;
		33685: Delta = 69'sb111111111101111111111111111111111111111111111111111111111111000000000;
		33840: Delta = 69'sb000000000100000000000000000000000000000000000000000000000001000000000;
		18045: Delta = 69'sb111111111100000000000000000000000000000000000000000000000001000000000;
		32816: Delta = 69'sb000000000011111111111111111111111111111111111111111111111111000000000;
		17021: Delta = 69'sb111111111011111111111111111111111111111111111111111111111111000000000;
		16307: Delta = 69'sb000000001000000000000000000000000000000000000000000000000001000000000;
		35578: Delta = 69'sb111111111000000000000000000000000000000000000000000000000001000000000;
		15283: Delta = 69'sb000000000111111111111111111111111111111111111111111111111111000000000;
		34554: Delta = 69'sb111111110111111111111111111111111111111111111111111111111111000000000;
		32102: Delta = 69'sb000000010000000000000000000000000000000000000000000000000001000000000;
		19783: Delta = 69'sb111111110000000000000000000000000000000000000000000000000001000000000;
		31078: Delta = 69'sb000000001111111111111111111111111111111111111111111111111111000000000;
		18759: Delta = 69'sb111111101111111111111111111111111111111111111111111111111111000000000;
		12831: Delta = 69'sb000000100000000000000000000000000000000000000000000000000001000000000;
		39054: Delta = 69'sb111111100000000000000000000000000000000000000000000000000001000000000;
		11807: Delta = 69'sb000000011111111111111111111111111111111111111111111111111111000000000;
		38030: Delta = 69'sb111111011111111111111111111111111111111111111111111111111111000000000;
		25150: Delta = 69'sb000001000000000000000000000000000000000000000000000000000001000000000;
		26735: Delta = 69'sb111111000000000000000000000000000000000000000000000000000001000000000;
		24126: Delta = 69'sb000000111111111111111111111111111111111111111111111111111111000000000;
		25711: Delta = 69'sb111110111111111111111111111111111111111111111111111111111111000000000;
		49788: Delta = 69'sb000010000000000000000000000000000000000000000000000000000001000000000;
		2097: Delta = 69'sb111110000000000000000000000000000000000000000000000000000001000000000;
		48764: Delta = 69'sb000001111111111111111111111111111111111111111111111111111111000000000;
		1073: Delta = 69'sb111101111111111111111111111111111111111111111111111111111111000000000;
		48203: Delta = 69'sb000100000000000000000000000000000000000000000000000000000001000000000;
		3682: Delta = 69'sb111100000000000000000000000000000000000000000000000000000001000000000;
		47179: Delta = 69'sb000011111111111111111111111111111111111111111111111111111111000000000;
		2658: Delta = 69'sb111011111111111111111111111111111111111111111111111111111111000000000;
		45033: Delta = 69'sb001000000000000000000000000000000000000000000000000000000001000000000;
		6852: Delta = 69'sb111000000000000000000000000000000000000000000000000000000001000000000;
		44009: Delta = 69'sb000111111111111111111111111111111111111111111111111111111111000000000;
		5828: Delta = 69'sb110111111111111111111111111111111111111111111111111111111111000000000;
		38693: Delta = 69'sb010000000000000000000000000000000000000000000000000000000001000000000;
		13192: Delta = 69'sb110000000000000000000000000000000000000000000000000000000001000000000;
		37669: Delta = 69'sb001111111111111111111111111111111111111111111111111111111111000000000;
		12168: Delta = 69'sb101111111111111111111111111111111111111111111111111111111111000000000;
		3072: Delta = 69'sb000000000000000000000000000000000000000000000000000000000110000000000;
		47789: Delta = 69'sb111111111111111111111111111111111111111111111111111111111010000000000;
		5120: Delta = 69'sb000000000000000000000000000000000000000000000000000000001010000000000;
		45741: Delta = 69'sb111111111111111111111111111111111111111111111111111111110110000000000;
		9216: Delta = 69'sb000000000000000000000000000000000000000000000000000000010010000000000;
		43693: Delta = 69'sb111111111111111111111111111111111111111111111111111111110010000000000;
		7168: Delta = 69'sb000000000000000000000000000000000000000000000000000000001110000000000;
		41645: Delta = 69'sb111111111111111111111111111111111111111111111111111111101110000000000;
		17408: Delta = 69'sb000000000000000000000000000000000000000000000000000000100010000000000;
		35501: Delta = 69'sb111111111111111111111111111111111111111111111111111111100010000000000;
		15360: Delta = 69'sb000000000000000000000000000000000000000000000000000000011110000000000;
		33453: Delta = 69'sb111111111111111111111111111111111111111111111111111111011110000000000;
		33792: Delta = 69'sb000000000000000000000000000000000000000000000000000001000010000000000;
		19117: Delta = 69'sb111111111111111111111111111111111111111111111111111111000010000000000;
		31744: Delta = 69'sb000000000000000000000000000000000000000000000000000000111110000000000;
		17069: Delta = 69'sb111111111111111111111111111111111111111111111111111110111110000000000;
		15699: Delta = 69'sb000000000000000000000000000000000000000000000000000010000010000000000;
		37210: Delta = 69'sb111111111111111111111111111111111111111111111111111110000010000000000;
		13651: Delta = 69'sb000000000000000000000000000000000000000000000000000001111110000000000;
		35162: Delta = 69'sb111111111111111111111111111111111111111111111111111101111110000000000;
		30374: Delta = 69'sb000000000000000000000000000000000000000000000000000100000010000000000;
		22535: Delta = 69'sb111111111111111111111111111111111111111111111111111100000010000000000;
		28326: Delta = 69'sb000000000000000000000000000000000000000000000000000011111110000000000;
		20487: Delta = 69'sb111111111111111111111111111111111111111111111111111011111110000000000;
		8863: Delta = 69'sb000000000000000000000000000000000000000000000000001000000010000000000;
		44046: Delta = 69'sb111111111111111111111111111111111111111111111111111000000010000000000;
		6815: Delta = 69'sb000000000000000000000000000000000000000000000000000111111110000000000;
		41998: Delta = 69'sb111111111111111111111111111111111111111111111111110111111110000000000;
		16702: Delta = 69'sb000000000000000000000000000000000000000000000000010000000010000000000;
		36207: Delta = 69'sb111111111111111111111111111111111111111111111111110000000010000000000;
		14654: Delta = 69'sb000000000000000000000000000000000000000000000000001111111110000000000;
		34159: Delta = 69'sb111111111111111111111111111111111111111111111111101111111110000000000;
		32380: Delta = 69'sb000000000000000000000000000000000000000000000000100000000010000000000;
		20529: Delta = 69'sb111111111111111111111111111111111111111111111111100000000010000000000;
		30332: Delta = 69'sb000000000000000000000000000000000000000000000000011111111110000000000;
		18481: Delta = 69'sb111111111111111111111111111111111111111111111111011111111110000000000;
		12875: Delta = 69'sb000000000000000000000000000000000000000000000001000000000010000000000;
		40034: Delta = 69'sb111111111111111111111111111111111111111111111111000000000010000000000;
		10827: Delta = 69'sb000000000000000000000000000000000000000000000000111111111110000000000;
		37986: Delta = 69'sb111111111111111111111111111111111111111111111110111111111110000000000;
		24726: Delta = 69'sb000000000000000000000000000000000000000000000010000000000010000000000;
		28183: Delta = 69'sb111111111111111111111111111111111111111111111110000000000010000000000;
		22678: Delta = 69'sb000000000000000000000000000000000000000000000001111111111110000000000;
		26135: Delta = 69'sb111111111111111111111111111111111111111111111101111111111110000000000;
		48428: Delta = 69'sb000000000000000000000000000000000000000000000100000000000010000000000;
		4481: Delta = 69'sb111111111111111111111111111111111111111111111100000000000010000000000;
		46380: Delta = 69'sb000000000000000000000000000000000000000000000011111111111110000000000;
		2433: Delta = 69'sb111111111111111111111111111111111111111111111011111111111110000000000;
		44971: Delta = 69'sb000000000000000000000000000000000000000000001000000000000010000000000;
		7938: Delta = 69'sb111111111111111111111111111111111111111111111000000000000010000000000;
		42923: Delta = 69'sb000000000000000000000000000000000000000000000111111111111110000000000;
		5890: Delta = 69'sb111111111111111111111111111111111111111111110111111111111110000000000;
		38057: Delta = 69'sb000000000000000000000000000000000000000000010000000000000010000000000;
		14852: Delta = 69'sb111111111111111111111111111111111111111111110000000000000010000000000;
		36009: Delta = 69'sb000000000000000000000000000000000000000000001111111111111110000000000;
		12804: Delta = 69'sb111111111111111111111111111111111111111111101111111111111110000000000;
		24229: Delta = 69'sb000000000000000000000000000000000000000000100000000000000010000000000;
		28680: Delta = 69'sb111111111111111111111111111111111111111111100000000000000010000000000;
		22181: Delta = 69'sb000000000000000000000000000000000000000000011111111111111110000000000;
		26632: Delta = 69'sb111111111111111111111111111111111111111111011111111111111110000000000;
		47434: Delta = 69'sb000000000000000000000000000000000000000001000000000000000010000000000;
		5475: Delta = 69'sb111111111111111111111111111111111111111111000000000000000010000000000;
		45386: Delta = 69'sb000000000000000000000000000000000000000000111111111111111110000000000;
		3427: Delta = 69'sb111111111111111111111111111111111111111110111111111111111110000000000;
		42983: Delta = 69'sb000000000000000000000000000000000000000010000000000000000010000000000;
		9926: Delta = 69'sb111111111111111111111111111111111111111110000000000000000010000000000;
		40935: Delta = 69'sb000000000000000000000000000000000000000001111111111111111110000000000;
		7878: Delta = 69'sb111111111111111111111111111111111111111101111111111111111110000000000;
		34081: Delta = 69'sb000000000000000000000000000000000000000100000000000000000010000000000;
		18828: Delta = 69'sb111111111111111111111111111111111111111100000000000000000010000000000;
		32033: Delta = 69'sb000000000000000000000000000000000000000011111111111111111110000000000;
		16780: Delta = 69'sb111111111111111111111111111111111111111011111111111111111110000000000;
		16277: Delta = 69'sb000000000000000000000000000000000000001000000000000000000010000000000;
		36632: Delta = 69'sb111111111111111111111111111111111111111000000000000000000010000000000;
		14229: Delta = 69'sb000000000000000000000000000000000000000111111111111111111110000000000;
		34584: Delta = 69'sb111111111111111111111111111111111111110111111111111111111110000000000;
		31530: Delta = 69'sb000000000000000000000000000000000000010000000000000000000010000000000;
		21379: Delta = 69'sb111111111111111111111111111111111111110000000000000000000010000000000;
		29482: Delta = 69'sb000000000000000000000000000000000000001111111111111111111110000000000;
		19331: Delta = 69'sb111111111111111111111111111111111111101111111111111111111110000000000;
		11175: Delta = 69'sb000000000000000000000000000000000000100000000000000000000010000000000;
		41734: Delta = 69'sb111111111111111111111111111111111111100000000000000000000010000000000;
		9127: Delta = 69'sb000000000000000000000000000000000000011111111111111111111110000000000;
		39686: Delta = 69'sb111111111111111111111111111111111111011111111111111111111110000000000;
		21326: Delta = 69'sb000000000000000000000000000000000001000000000000000000000010000000000;
		31583: Delta = 69'sb111111111111111111111111111111111111000000000000000000000010000000000;
		19278: Delta = 69'sb000000000000000000000000000000000000111111111111111111111110000000000;
		29535: Delta = 69'sb111111111111111111111111111111111110111111111111111111111110000000000;
		41628: Delta = 69'sb000000000000000000000000000000000010000000000000000000000010000000000;
		11281: Delta = 69'sb111111111111111111111111111111111110000000000000000000000010000000000;
		39580: Delta = 69'sb000000000000000000000000000000000001111111111111111111111110000000000;
		9233: Delta = 69'sb111111111111111111111111111111111101111111111111111111111110000000000;
		31371: Delta = 69'sb000000000000000000000000000000000100000000000000000000000010000000000;
		21538: Delta = 69'sb111111111111111111111111111111111100000000000000000000000010000000000;
		29323: Delta = 69'sb000000000000000000000000000000000011111111111111111111111110000000000;
		19490: Delta = 69'sb111111111111111111111111111111111011111111111111111111111110000000000;
		10857: Delta = 69'sb000000000000000000000000000000001000000000000000000000000010000000000;
		42052: Delta = 69'sb111111111111111111111111111111111000000000000000000000000010000000000;
		8809: Delta = 69'sb000000000000000000000000000000000111111111111111111111111110000000000;
		40004: Delta = 69'sb111111111111111111111111111111110111111111111111111111111110000000000;
		20690: Delta = 69'sb000000000000000000000000000000010000000000000000000000000010000000000;
		32219: Delta = 69'sb111111111111111111111111111111110000000000000000000000000010000000000;
		18642: Delta = 69'sb000000000000000000000000000000001111111111111111111111111110000000000;
		30171: Delta = 69'sb111111111111111111111111111111101111111111111111111111111110000000000;
		40356: Delta = 69'sb000000000000000000000000000000100000000000000000000000000010000000000;
		12553: Delta = 69'sb111111111111111111111111111111100000000000000000000000000010000000000;
		38308: Delta = 69'sb000000000000000000000000000000011111111111111111111111111110000000000;
		10505: Delta = 69'sb111111111111111111111111111111011111111111111111111111111110000000000;
		28827: Delta = 69'sb000000000000000000000000000001000000000000000000000000000010000000000;
		24082: Delta = 69'sb111111111111111111111111111111000000000000000000000000000010000000000;
		26779: Delta = 69'sb000000000000000000000000000000111111111111111111111111111110000000000;
		22034: Delta = 69'sb111111111111111111111111111110111111111111111111111111111110000000000;
		5769: Delta = 69'sb000000000000000000000000000010000000000000000000000000000010000000000;
		47140: Delta = 69'sb111111111111111111111111111110000000000000000000000000000010000000000;
		3721: Delta = 69'sb000000000000000000000000000001111111111111111111111111111110000000000;
		45092: Delta = 69'sb111111111111111111111111111101111111111111111111111111111110000000000;
		10514: Delta = 69'sb000000000000000000000000000100000000000000000000000000000010000000000;
		42395: Delta = 69'sb111111111111111111111111111100000000000000000000000000000010000000000;
		8466: Delta = 69'sb000000000000000000000000000011111111111111111111111111111110000000000;
		40347: Delta = 69'sb111111111111111111111111111011111111111111111111111111111110000000000;
		20004: Delta = 69'sb000000000000000000000000001000000000000000000000000000000010000000000;
		32905: Delta = 69'sb111111111111111111111111111000000000000000000000000000000010000000000;
		17956: Delta = 69'sb000000000000000000000000000111111111111111111111111111111110000000000;
		30857: Delta = 69'sb111111111111111111111111110111111111111111111111111111111110000000000;
		38984: Delta = 69'sb000000000000000000000000010000000000000000000000000000000010000000000;
		13925: Delta = 69'sb111111111111111111111111110000000000000000000000000000000010000000000;
		36936: Delta = 69'sb000000000000000000000000001111111111111111111111111111111110000000000;
		11877: Delta = 69'sb111111111111111111111111101111111111111111111111111111111110000000000;
		26083: Delta = 69'sb000000000000000000000000100000000000000000000000000000000010000000000;
		26826: Delta = 69'sb111111111111111111111111100000000000000000000000000000000010000000000;
		24035: Delta = 69'sb000000000000000000000000011111111111111111111111111111111110000000000;
		24778: Delta = 69'sb111111111111111111111111011111111111111111111111111111111110000000000;
		281: Delta = 69'sb000000000000000000000001000000000000000000000000000000000010000000000;
		1767: Delta = 69'sb111111111111111111111111000000000000000000000000000000000010000000000;
		49094: Delta = 69'sb000000000000000000000000111111111111111111111111111111111110000000000;
		50580: Delta = 69'sb111111111111111111111110111111111111111111111111111111111110000000000;
		50399: Delta = 69'sb000000000000000000000010000000000000000000000000000000000010000000000;
		2510: Delta = 69'sb111111111111111111111110000000000000000000000000000000000010000000000;
		48351: Delta = 69'sb000000000000000000000001111111111111111111111111111111111110000000000;
		462: Delta = 69'sb111111111111111111111101111111111111111111111111111111111110000000000;
		48913: Delta = 69'sb000000000000000000000100000000000000000000000000000000000010000000000;
		3996: Delta = 69'sb111111111111111111111100000000000000000000000000000000000010000000000;
		46865: Delta = 69'sb000000000000000000000011111111111111111111111111111111111110000000000;
		1948: Delta = 69'sb111111111111111111111011111111111111111111111111111111111110000000000;
		45941: Delta = 69'sb000000000000000000001000000000000000000000000000000000000010000000000;
		6968: Delta = 69'sb111111111111111111111000000000000000000000000000000000000010000000000;
		43893: Delta = 69'sb000000000000000000000111111111111111111111111111111111111110000000000;
		4920: Delta = 69'sb111111111111111111110111111111111111111111111111111111111110000000000;
		39997: Delta = 69'sb000000000000000000010000000000000000000000000000000000000010000000000;
		12912: Delta = 69'sb111111111111111111110000000000000000000000000000000000000010000000000;
		37949: Delta = 69'sb000000000000000000001111111111111111111111111111111111111110000000000;
		10864: Delta = 69'sb111111111111111111101111111111111111111111111111111111111110000000000;
		28109: Delta = 69'sb000000000000000000100000000000000000000000000000000000000010000000000;
		24800: Delta = 69'sb111111111111111111100000000000000000000000000000000000000010000000000;
		26061: Delta = 69'sb000000000000000000011111111111111111111111111111111111111110000000000;
		22752: Delta = 69'sb111111111111111111011111111111111111111111111111111111111110000000000;
		4333: Delta = 69'sb000000000000000001000000000000000000000000000000000000000010000000000;
		48576: Delta = 69'sb111111111111111111000000000000000000000000000000000000000010000000000;
		2285: Delta = 69'sb000000000000000000111111111111111111111111111111111111111110000000000;
		46528: Delta = 69'sb111111111111111110111111111111111111111111111111111111111110000000000;
		7642: Delta = 69'sb000000000000000010000000000000000000000000000000000000000010000000000;
		45267: Delta = 69'sb111111111111111110000000000000000000000000000000000000000010000000000;
		5594: Delta = 69'sb000000000000000001111111111111111111111111111111111111111110000000000;
		43219: Delta = 69'sb111111111111111101111111111111111111111111111111111111111110000000000;
		14260: Delta = 69'sb000000000000000100000000000000000000000000000000000000000010000000000;
		38649: Delta = 69'sb111111111111111100000000000000000000000000000000000000000010000000000;
		12212: Delta = 69'sb000000000000000011111111111111111111111111111111111111111110000000000;
		36601: Delta = 69'sb111111111111111011111111111111111111111111111111111111111110000000000;
		27496: Delta = 69'sb000000000000001000000000000000000000000000000000000000000010000000000;
		25413: Delta = 69'sb111111111111111000000000000000000000000000000000000000000010000000000;
		25448: Delta = 69'sb000000000000000111111111111111111111111111111111111111111110000000000;
		23365: Delta = 69'sb111111111111110111111111111111111111111111111111111111111110000000000;
		3107: Delta = 69'sb000000000000010000000000000000000000000000000000000000000010000000000;
		49802: Delta = 69'sb111111111111110000000000000000000000000000000000000000000010000000000;
		1059: Delta = 69'sb000000000000001111111111111111111111111111111111111111111110000000000;
		47754: Delta = 69'sb111111111111101111111111111111111111111111111111111111111110000000000;
		5190: Delta = 69'sb000000000000100000000000000000000000000000000000000000000010000000000;
		47719: Delta = 69'sb111111111111100000000000000000000000000000000000000000000010000000000;
		3142: Delta = 69'sb000000000000011111111111111111111111111111111111111111111110000000000;
		45671: Delta = 69'sb111111111111011111111111111111111111111111111111111111111110000000000;
		9356: Delta = 69'sb000000000001000000000000000000000000000000000000000000000010000000000;
		43553: Delta = 69'sb111111111111000000000000000000000000000000000000000000000010000000000;
		7308: Delta = 69'sb000000000000111111111111111111111111111111111111111111111110000000000;
		41505: Delta = 69'sb111111111110111111111111111111111111111111111111111111111110000000000;
		17688: Delta = 69'sb000000000010000000000000000000000000000000000000000000000010000000000;
		35221: Delta = 69'sb111111111110000000000000000000000000000000000000000000000010000000000;
		15640: Delta = 69'sb000000000001111111111111111111111111111111111111111111111110000000000;
		33173: Delta = 69'sb111111111101111111111111111111111111111111111111111111111110000000000;
		34352: Delta = 69'sb000000000100000000000000000000000000000000000000000000000010000000000;
		18557: Delta = 69'sb111111111100000000000000000000000000000000000000000000000010000000000;
		32304: Delta = 69'sb000000000011111111111111111111111111111111111111111111111110000000000;
		16509: Delta = 69'sb111111111011111111111111111111111111111111111111111111111110000000000;
		16819: Delta = 69'sb000000001000000000000000000000000000000000000000000000000010000000000;
		36090: Delta = 69'sb111111111000000000000000000000000000000000000000000000000010000000000;
		14771: Delta = 69'sb000000000111111111111111111111111111111111111111111111111110000000000;
		34042: Delta = 69'sb111111110111111111111111111111111111111111111111111111111110000000000;
		32614: Delta = 69'sb000000010000000000000000000000000000000000000000000000000010000000000;
		20295: Delta = 69'sb111111110000000000000000000000000000000000000000000000000010000000000;
		30566: Delta = 69'sb000000001111111111111111111111111111111111111111111111111110000000000;
		18247: Delta = 69'sb111111101111111111111111111111111111111111111111111111111110000000000;
		13343: Delta = 69'sb000000100000000000000000000000000000000000000000000000000010000000000;
		39566: Delta = 69'sb111111100000000000000000000000000000000000000000000000000010000000000;
		11295: Delta = 69'sb000000011111111111111111111111111111111111111111111111111110000000000;
		37518: Delta = 69'sb111111011111111111111111111111111111111111111111111111111110000000000;
		25662: Delta = 69'sb000001000000000000000000000000000000000000000000000000000010000000000;
		27247: Delta = 69'sb111111000000000000000000000000000000000000000000000000000010000000000;
		23614: Delta = 69'sb000000111111111111111111111111111111111111111111111111111110000000000;
		25199: Delta = 69'sb111110111111111111111111111111111111111111111111111111111110000000000;
		50300: Delta = 69'sb000010000000000000000000000000000000000000000000000000000010000000000;
		2609: Delta = 69'sb111110000000000000000000000000000000000000000000000000000010000000000;
		48252: Delta = 69'sb000001111111111111111111111111111111111111111111111111111110000000000;
		561: Delta = 69'sb111101111111111111111111111111111111111111111111111111111110000000000;
		48715: Delta = 69'sb000100000000000000000000000000000000000000000000000000000010000000000;
		4194: Delta = 69'sb111100000000000000000000000000000000000000000000000000000010000000000;
		46667: Delta = 69'sb000011111111111111111111111111111111111111111111111111111110000000000;
		2146: Delta = 69'sb111011111111111111111111111111111111111111111111111111111110000000000;
		45545: Delta = 69'sb001000000000000000000000000000000000000000000000000000000010000000000;
		7364: Delta = 69'sb111000000000000000000000000000000000000000000000000000000010000000000;
		43497: Delta = 69'sb000111111111111111111111111111111111111111111111111111111110000000000;
		5316: Delta = 69'sb110111111111111111111111111111111111111111111111111111111110000000000;
		39205: Delta = 69'sb010000000000000000000000000000000000000000000000000000000010000000000;
		13704: Delta = 69'sb110000000000000000000000000000000000000000000000000000000010000000000;
		37157: Delta = 69'sb001111111111111111111111111111111111111111111111111111111110000000000;
		11656: Delta = 69'sb101111111111111111111111111111111111111111111111111111111110000000000;
		6144: Delta = 69'sb000000000000000000000000000000000000000000000000000000001100000000000;
		44717: Delta = 69'sb111111111111111111111111111111111111111111111111111111110100000000000;
		10240: Delta = 69'sb000000000000000000000000000000000000000000000000000000010100000000000;
		40621: Delta = 69'sb111111111111111111111111111111111111111111111111111111101100000000000;
		18432: Delta = 69'sb000000000000000000000000000000000000000000000000000000100100000000000;
		36525: Delta = 69'sb111111111111111111111111111111111111111111111111111111100100000000000;
		14336: Delta = 69'sb000000000000000000000000000000000000000000000000000000011100000000000;
		32429: Delta = 69'sb111111111111111111111111111111111111111111111111111111011100000000000;
		34816: Delta = 69'sb000000000000000000000000000000000000000000000000000001000100000000000;
		20141: Delta = 69'sb111111111111111111111111111111111111111111111111111111000100000000000;
		30720: Delta = 69'sb000000000000000000000000000000000000000000000000000000111100000000000;
		16045: Delta = 69'sb111111111111111111111111111111111111111111111111111110111100000000000;
		16723: Delta = 69'sb000000000000000000000000000000000000000000000000000010000100000000000;
		38234: Delta = 69'sb111111111111111111111111111111111111111111111111111110000100000000000;
		12627: Delta = 69'sb000000000000000000000000000000000000000000000000000001111100000000000;
		34138: Delta = 69'sb111111111111111111111111111111111111111111111111111101111100000000000;
		31398: Delta = 69'sb000000000000000000000000000000000000000000000000000100000100000000000;
		23559: Delta = 69'sb111111111111111111111111111111111111111111111111111100000100000000000;
		27302: Delta = 69'sb000000000000000000000000000000000000000000000000000011111100000000000;
		19463: Delta = 69'sb111111111111111111111111111111111111111111111111111011111100000000000;
		9887: Delta = 69'sb000000000000000000000000000000000000000000000000001000000100000000000;
		45070: Delta = 69'sb111111111111111111111111111111111111111111111111111000000100000000000;
		5791: Delta = 69'sb000000000000000000000000000000000000000000000000000111111100000000000;
		40974: Delta = 69'sb111111111111111111111111111111111111111111111111110111111100000000000;
		17726: Delta = 69'sb000000000000000000000000000000000000000000000000010000000100000000000;
		37231: Delta = 69'sb111111111111111111111111111111111111111111111111110000000100000000000;
		13630: Delta = 69'sb000000000000000000000000000000000000000000000000001111111100000000000;
		33135: Delta = 69'sb111111111111111111111111111111111111111111111111101111111100000000000;
		33404: Delta = 69'sb000000000000000000000000000000000000000000000000100000000100000000000;
		21553: Delta = 69'sb111111111111111111111111111111111111111111111111100000000100000000000;
		29308: Delta = 69'sb000000000000000000000000000000000000000000000000011111111100000000000;
		17457: Delta = 69'sb111111111111111111111111111111111111111111111111011111111100000000000;
		13899: Delta = 69'sb000000000000000000000000000000000000000000000001000000000100000000000;
		41058: Delta = 69'sb111111111111111111111111111111111111111111111111000000000100000000000;
		9803: Delta = 69'sb000000000000000000000000000000000000000000000000111111111100000000000;
		36962: Delta = 69'sb111111111111111111111111111111111111111111111110111111111100000000000;
		25750: Delta = 69'sb000000000000000000000000000000000000000000000010000000000100000000000;
		29207: Delta = 69'sb111111111111111111111111111111111111111111111110000000000100000000000;
		21654: Delta = 69'sb000000000000000000000000000000000000000000000001111111111100000000000;
		25111: Delta = 69'sb111111111111111111111111111111111111111111111101111111111100000000000;
		49452: Delta = 69'sb000000000000000000000000000000000000000000000100000000000100000000000;
		5505: Delta = 69'sb111111111111111111111111111111111111111111111100000000000100000000000;
		45356: Delta = 69'sb000000000000000000000000000000000000000000000011111111111100000000000;
		1409: Delta = 69'sb111111111111111111111111111111111111111111111011111111111100000000000;
		45995: Delta = 69'sb000000000000000000000000000000000000000000001000000000000100000000000;
		8962: Delta = 69'sb111111111111111111111111111111111111111111111000000000000100000000000;
		41899: Delta = 69'sb000000000000000000000000000000000000000000000111111111111100000000000;
		4866: Delta = 69'sb111111111111111111111111111111111111111111110111111111111100000000000;
		39081: Delta = 69'sb000000000000000000000000000000000000000000010000000000000100000000000;
		15876: Delta = 69'sb111111111111111111111111111111111111111111110000000000000100000000000;
		34985: Delta = 69'sb000000000000000000000000000000000000000000001111111111111100000000000;
		11780: Delta = 69'sb111111111111111111111111111111111111111111101111111111111100000000000;
		25253: Delta = 69'sb000000000000000000000000000000000000000000100000000000000100000000000;
		29704: Delta = 69'sb111111111111111111111111111111111111111111100000000000000100000000000;
		21157: Delta = 69'sb000000000000000000000000000000000000000000011111111111111100000000000;
		25608: Delta = 69'sb111111111111111111111111111111111111111111011111111111111100000000000;
		48458: Delta = 69'sb000000000000000000000000000000000000000001000000000000000100000000000;
		6499: Delta = 69'sb111111111111111111111111111111111111111111000000000000000100000000000;
		44362: Delta = 69'sb000000000000000000000000000000000000000000111111111111111100000000000;
		2403: Delta = 69'sb111111111111111111111111111111111111111110111111111111111100000000000;
		44007: Delta = 69'sb000000000000000000000000000000000000000010000000000000000100000000000;
		10950: Delta = 69'sb111111111111111111111111111111111111111110000000000000000100000000000;
		39911: Delta = 69'sb000000000000000000000000000000000000000001111111111111111100000000000;
		6854: Delta = 69'sb111111111111111111111111111111111111111101111111111111111100000000000;
		35105: Delta = 69'sb000000000000000000000000000000000000000100000000000000000100000000000;
		19852: Delta = 69'sb111111111111111111111111111111111111111100000000000000000100000000000;
		31009: Delta = 69'sb000000000000000000000000000000000000000011111111111111111100000000000;
		15756: Delta = 69'sb111111111111111111111111111111111111111011111111111111111100000000000;
		17301: Delta = 69'sb000000000000000000000000000000000000001000000000000000000100000000000;
		37656: Delta = 69'sb111111111111111111111111111111111111111000000000000000000100000000000;
		13205: Delta = 69'sb000000000000000000000000000000000000000111111111111111111100000000000;
		33560: Delta = 69'sb111111111111111111111111111111111111110111111111111111111100000000000;
		32554: Delta = 69'sb000000000000000000000000000000000000010000000000000000000100000000000;
		22403: Delta = 69'sb111111111111111111111111111111111111110000000000000000000100000000000;
		28458: Delta = 69'sb000000000000000000000000000000000000001111111111111111111100000000000;
		18307: Delta = 69'sb111111111111111111111111111111111111101111111111111111111100000000000;
		12199: Delta = 69'sb000000000000000000000000000000000000100000000000000000000100000000000;
		42758: Delta = 69'sb111111111111111111111111111111111111100000000000000000000100000000000;
		8103: Delta = 69'sb000000000000000000000000000000000000011111111111111111111100000000000;
		38662: Delta = 69'sb111111111111111111111111111111111111011111111111111111111100000000000;
		22350: Delta = 69'sb000000000000000000000000000000000001000000000000000000000100000000000;
		32607: Delta = 69'sb111111111111111111111111111111111111000000000000000000000100000000000;
		18254: Delta = 69'sb000000000000000000000000000000000000111111111111111111111100000000000;
		28511: Delta = 69'sb111111111111111111111111111111111110111111111111111111111100000000000;
		42652: Delta = 69'sb000000000000000000000000000000000010000000000000000000000100000000000;
		12305: Delta = 69'sb111111111111111111111111111111111110000000000000000000000100000000000;
		38556: Delta = 69'sb000000000000000000000000000000000001111111111111111111111100000000000;
		8209: Delta = 69'sb111111111111111111111111111111111101111111111111111111111100000000000;
		32395: Delta = 69'sb000000000000000000000000000000000100000000000000000000000100000000000;
		22562: Delta = 69'sb111111111111111111111111111111111100000000000000000000000100000000000;
		28299: Delta = 69'sb000000000000000000000000000000000011111111111111111111111100000000000;
		18466: Delta = 69'sb111111111111111111111111111111111011111111111111111111111100000000000;
		11881: Delta = 69'sb000000000000000000000000000000001000000000000000000000000100000000000;
		43076: Delta = 69'sb111111111111111111111111111111111000000000000000000000000100000000000;
		7785: Delta = 69'sb000000000000000000000000000000000111111111111111111111111100000000000;
		38980: Delta = 69'sb111111111111111111111111111111110111111111111111111111111100000000000;
		21714: Delta = 69'sb000000000000000000000000000000010000000000000000000000000100000000000;
		33243: Delta = 69'sb111111111111111111111111111111110000000000000000000000000100000000000;
		17618: Delta = 69'sb000000000000000000000000000000001111111111111111111111111100000000000;
		29147: Delta = 69'sb111111111111111111111111111111101111111111111111111111111100000000000;
		41380: Delta = 69'sb000000000000000000000000000000100000000000000000000000000100000000000;
		13577: Delta = 69'sb111111111111111111111111111111100000000000000000000000000100000000000;
		37284: Delta = 69'sb000000000000000000000000000000011111111111111111111111111100000000000;
		9481: Delta = 69'sb111111111111111111111111111111011111111111111111111111111100000000000;
		29851: Delta = 69'sb000000000000000000000000000001000000000000000000000000000100000000000;
		25106: Delta = 69'sb111111111111111111111111111111000000000000000000000000000100000000000;
		25755: Delta = 69'sb000000000000000000000000000000111111111111111111111111111100000000000;
		21010: Delta = 69'sb111111111111111111111111111110111111111111111111111111111100000000000;
		6793: Delta = 69'sb000000000000000000000000000010000000000000000000000000000100000000000;
		48164: Delta = 69'sb111111111111111111111111111110000000000000000000000000000100000000000;
		2697: Delta = 69'sb000000000000000000000000000001111111111111111111111111111100000000000;
		44068: Delta = 69'sb111111111111111111111111111101111111111111111111111111111100000000000;
		11538: Delta = 69'sb000000000000000000000000000100000000000000000000000000000100000000000;
		43419: Delta = 69'sb111111111111111111111111111100000000000000000000000000000100000000000;
		7442: Delta = 69'sb000000000000000000000000000011111111111111111111111111111100000000000;
		39323: Delta = 69'sb111111111111111111111111111011111111111111111111111111111100000000000;
		21028: Delta = 69'sb000000000000000000000000001000000000000000000000000000000100000000000;
		33929: Delta = 69'sb111111111111111111111111111000000000000000000000000000000100000000000;
		16932: Delta = 69'sb000000000000000000000000000111111111111111111111111111111100000000000;
		29833: Delta = 69'sb111111111111111111111111110111111111111111111111111111111100000000000;
		40008: Delta = 69'sb000000000000000000000000010000000000000000000000000000000100000000000;
		14949: Delta = 69'sb111111111111111111111111110000000000000000000000000000000100000000000;
		35912: Delta = 69'sb000000000000000000000000001111111111111111111111111111111100000000000;
		10853: Delta = 69'sb111111111111111111111111101111111111111111111111111111111100000000000;
		27107: Delta = 69'sb000000000000000000000000100000000000000000000000000000000100000000000;
		27850: Delta = 69'sb111111111111111111111111100000000000000000000000000000000100000000000;
		23011: Delta = 69'sb000000000000000000000000011111111111111111111111111111111100000000000;
		23754: Delta = 69'sb111111111111111111111111011111111111111111111111111111111100000000000;
		1305: Delta = 69'sb000000000000000000000001000000000000000000000000000000000100000000000;
		2791: Delta = 69'sb111111111111111111111111000000000000000000000000000000000100000000000;
		48070: Delta = 69'sb000000000000000000000000111111111111111111111111111111111100000000000;
		49556: Delta = 69'sb111111111111111111111110111111111111111111111111111111111100000000000;
		562: Delta = 69'sb000000000000000000000010000000000000000000000000000000000100000000000;
		3534: Delta = 69'sb111111111111111111111110000000000000000000000000000000000100000000000;
		47327: Delta = 69'sb000000000000000000000001111111111111111111111111111111111100000000000;
		50299: Delta = 69'sb111111111111111111111101111111111111111111111111111111111100000000000;
		49937: Delta = 69'sb000000000000000000000100000000000000000000000000000000000100000000000;
		5020: Delta = 69'sb111111111111111111111100000000000000000000000000000000000100000000000;
		45841: Delta = 69'sb000000000000000000000011111111111111111111111111111111111100000000000;
		924: Delta = 69'sb111111111111111111111011111111111111111111111111111111111100000000000;
		46965: Delta = 69'sb000000000000000000001000000000000000000000000000000000000100000000000;
		7992: Delta = 69'sb111111111111111111111000000000000000000000000000000000000100000000000;
		42869: Delta = 69'sb000000000000000000000111111111111111111111111111111111111100000000000;
		3896: Delta = 69'sb111111111111111111110111111111111111111111111111111111111100000000000;
		41021: Delta = 69'sb000000000000000000010000000000000000000000000000000000000100000000000;
		13936: Delta = 69'sb111111111111111111110000000000000000000000000000000000000100000000000;
		36925: Delta = 69'sb000000000000000000001111111111111111111111111111111111111100000000000;
		9840: Delta = 69'sb111111111111111111101111111111111111111111111111111111111100000000000;
		29133: Delta = 69'sb000000000000000000100000000000000000000000000000000000000100000000000;
		25824: Delta = 69'sb111111111111111111100000000000000000000000000000000000000100000000000;
		25037: Delta = 69'sb000000000000000000011111111111111111111111111111111111111100000000000;
		21728: Delta = 69'sb111111111111111111011111111111111111111111111111111111111100000000000;
		5357: Delta = 69'sb000000000000000001000000000000000000000000000000000000000100000000000;
		49600: Delta = 69'sb111111111111111111000000000000000000000000000000000000000100000000000;
		1261: Delta = 69'sb000000000000000000111111111111111111111111111111111111111100000000000;
		45504: Delta = 69'sb111111111111111110111111111111111111111111111111111111111100000000000;
		8666: Delta = 69'sb000000000000000010000000000000000000000000000000000000000100000000000;
		46291: Delta = 69'sb111111111111111110000000000000000000000000000000000000000100000000000;
		4570: Delta = 69'sb000000000000000001111111111111111111111111111111111111111100000000000;
		42195: Delta = 69'sb111111111111111101111111111111111111111111111111111111111100000000000;
		15284: Delta = 69'sb000000000000000100000000000000000000000000000000000000000100000000000;
		39673: Delta = 69'sb111111111111111100000000000000000000000000000000000000000100000000000;
		11188: Delta = 69'sb000000000000000011111111111111111111111111111111111111111100000000000;
		35577: Delta = 69'sb111111111111111011111111111111111111111111111111111111111100000000000;
		28520: Delta = 69'sb000000000000001000000000000000000000000000000000000000000100000000000;
		26437: Delta = 69'sb111111111111111000000000000000000000000000000000000000000100000000000;
		24424: Delta = 69'sb000000000000000111111111111111111111111111111111111111111100000000000;
		22341: Delta = 69'sb111111111111110111111111111111111111111111111111111111111100000000000;
		4131: Delta = 69'sb000000000000010000000000000000000000000000000000000000000100000000000;
		50826: Delta = 69'sb111111111111110000000000000000000000000000000000000000000100000000000;
		35: Delta = 69'sb000000000000001111111111111111111111111111111111111111111100000000000;
		46730: Delta = 69'sb111111111111101111111111111111111111111111111111111111111100000000000;
		6214: Delta = 69'sb000000000000100000000000000000000000000000000000000000000100000000000;
		48743: Delta = 69'sb111111111111100000000000000000000000000000000000000000000100000000000;
		2118: Delta = 69'sb000000000000011111111111111111111111111111111111111111111100000000000;
		44647: Delta = 69'sb111111111111011111111111111111111111111111111111111111111100000000000;
		10380: Delta = 69'sb000000000001000000000000000000000000000000000000000000000100000000000;
		44577: Delta = 69'sb111111111111000000000000000000000000000000000000000000000100000000000;
		6284: Delta = 69'sb000000000000111111111111111111111111111111111111111111111100000000000;
		40481: Delta = 69'sb111111111110111111111111111111111111111111111111111111111100000000000;
		18712: Delta = 69'sb000000000010000000000000000000000000000000000000000000000100000000000;
		36245: Delta = 69'sb111111111110000000000000000000000000000000000000000000000100000000000;
		14616: Delta = 69'sb000000000001111111111111111111111111111111111111111111111100000000000;
		32149: Delta = 69'sb111111111101111111111111111111111111111111111111111111111100000000000;
		35376: Delta = 69'sb000000000100000000000000000000000000000000000000000000000100000000000;
		19581: Delta = 69'sb111111111100000000000000000000000000000000000000000000000100000000000;
		31280: Delta = 69'sb000000000011111111111111111111111111111111111111111111111100000000000;
		15485: Delta = 69'sb111111111011111111111111111111111111111111111111111111111100000000000;
		17843: Delta = 69'sb000000001000000000000000000000000000000000000000000000000100000000000;
		37114: Delta = 69'sb111111111000000000000000000000000000000000000000000000000100000000000;
		13747: Delta = 69'sb000000000111111111111111111111111111111111111111111111111100000000000;
		33018: Delta = 69'sb111111110111111111111111111111111111111111111111111111111100000000000;
		33638: Delta = 69'sb000000010000000000000000000000000000000000000000000000000100000000000;
		21319: Delta = 69'sb111111110000000000000000000000000000000000000000000000000100000000000;
		29542: Delta = 69'sb000000001111111111111111111111111111111111111111111111111100000000000;
		17223: Delta = 69'sb111111101111111111111111111111111111111111111111111111111100000000000;
		14367: Delta = 69'sb000000100000000000000000000000000000000000000000000000000100000000000;
		40590: Delta = 69'sb111111100000000000000000000000000000000000000000000000000100000000000;
		10271: Delta = 69'sb000000011111111111111111111111111111111111111111111111111100000000000;
		36494: Delta = 69'sb111111011111111111111111111111111111111111111111111111111100000000000;
		26686: Delta = 69'sb000001000000000000000000000000000000000000000000000000000100000000000;
		28271: Delta = 69'sb111111000000000000000000000000000000000000000000000000000100000000000;
		22590: Delta = 69'sb000000111111111111111111111111111111111111111111111111111100000000000;
		24175: Delta = 69'sb111110111111111111111111111111111111111111111111111111111100000000000;
		463: Delta = 69'sb000010000000000000000000000000000000000000000000000000000100000000000;
		3633: Delta = 69'sb111110000000000000000000000000000000000000000000000000000100000000000;
		47228: Delta = 69'sb000001111111111111111111111111111111111111111111111111111100000000000;
		50398: Delta = 69'sb111101111111111111111111111111111111111111111111111111111100000000000;
		49739: Delta = 69'sb000100000000000000000000000000000000000000000000000000000100000000000;
		5218: Delta = 69'sb111100000000000000000000000000000000000000000000000000000100000000000;
		45643: Delta = 69'sb000011111111111111111111111111111111111111111111111111111100000000000;
		1122: Delta = 69'sb111011111111111111111111111111111111111111111111111111111100000000000;
		46569: Delta = 69'sb001000000000000000000000000000000000000000000000000000000100000000000;
		8388: Delta = 69'sb111000000000000000000000000000000000000000000000000000000100000000000;
		42473: Delta = 69'sb000111111111111111111111111111111111111111111111111111111100000000000;
		4292: Delta = 69'sb110111111111111111111111111111111111111111111111111111111100000000000;
		40229: Delta = 69'sb010000000000000000000000000000000000000000000000000000000100000000000;
		14728: Delta = 69'sb110000000000000000000000000000000000000000000000000000000100000000000;
		36133: Delta = 69'sb001111111111111111111111111111111111111111111111111111111100000000000;
		10632: Delta = 69'sb101111111111111111111111111111111111111111111111111111111100000000000;
		12288: Delta = 69'sb000000000000000000000000000000000000000000000000000000011000000000000;
		38573: Delta = 69'sb111111111111111111111111111111111111111111111111111111101000000000000;
		20480: Delta = 69'sb000000000000000000000000000000000000000000000000000000101000000000000;
		30381: Delta = 69'sb111111111111111111111111111111111111111111111111111111011000000000000;
		36864: Delta = 69'sb000000000000000000000000000000000000000000000000000001001000000000000;
		22189: Delta = 69'sb111111111111111111111111111111111111111111111111111111001000000000000;
		28672: Delta = 69'sb000000000000000000000000000000000000000000000000000000111000000000000;
		13997: Delta = 69'sb111111111111111111111111111111111111111111111111111110111000000000000;
		18771: Delta = 69'sb000000000000000000000000000000000000000000000000000010001000000000000;
		40282: Delta = 69'sb111111111111111111111111111111111111111111111111111110001000000000000;
		10579: Delta = 69'sb000000000000000000000000000000000000000000000000000001111000000000000;
		32090: Delta = 69'sb111111111111111111111111111111111111111111111111111101111000000000000;
		33446: Delta = 69'sb000000000000000000000000000000000000000000000000000100001000000000000;
		25607: Delta = 69'sb111111111111111111111111111111111111111111111111111100001000000000000;
		25254: Delta = 69'sb000000000000000000000000000000000000000000000000000011111000000000000;
		17415: Delta = 69'sb111111111111111111111111111111111111111111111111111011111000000000000;
		11935: Delta = 69'sb000000000000000000000000000000000000000000000000001000001000000000000;
		47118: Delta = 69'sb111111111111111111111111111111111111111111111111111000001000000000000;
		3743: Delta = 69'sb000000000000000000000000000000000000000000000000000111111000000000000;
		38926: Delta = 69'sb111111111111111111111111111111111111111111111111110111111000000000000;
		19774: Delta = 69'sb000000000000000000000000000000000000000000000000010000001000000000000;
		39279: Delta = 69'sb111111111111111111111111111111111111111111111111110000001000000000000;
		11582: Delta = 69'sb000000000000000000000000000000000000000000000000001111111000000000000;
		31087: Delta = 69'sb111111111111111111111111111111111111111111111111101111111000000000000;
		35452: Delta = 69'sb000000000000000000000000000000000000000000000000100000001000000000000;
		23601: Delta = 69'sb111111111111111111111111111111111111111111111111100000001000000000000;
		27260: Delta = 69'sb000000000000000000000000000000000000000000000000011111111000000000000;
		15409: Delta = 69'sb111111111111111111111111111111111111111111111111011111111000000000000;
		15947: Delta = 69'sb000000000000000000000000000000000000000000000001000000001000000000000;
		43106: Delta = 69'sb111111111111111111111111111111111111111111111111000000001000000000000;
		7755: Delta = 69'sb000000000000000000000000000000000000000000000000111111111000000000000;
		34914: Delta = 69'sb111111111111111111111111111111111111111111111110111111111000000000000;
		27798: Delta = 69'sb000000000000000000000000000000000000000000000010000000001000000000000;
		31255: Delta = 69'sb111111111111111111111111111111111111111111111110000000001000000000000;
		19606: Delta = 69'sb000000000000000000000000000000000000000000000001111111111000000000000;
		23063: Delta = 69'sb111111111111111111111111111111111111111111111101111111111000000000000;
		639: Delta = 69'sb000000000000000000000000000000000000000000000100000000001000000000000;
		7553: Delta = 69'sb111111111111111111111111111111111111111111111100000000001000000000000;
		43308: Delta = 69'sb000000000000000000000000000000000000000000000011111111111000000000000;
		50222: Delta = 69'sb111111111111111111111111111111111111111111111011111111111000000000000;
		48043: Delta = 69'sb000000000000000000000000000000000000000000001000000000001000000000000;
		11010: Delta = 69'sb111111111111111111111111111111111111111111111000000000001000000000000;
		39851: Delta = 69'sb000000000000000000000000000000000000000000000111111111111000000000000;
		2818: Delta = 69'sb111111111111111111111111111111111111111111110111111111111000000000000;
		41129: Delta = 69'sb000000000000000000000000000000000000000000010000000000001000000000000;
		17924: Delta = 69'sb111111111111111111111111111111111111111111110000000000001000000000000;
		32937: Delta = 69'sb000000000000000000000000000000000000000000001111111111111000000000000;
		9732: Delta = 69'sb111111111111111111111111111111111111111111101111111111111000000000000;
		27301: Delta = 69'sb000000000000000000000000000000000000000000100000000000001000000000000;
		31752: Delta = 69'sb111111111111111111111111111111111111111111100000000000001000000000000;
		19109: Delta = 69'sb000000000000000000000000000000000000000000011111111111111000000000000;
		23560: Delta = 69'sb111111111111111111111111111111111111111111011111111111111000000000000;
		50506: Delta = 69'sb000000000000000000000000000000000000000001000000000000001000000000000;
		8547: Delta = 69'sb111111111111111111111111111111111111111111000000000000001000000000000;
		42314: Delta = 69'sb000000000000000000000000000000000000000000111111111111111000000000000;
		355: Delta = 69'sb111111111111111111111111111111111111111110111111111111111000000000000;
		46055: Delta = 69'sb000000000000000000000000000000000000000010000000000000001000000000000;
		12998: Delta = 69'sb111111111111111111111111111111111111111110000000000000001000000000000;
		37863: Delta = 69'sb000000000000000000000000000000000000000001111111111111111000000000000;
		4806: Delta = 69'sb111111111111111111111111111111111111111101111111111111111000000000000;
		37153: Delta = 69'sb000000000000000000000000000000000000000100000000000000001000000000000;
		21900: Delta = 69'sb111111111111111111111111111111111111111100000000000000001000000000000;
		28961: Delta = 69'sb000000000000000000000000000000000000000011111111111111111000000000000;
		13708: Delta = 69'sb111111111111111111111111111111111111111011111111111111111000000000000;
		19349: Delta = 69'sb000000000000000000000000000000000000001000000000000000001000000000000;
		39704: Delta = 69'sb111111111111111111111111111111111111111000000000000000001000000000000;
		11157: Delta = 69'sb000000000000000000000000000000000000000111111111111111111000000000000;
		31512: Delta = 69'sb111111111111111111111111111111111111110111111111111111111000000000000;
		34602: Delta = 69'sb000000000000000000000000000000000000010000000000000000001000000000000;
		24451: Delta = 69'sb111111111111111111111111111111111111110000000000000000001000000000000;
		26410: Delta = 69'sb000000000000000000000000000000000000001111111111111111111000000000000;
		16259: Delta = 69'sb111111111111111111111111111111111111101111111111111111111000000000000;
		14247: Delta = 69'sb000000000000000000000000000000000000100000000000000000001000000000000;
		44806: Delta = 69'sb111111111111111111111111111111111111100000000000000000001000000000000;
		6055: Delta = 69'sb000000000000000000000000000000000000011111111111111111111000000000000;
		36614: Delta = 69'sb111111111111111111111111111111111111011111111111111111111000000000000;
		24398: Delta = 69'sb000000000000000000000000000000000001000000000000000000001000000000000;
		34655: Delta = 69'sb111111111111111111111111111111111111000000000000000000001000000000000;
		16206: Delta = 69'sb000000000000000000000000000000000000111111111111111111111000000000000;
		26463: Delta = 69'sb111111111111111111111111111111111110111111111111111111111000000000000;
		44700: Delta = 69'sb000000000000000000000000000000000010000000000000000000001000000000000;
		14353: Delta = 69'sb111111111111111111111111111111111110000000000000000000001000000000000;
		36508: Delta = 69'sb000000000000000000000000000000000001111111111111111111111000000000000;
		6161: Delta = 69'sb111111111111111111111111111111111101111111111111111111111000000000000;
		34443: Delta = 69'sb000000000000000000000000000000000100000000000000000000001000000000000;
		24610: Delta = 69'sb111111111111111111111111111111111100000000000000000000001000000000000;
		26251: Delta = 69'sb000000000000000000000000000000000011111111111111111111111000000000000;
		16418: Delta = 69'sb111111111111111111111111111111111011111111111111111111111000000000000;
		13929: Delta = 69'sb000000000000000000000000000000001000000000000000000000001000000000000;
		45124: Delta = 69'sb111111111111111111111111111111111000000000000000000000001000000000000;
		5737: Delta = 69'sb000000000000000000000000000000000111111111111111111111111000000000000;
		36932: Delta = 69'sb111111111111111111111111111111110111111111111111111111111000000000000;
		23762: Delta = 69'sb000000000000000000000000000000010000000000000000000000001000000000000;
		35291: Delta = 69'sb111111111111111111111111111111110000000000000000000000001000000000000;
		15570: Delta = 69'sb000000000000000000000000000000001111111111111111111111111000000000000;
		27099: Delta = 69'sb111111111111111111111111111111101111111111111111111111111000000000000;
		43428: Delta = 69'sb000000000000000000000000000000100000000000000000000000001000000000000;
		15625: Delta = 69'sb111111111111111111111111111111100000000000000000000000001000000000000;
		35236: Delta = 69'sb000000000000000000000000000000011111111111111111111111111000000000000;
		7433: Delta = 69'sb111111111111111111111111111111011111111111111111111111111000000000000;
		31899: Delta = 69'sb000000000000000000000000000001000000000000000000000000001000000000000;
		27154: Delta = 69'sb111111111111111111111111111111000000000000000000000000001000000000000;
		23707: Delta = 69'sb000000000000000000000000000000111111111111111111111111111000000000000;
		18962: Delta = 69'sb111111111111111111111111111110111111111111111111111111111000000000000;
		8841: Delta = 69'sb000000000000000000000000000010000000000000000000000000001000000000000;
		50212: Delta = 69'sb111111111111111111111111111110000000000000000000000000001000000000000;
		649: Delta = 69'sb000000000000000000000000000001111111111111111111111111111000000000000;
		42020: Delta = 69'sb111111111111111111111111111101111111111111111111111111111000000000000;
		13586: Delta = 69'sb000000000000000000000000000100000000000000000000000000001000000000000;
		45467: Delta = 69'sb111111111111111111111111111100000000000000000000000000001000000000000;
		5394: Delta = 69'sb000000000000000000000000000011111111111111111111111111111000000000000;
		37275: Delta = 69'sb111111111111111111111111111011111111111111111111111111111000000000000;
		23076: Delta = 69'sb000000000000000000000000001000000000000000000000000000001000000000000;
		35977: Delta = 69'sb111111111111111111111111111000000000000000000000000000001000000000000;
		14884: Delta = 69'sb000000000000000000000000000111111111111111111111111111111000000000000;
		27785: Delta = 69'sb111111111111111111111111110111111111111111111111111111111000000000000;
		42056: Delta = 69'sb000000000000000000000000010000000000000000000000000000001000000000000;
		16997: Delta = 69'sb111111111111111111111111110000000000000000000000000000001000000000000;
		33864: Delta = 69'sb000000000000000000000000001111111111111111111111111111111000000000000;
		8805: Delta = 69'sb111111111111111111111111101111111111111111111111111111111000000000000;
		29155: Delta = 69'sb000000000000000000000000100000000000000000000000000000001000000000000;
		29898: Delta = 69'sb111111111111111111111111100000000000000000000000000000001000000000000;
		20963: Delta = 69'sb000000000000000000000000011111111111111111111111111111111000000000000;
		21706: Delta = 69'sb111111111111111111111111011111111111111111111111111111111000000000000;
		3353: Delta = 69'sb000000000000000000000001000000000000000000000000000000001000000000000;
		4839: Delta = 69'sb111111111111111111111111000000000000000000000000000000001000000000000;
		46022: Delta = 69'sb000000000000000000000000111111111111111111111111111111111000000000000;
		47508: Delta = 69'sb111111111111111111111110111111111111111111111111111111111000000000000;
		2610: Delta = 69'sb000000000000000000000010000000000000000000000000000000001000000000000;
		5582: Delta = 69'sb111111111111111111111110000000000000000000000000000000001000000000000;
		45279: Delta = 69'sb000000000000000000000001111111111111111111111111111111111000000000000;
		48251: Delta = 69'sb111111111111111111111101111111111111111111111111111111111000000000000;
		1124: Delta = 69'sb000000000000000000000100000000000000000000000000000000001000000000000;
		7068: Delta = 69'sb111111111111111111111100000000000000000000000000000000001000000000000;
		43793: Delta = 69'sb000000000000000000000011111111111111111111111111111111111000000000000;
		49737: Delta = 69'sb111111111111111111111011111111111111111111111111111111111000000000000;
		49013: Delta = 69'sb000000000000000000001000000000000000000000000000000000001000000000000;
		10040: Delta = 69'sb111111111111111111111000000000000000000000000000000000001000000000000;
		40821: Delta = 69'sb000000000000000000000111111111111111111111111111111111111000000000000;
		1848: Delta = 69'sb111111111111111111110111111111111111111111111111111111111000000000000;
		43069: Delta = 69'sb000000000000000000010000000000000000000000000000000000001000000000000;
		15984: Delta = 69'sb111111111111111111110000000000000000000000000000000000001000000000000;
		34877: Delta = 69'sb000000000000000000001111111111111111111111111111111111111000000000000;
		7792: Delta = 69'sb111111111111111111101111111111111111111111111111111111111000000000000;
		31181: Delta = 69'sb000000000000000000100000000000000000000000000000000000001000000000000;
		27872: Delta = 69'sb111111111111111111100000000000000000000000000000000000001000000000000;
		22989: Delta = 69'sb000000000000000000011111111111111111111111111111111111111000000000000;
		19680: Delta = 69'sb111111111111111111011111111111111111111111111111111111111000000000000;
		7405: Delta = 69'sb000000000000000001000000000000000000000000000000000000001000000000000;
		787: Delta = 69'sb111111111111111111000000000000000000000000000000000000001000000000000;
		50074: Delta = 69'sb000000000000000000111111111111111111111111111111111111111000000000000;
		43456: Delta = 69'sb111111111111111110111111111111111111111111111111111111111000000000000;
		10714: Delta = 69'sb000000000000000010000000000000000000000000000000000000001000000000000;
		48339: Delta = 69'sb111111111111111110000000000000000000000000000000000000001000000000000;
		2522: Delta = 69'sb000000000000000001111111111111111111111111111111111111111000000000000;
		40147: Delta = 69'sb111111111111111101111111111111111111111111111111111111111000000000000;
		17332: Delta = 69'sb000000000000000100000000000000000000000000000000000000001000000000000;
		41721: Delta = 69'sb111111111111111100000000000000000000000000000000000000001000000000000;
		9140: Delta = 69'sb000000000000000011111111111111111111111111111111111111111000000000000;
		33529: Delta = 69'sb111111111111111011111111111111111111111111111111111111111000000000000;
		30568: Delta = 69'sb000000000000001000000000000000000000000000000000000000001000000000000;
		28485: Delta = 69'sb111111111111111000000000000000000000000000000000000000001000000000000;
		22376: Delta = 69'sb000000000000000111111111111111111111111111111111111111111000000000000;
		20293: Delta = 69'sb111111111111110111111111111111111111111111111111111111111000000000000;
		6179: Delta = 69'sb000000000000010000000000000000000000000000000000000000001000000000000;
		2013: Delta = 69'sb111111111111110000000000000000000000000000000000000000001000000000000;
		48848: Delta = 69'sb000000000000001111111111111111111111111111111111111111111000000000000;
		44682: Delta = 69'sb111111111111101111111111111111111111111111111111111111111000000000000;
		8262: Delta = 69'sb000000000000100000000000000000000000000000000000000000001000000000000;
		50791: Delta = 69'sb111111111111100000000000000000000000000000000000000000001000000000000;
		70: Delta = 69'sb000000000000011111111111111111111111111111111111111111111000000000000;
		42599: Delta = 69'sb111111111111011111111111111111111111111111111111111111111000000000000;
		12428: Delta = 69'sb000000000001000000000000000000000000000000000000000000001000000000000;
		46625: Delta = 69'sb111111111111000000000000000000000000000000000000000000001000000000000;
		4236: Delta = 69'sb000000000000111111111111111111111111111111111111111111111000000000000;
		38433: Delta = 69'sb111111111110111111111111111111111111111111111111111111111000000000000;
		20760: Delta = 69'sb000000000010000000000000000000000000000000000000000000001000000000000;
		38293: Delta = 69'sb111111111110000000000000000000000000000000000000000000001000000000000;
		12568: Delta = 69'sb000000000001111111111111111111111111111111111111111111111000000000000;
		30101: Delta = 69'sb111111111101111111111111111111111111111111111111111111111000000000000;
		37424: Delta = 69'sb000000000100000000000000000000000000000000000000000000001000000000000;
		21629: Delta = 69'sb111111111100000000000000000000000000000000000000000000001000000000000;
		29232: Delta = 69'sb000000000011111111111111111111111111111111111111111111111000000000000;
		13437: Delta = 69'sb111111111011111111111111111111111111111111111111111111111000000000000;
		19891: Delta = 69'sb000000001000000000000000000000000000000000000000000000001000000000000;
		39162: Delta = 69'sb111111111000000000000000000000000000000000000000000000001000000000000;
		11699: Delta = 69'sb000000000111111111111111111111111111111111111111111111111000000000000;
		30970: Delta = 69'sb111111110111111111111111111111111111111111111111111111111000000000000;
		35686: Delta = 69'sb000000010000000000000000000000000000000000000000000000001000000000000;
		23367: Delta = 69'sb111111110000000000000000000000000000000000000000000000001000000000000;
		27494: Delta = 69'sb000000001111111111111111111111111111111111111111111111111000000000000;
		15175: Delta = 69'sb111111101111111111111111111111111111111111111111111111111000000000000;
		16415: Delta = 69'sb000000100000000000000000000000000000000000000000000000001000000000000;
		42638: Delta = 69'sb111111100000000000000000000000000000000000000000000000001000000000000;
		8223: Delta = 69'sb000000011111111111111111111111111111111111111111111111111000000000000;
		34446: Delta = 69'sb111111011111111111111111111111111111111111111111111111111000000000000;
		28734: Delta = 69'sb000001000000000000000000000000000000000000000000000000001000000000000;
		30319: Delta = 69'sb111111000000000000000000000000000000000000000000000000001000000000000;
		20542: Delta = 69'sb000000111111111111111111111111111111111111111111111111111000000000000;
		22127: Delta = 69'sb111110111111111111111111111111111111111111111111111111111000000000000;
		2511: Delta = 69'sb000010000000000000000000000000000000000000000000000000001000000000000;
		5681: Delta = 69'sb111110000000000000000000000000000000000000000000000000001000000000000;
		45180: Delta = 69'sb000001111111111111111111111111111111111111111111111111111000000000000;
		48350: Delta = 69'sb111101111111111111111111111111111111111111111111111111111000000000000;
		926: Delta = 69'sb000100000000000000000000000000000000000000000000000000001000000000000;
		7266: Delta = 69'sb111100000000000000000000000000000000000000000000000000001000000000000;
		43595: Delta = 69'sb000011111111111111111111111111111111111111111111111111111000000000000;
		49935: Delta = 69'sb111011111111111111111111111111111111111111111111111111111000000000000;
		48617: Delta = 69'sb001000000000000000000000000000000000000000000000000000001000000000000;
		10436: Delta = 69'sb111000000000000000000000000000000000000000000000000000001000000000000;
		40425: Delta = 69'sb000111111111111111111111111111111111111111111111111111111000000000000;
		2244: Delta = 69'sb110111111111111111111111111111111111111111111111111111111000000000000;
		42277: Delta = 69'sb010000000000000000000000000000000000000000000000000000001000000000000;
		16776: Delta = 69'sb110000000000000000000000000000000000000000000000000000001000000000000;
		34085: Delta = 69'sb001111111111111111111111111111111111111111111111111111111000000000000;
		8584: Delta = 69'sb101111111111111111111111111111111111111111111111111111111000000000000;
		24576: Delta = 69'sb000000000000000000000000000000000000000000000000000000110000000000000;
		26285: Delta = 69'sb111111111111111111111111111111111111111111111111111111010000000000000;
		40960: Delta = 69'sb000000000000000000000000000000000000000000000000000001010000000000000;
		9901: Delta = 69'sb111111111111111111111111111111111111111111111111111110110000000000000;
		22867: Delta = 69'sb000000000000000000000000000000000000000000000000000010010000000000000;
		44378: Delta = 69'sb111111111111111111111111111111111111111111111111111110010000000000000;
		6483: Delta = 69'sb000000000000000000000000000000000000000000000000000001110000000000000;
		27994: Delta = 69'sb111111111111111111111111111111111111111111111111111101110000000000000;
		37542: Delta = 69'sb000000000000000000000000000000000000000000000000000100010000000000000;
		29703: Delta = 69'sb111111111111111111111111111111111111111111111111111100010000000000000;
		21158: Delta = 69'sb000000000000000000000000000000000000000000000000000011110000000000000;
		13319: Delta = 69'sb111111111111111111111111111111111111111111111111111011110000000000000;
		16031: Delta = 69'sb000000000000000000000000000000000000000000000000001000010000000000000;
		353: Delta = 69'sb111111111111111111111111111111111111111111111111111000010000000000000;
		50508: Delta = 69'sb000000000000000000000000000000000000000000000000000111110000000000000;
		34830: Delta = 69'sb111111111111111111111111111111111111111111111111110111110000000000000;
		23870: Delta = 69'sb000000000000000000000000000000000000000000000000010000010000000000000;
		43375: Delta = 69'sb111111111111111111111111111111111111111111111111110000010000000000000;
		7486: Delta = 69'sb000000000000000000000000000000000000000000000000001111110000000000000;
		26991: Delta = 69'sb111111111111111111111111111111111111111111111111101111110000000000000;
		39548: Delta = 69'sb000000000000000000000000000000000000000000000000100000010000000000000;
		27697: Delta = 69'sb111111111111111111111111111111111111111111111111100000010000000000000;
		23164: Delta = 69'sb000000000000000000000000000000000000000000000000011111110000000000000;
		11313: Delta = 69'sb111111111111111111111111111111111111111111111111011111110000000000000;
		20043: Delta = 69'sb000000000000000000000000000000000000000000000001000000010000000000000;
		47202: Delta = 69'sb111111111111111111111111111111111111111111111111000000010000000000000;
		3659: Delta = 69'sb000000000000000000000000000000000000000000000000111111110000000000000;
		30818: Delta = 69'sb111111111111111111111111111111111111111111111110111111110000000000000;
		31894: Delta = 69'sb000000000000000000000000000000000000000000000010000000010000000000000;
		35351: Delta = 69'sb111111111111111111111111111111111111111111111110000000010000000000000;
		15510: Delta = 69'sb000000000000000000000000000000000000000000000001111111110000000000000;
		18967: Delta = 69'sb111111111111111111111111111111111111111111111101111111110000000000000;
		4735: Delta = 69'sb000000000000000000000000000000000000000000000100000000010000000000000;
		11649: Delta = 69'sb111111111111111111111111111111111111111111111100000000010000000000000;
		39212: Delta = 69'sb000000000000000000000000000000000000000000000011111111110000000000000;
		46126: Delta = 69'sb111111111111111111111111111111111111111111111011111111110000000000000;
		1278: Delta = 69'sb000000000000000000000000000000000000000000001000000000010000000000000;
		15106: Delta = 69'sb111111111111111111111111111111111111111111111000000000010000000000000;
		35755: Delta = 69'sb000000000000000000000000000000000000000000000111111111110000000000000;
		49583: Delta = 69'sb111111111111111111111111111111111111111111110111111111110000000000000;
		45225: Delta = 69'sb000000000000000000000000000000000000000000010000000000010000000000000;
		22020: Delta = 69'sb111111111111111111111111111111111111111111110000000000010000000000000;
		28841: Delta = 69'sb000000000000000000000000000000000000000000001111111111110000000000000;
		5636: Delta = 69'sb111111111111111111111111111111111111111111101111111111110000000000000;
		31397: Delta = 69'sb000000000000000000000000000000000000000000100000000000010000000000000;
		35848: Delta = 69'sb111111111111111111111111111111111111111111100000000000010000000000000;
		15013: Delta = 69'sb000000000000000000000000000000000000000000011111111111110000000000000;
		19464: Delta = 69'sb111111111111111111111111111111111111111111011111111111110000000000000;
		3741: Delta = 69'sb000000000000000000000000000000000000000001000000000000010000000000000;
		12643: Delta = 69'sb111111111111111111111111111111111111111111000000000000010000000000000;
		38218: Delta = 69'sb000000000000000000000000000000000000000000111111111111110000000000000;
		47120: Delta = 69'sb111111111111111111111111111111111111111110111111111111110000000000000;
		50151: Delta = 69'sb000000000000000000000000000000000000000010000000000000010000000000000;
		17094: Delta = 69'sb111111111111111111111111111111111111111110000000000000010000000000000;
		33767: Delta = 69'sb000000000000000000000000000000000000000001111111111111110000000000000;
		710: Delta = 69'sb111111111111111111111111111111111111111101111111111111110000000000000;
		41249: Delta = 69'sb000000000000000000000000000000000000000100000000000000010000000000000;
		25996: Delta = 69'sb111111111111111111111111111111111111111100000000000000010000000000000;
		24865: Delta = 69'sb000000000000000000000000000000000000000011111111111111110000000000000;
		9612: Delta = 69'sb111111111111111111111111111111111111111011111111111111110000000000000;
		23445: Delta = 69'sb000000000000000000000000000000000000001000000000000000010000000000000;
		43800: Delta = 69'sb111111111111111111111111111111111111111000000000000000010000000000000;
		7061: Delta = 69'sb000000000000000000000000000000000000000111111111111111110000000000000;
		27416: Delta = 69'sb111111111111111111111111111111111111110111111111111111110000000000000;
		38698: Delta = 69'sb000000000000000000000000000000000000010000000000000000010000000000000;
		28547: Delta = 69'sb111111111111111111111111111111111111110000000000000000010000000000000;
		22314: Delta = 69'sb000000000000000000000000000000000000001111111111111111110000000000000;
		12163: Delta = 69'sb111111111111111111111111111111111111101111111111111111110000000000000;
		18343: Delta = 69'sb000000000000000000000000000000000000100000000000000000010000000000000;
		48902: Delta = 69'sb111111111111111111111111111111111111100000000000000000010000000000000;
		1959: Delta = 69'sb000000000000000000000000000000000000011111111111111111110000000000000;
		32518: Delta = 69'sb111111111111111111111111111111111111011111111111111111110000000000000;
		28494: Delta = 69'sb000000000000000000000000000000000001000000000000000000010000000000000;
		38751: Delta = 69'sb111111111111111111111111111111111111000000000000000000010000000000000;
		12110: Delta = 69'sb000000000000000000000000000000000000111111111111111111110000000000000;
		22367: Delta = 69'sb111111111111111111111111111111111110111111111111111111110000000000000;
		48796: Delta = 69'sb000000000000000000000000000000000010000000000000000000010000000000000;
		18449: Delta = 69'sb111111111111111111111111111111111110000000000000000000010000000000000;
		32412: Delta = 69'sb000000000000000000000000000000000001111111111111111111110000000000000;
		2065: Delta = 69'sb111111111111111111111111111111111101111111111111111111110000000000000;
		38539: Delta = 69'sb000000000000000000000000000000000100000000000000000000010000000000000;
		28706: Delta = 69'sb111111111111111111111111111111111100000000000000000000010000000000000;
		22155: Delta = 69'sb000000000000000000000000000000000011111111111111111111110000000000000;
		12322: Delta = 69'sb111111111111111111111111111111111011111111111111111111110000000000000;
		18025: Delta = 69'sb000000000000000000000000000000001000000000000000000000010000000000000;
		49220: Delta = 69'sb111111111111111111111111111111111000000000000000000000010000000000000;
		1641: Delta = 69'sb000000000000000000000000000000000111111111111111111111110000000000000;
		32836: Delta = 69'sb111111111111111111111111111111110111111111111111111111110000000000000;
		27858: Delta = 69'sb000000000000000000000000000000010000000000000000000000010000000000000;
		39387: Delta = 69'sb111111111111111111111111111111110000000000000000000000010000000000000;
		11474: Delta = 69'sb000000000000000000000000000000001111111111111111111111110000000000000;
		23003: Delta = 69'sb111111111111111111111111111111101111111111111111111111110000000000000;
		47524: Delta = 69'sb000000000000000000000000000000100000000000000000000000010000000000000;
		19721: Delta = 69'sb111111111111111111111111111111100000000000000000000000010000000000000;
		31140: Delta = 69'sb000000000000000000000000000000011111111111111111111111110000000000000;
		3337: Delta = 69'sb111111111111111111111111111111011111111111111111111111110000000000000;
		35995: Delta = 69'sb000000000000000000000000000001000000000000000000000000010000000000000;
		31250: Delta = 69'sb111111111111111111111111111111000000000000000000000000010000000000000;
		19611: Delta = 69'sb000000000000000000000000000000111111111111111111111111110000000000000;
		14866: Delta = 69'sb111111111111111111111111111110111111111111111111111111110000000000000;
		12937: Delta = 69'sb000000000000000000000000000010000000000000000000000000010000000000000;
		3447: Delta = 69'sb111111111111111111111111111110000000000000000000000000010000000000000;
		47414: Delta = 69'sb000000000000000000000000000001111111111111111111111111110000000000000;
		37924: Delta = 69'sb111111111111111111111111111101111111111111111111111111110000000000000;
		17682: Delta = 69'sb000000000000000000000000000100000000000000000000000000010000000000000;
		49563: Delta = 69'sb111111111111111111111111111100000000000000000000000000010000000000000;
		1298: Delta = 69'sb000000000000000000000000000011111111111111111111111111110000000000000;
		33179: Delta = 69'sb111111111111111111111111111011111111111111111111111111110000000000000;
		27172: Delta = 69'sb000000000000000000000000001000000000000000000000000000010000000000000;
		40073: Delta = 69'sb111111111111111111111111111000000000000000000000000000010000000000000;
		10788: Delta = 69'sb000000000000000000000000000111111111111111111111111111110000000000000;
		23689: Delta = 69'sb111111111111111111111111110111111111111111111111111111110000000000000;
		46152: Delta = 69'sb000000000000000000000000010000000000000000000000000000010000000000000;
		21093: Delta = 69'sb111111111111111111111111110000000000000000000000000000010000000000000;
		29768: Delta = 69'sb000000000000000000000000001111111111111111111111111111110000000000000;
		4709: Delta = 69'sb111111111111111111111111101111111111111111111111111111110000000000000;
		33251: Delta = 69'sb000000000000000000000000100000000000000000000000000000010000000000000;
		33994: Delta = 69'sb111111111111111111111111100000000000000000000000000000010000000000000;
		16867: Delta = 69'sb000000000000000000000000011111111111111111111111111111110000000000000;
		17610: Delta = 69'sb111111111111111111111111011111111111111111111111111111110000000000000;
		7449: Delta = 69'sb000000000000000000000001000000000000000000000000000000010000000000000;
		8935: Delta = 69'sb111111111111111111111111000000000000000000000000000000010000000000000;
		41926: Delta = 69'sb000000000000000000000000111111111111111111111111111111110000000000000;
		43412: Delta = 69'sb111111111111111111111110111111111111111111111111111111110000000000000;
		6706: Delta = 69'sb000000000000000000000010000000000000000000000000000000010000000000000;
		9678: Delta = 69'sb111111111111111111111110000000000000000000000000000000010000000000000;
		41183: Delta = 69'sb000000000000000000000001111111111111111111111111111111110000000000000;
		44155: Delta = 69'sb111111111111111111111101111111111111111111111111111111110000000000000;
		5220: Delta = 69'sb000000000000000000000100000000000000000000000000000000010000000000000;
		11164: Delta = 69'sb111111111111111111111100000000000000000000000000000000010000000000000;
		39697: Delta = 69'sb000000000000000000000011111111111111111111111111111111110000000000000;
		45641: Delta = 69'sb111111111111111111111011111111111111111111111111111111110000000000000;
		2248: Delta = 69'sb000000000000000000001000000000000000000000000000000000010000000000000;
		14136: Delta = 69'sb111111111111111111111000000000000000000000000000000000010000000000000;
		36725: Delta = 69'sb000000000000000000000111111111111111111111111111111111110000000000000;
		48613: Delta = 69'sb111111111111111111110111111111111111111111111111111111110000000000000;
		47165: Delta = 69'sb000000000000000000010000000000000000000000000000000000010000000000000;
		20080: Delta = 69'sb111111111111111111110000000000000000000000000000000000010000000000000;
		30781: Delta = 69'sb000000000000000000001111111111111111111111111111111111110000000000000;
		3696: Delta = 69'sb111111111111111111101111111111111111111111111111111111110000000000000;
		35277: Delta = 69'sb000000000000000000100000000000000000000000000000000000010000000000000;
		31968: Delta = 69'sb111111111111111111100000000000000000000000000000000000010000000000000;
		18893: Delta = 69'sb000000000000000000011111111111111111111111111111111111110000000000000;
		15584: Delta = 69'sb111111111111111111011111111111111111111111111111111111110000000000000;
		11501: Delta = 69'sb000000000000000001000000000000000000000000000000000000010000000000000;
		4883: Delta = 69'sb111111111111111111000000000000000000000000000000000000010000000000000;
		45978: Delta = 69'sb000000000000000000111111111111111111111111111111111111110000000000000;
		39360: Delta = 69'sb111111111111111110111111111111111111111111111111111111110000000000000;
		14810: Delta = 69'sb000000000000000010000000000000000000000000000000000000010000000000000;
		1574: Delta = 69'sb111111111111111110000000000000000000000000000000000000010000000000000;
		49287: Delta = 69'sb000000000000000001111111111111111111111111111111111111110000000000000;
		36051: Delta = 69'sb111111111111111101111111111111111111111111111111111111110000000000000;
		21428: Delta = 69'sb000000000000000100000000000000000000000000000000000000010000000000000;
		45817: Delta = 69'sb111111111111111100000000000000000000000000000000000000010000000000000;
		5044: Delta = 69'sb000000000000000011111111111111111111111111111111111111110000000000000;
		29433: Delta = 69'sb111111111111111011111111111111111111111111111111111111110000000000000;
		34664: Delta = 69'sb000000000000001000000000000000000000000000000000000000010000000000000;
		32581: Delta = 69'sb111111111111111000000000000000000000000000000000000000010000000000000;
		18280: Delta = 69'sb000000000000000111111111111111111111111111111111111111110000000000000;
		16197: Delta = 69'sb111111111111110111111111111111111111111111111111111111110000000000000;
		10275: Delta = 69'sb000000000000010000000000000000000000000000000000000000010000000000000;
		6109: Delta = 69'sb111111111111110000000000000000000000000000000000000000010000000000000;
		44752: Delta = 69'sb000000000000001111111111111111111111111111111111111111110000000000000;
		40586: Delta = 69'sb111111111111101111111111111111111111111111111111111111110000000000000;
		12358: Delta = 69'sb000000000000100000000000000000000000000000000000000000010000000000000;
		4026: Delta = 69'sb111111111111100000000000000000000000000000000000000000010000000000000;
		46835: Delta = 69'sb000000000000011111111111111111111111111111111111111111110000000000000;
		38503: Delta = 69'sb111111111111011111111111111111111111111111111111111111110000000000000;
		16524: Delta = 69'sb000000000001000000000000000000000000000000000000000000010000000000000;
		50721: Delta = 69'sb111111111111000000000000000000000000000000000000000000010000000000000;
		140: Delta = 69'sb000000000000111111111111111111111111111111111111111111110000000000000;
		34337: Delta = 69'sb111111111110111111111111111111111111111111111111111111110000000000000;
		24856: Delta = 69'sb000000000010000000000000000000000000000000000000000000010000000000000;
		42389: Delta = 69'sb111111111110000000000000000000000000000000000000000000010000000000000;
		8472: Delta = 69'sb000000000001111111111111111111111111111111111111111111110000000000000;
		26005: Delta = 69'sb111111111101111111111111111111111111111111111111111111110000000000000;
		41520: Delta = 69'sb000000000100000000000000000000000000000000000000000000010000000000000;
		25725: Delta = 69'sb111111111100000000000000000000000000000000000000000000010000000000000;
		25136: Delta = 69'sb000000000011111111111111111111111111111111111111111111110000000000000;
		9341: Delta = 69'sb111111111011111111111111111111111111111111111111111111110000000000000;
		23987: Delta = 69'sb000000001000000000000000000000000000000000000000000000010000000000000;
		43258: Delta = 69'sb111111111000000000000000000000000000000000000000000000010000000000000;
		7603: Delta = 69'sb000000000111111111111111111111111111111111111111111111110000000000000;
		26874: Delta = 69'sb111111110111111111111111111111111111111111111111111111110000000000000;
		39782: Delta = 69'sb000000010000000000000000000000000000000000000000000000010000000000000;
		27463: Delta = 69'sb111111110000000000000000000000000000000000000000000000010000000000000;
		23398: Delta = 69'sb000000001111111111111111111111111111111111111111111111110000000000000;
		11079: Delta = 69'sb111111101111111111111111111111111111111111111111111111110000000000000;
		20511: Delta = 69'sb000000100000000000000000000000000000000000000000000000010000000000000;
		46734: Delta = 69'sb111111100000000000000000000000000000000000000000000000010000000000000;
		4127: Delta = 69'sb000000011111111111111111111111111111111111111111111111110000000000000;
		30350: Delta = 69'sb111111011111111111111111111111111111111111111111111111110000000000000;
		32830: Delta = 69'sb000001000000000000000000000000000000000000000000000000010000000000000;
		34415: Delta = 69'sb111111000000000000000000000000000000000000000000000000010000000000000;
		16446: Delta = 69'sb000000111111111111111111111111111111111111111111111111110000000000000;
		18031: Delta = 69'sb111110111111111111111111111111111111111111111111111111110000000000000;
		6607: Delta = 69'sb000010000000000000000000000000000000000000000000000000010000000000000;
		9777: Delta = 69'sb111110000000000000000000000000000000000000000000000000010000000000000;
		41084: Delta = 69'sb000001111111111111111111111111111111111111111111111111110000000000000;
		44254: Delta = 69'sb111101111111111111111111111111111111111111111111111111110000000000000;
		5022: Delta = 69'sb000100000000000000000000000000000000000000000000000000010000000000000;
		11362: Delta = 69'sb111100000000000000000000000000000000000000000000000000010000000000000;
		39499: Delta = 69'sb000011111111111111111111111111111111111111111111111111110000000000000;
		45839: Delta = 69'sb111011111111111111111111111111111111111111111111111111110000000000000;
		1852: Delta = 69'sb001000000000000000000000000000000000000000000000000000010000000000000;
		14532: Delta = 69'sb111000000000000000000000000000000000000000000000000000010000000000000;
		36329: Delta = 69'sb000111111111111111111111111111111111111111111111111111110000000000000;
		49009: Delta = 69'sb110111111111111111111111111111111111111111111111111111110000000000000;
		46373: Delta = 69'sb010000000000000000000000000000000000000000000000000000010000000000000;
		20872: Delta = 69'sb110000000000000000000000000000000000000000000000000000010000000000000;
		29989: Delta = 69'sb001111111111111111111111111111111111111111111111111111110000000000000;
		4488: Delta = 69'sb101111111111111111111111111111111111111111111111111111110000000000000;
		49152: Delta = 69'sb000000000000000000000000000000000000000000000000000001100000000000000;
		1709: Delta = 69'sb111111111111111111111111111111111111111111111111111110100000000000000;
		31059: Delta = 69'sb000000000000000000000000000000000000000000000000000010100000000000000;
		19802: Delta = 69'sb111111111111111111111111111111111111111111111111111101100000000000000;
		45734: Delta = 69'sb000000000000000000000000000000000000000000000000000100100000000000000;
		37895: Delta = 69'sb111111111111111111111111111111111111111111111111111100100000000000000;
		12966: Delta = 69'sb000000000000000000000000000000000000000000000000000011100000000000000;
		5127: Delta = 69'sb111111111111111111111111111111111111111111111111111011100000000000000;
		24223: Delta = 69'sb000000000000000000000000000000000000000000000000001000100000000000000;
		8545: Delta = 69'sb111111111111111111111111111111111111111111111111111000100000000000000;
		42316: Delta = 69'sb000000000000000000000000000000000000000000000000000111100000000000000;
		26638: Delta = 69'sb111111111111111111111111111111111111111111111111110111100000000000000;
		32062: Delta = 69'sb000000000000000000000000000000000000000000000000010000100000000000000;
		706: Delta = 69'sb111111111111111111111111111111111111111111111111110000100000000000000;
		50155: Delta = 69'sb000000000000000000000000000000000000000000000000001111100000000000000;
		18799: Delta = 69'sb111111111111111111111111111111111111111111111111101111100000000000000;
		47740: Delta = 69'sb000000000000000000000000000000000000000000000000100000100000000000000;
		35889: Delta = 69'sb111111111111111111111111111111111111111111111111100000100000000000000;
		14972: Delta = 69'sb000000000000000000000000000000000000000000000000011111100000000000000;
		3121: Delta = 69'sb111111111111111111111111111111111111111111111111011111100000000000000;
		28235: Delta = 69'sb000000000000000000000000000000000000000000000001000000100000000000000;
		4533: Delta = 69'sb111111111111111111111111111111111111111111111111000000100000000000000;
		46328: Delta = 69'sb000000000000000000000000000000000000000000000000111111100000000000000;
		22626: Delta = 69'sb111111111111111111111111111111111111111111111110111111100000000000000;
		40086: Delta = 69'sb000000000000000000000000000000000000000000000010000000100000000000000;
		43543: Delta = 69'sb111111111111111111111111111111111111111111111110000000100000000000000;
		7318: Delta = 69'sb000000000000000000000000000000000000000000000001111111100000000000000;
		10775: Delta = 69'sb111111111111111111111111111111111111111111111101111111100000000000000;
		12927: Delta = 69'sb000000000000000000000000000000000000000000000100000000100000000000000;
		19841: Delta = 69'sb111111111111111111111111111111111111111111111100000000100000000000000;
		31020: Delta = 69'sb000000000000000000000000000000000000000000000011111111100000000000000;
		37934: Delta = 69'sb111111111111111111111111111111111111111111111011111111100000000000000;
		9470: Delta = 69'sb000000000000000000000000000000000000000000001000000000100000000000000;
		23298: Delta = 69'sb111111111111111111111111111111111111111111111000000000100000000000000;
		27563: Delta = 69'sb000000000000000000000000000000000000000000000111111111100000000000000;
		41391: Delta = 69'sb111111111111111111111111111111111111111111110111111111100000000000000;
		2556: Delta = 69'sb000000000000000000000000000000000000000000010000000000100000000000000;
		30212: Delta = 69'sb111111111111111111111111111111111111111111110000000000100000000000000;
		20649: Delta = 69'sb000000000000000000000000000000000000000000001111111111100000000000000;
		48305: Delta = 69'sb111111111111111111111111111111111111111111101111111111100000000000000;
		39589: Delta = 69'sb000000000000000000000000000000000000000000100000000000100000000000000;
		44040: Delta = 69'sb111111111111111111111111111111111111111111100000000000100000000000000;
		6821: Delta = 69'sb000000000000000000000000000000000000000000011111111111100000000000000;
		11272: Delta = 69'sb111111111111111111111111111111111111111111011111111111100000000000000;
		11933: Delta = 69'sb000000000000000000000000000000000000000001000000000000100000000000000;
		20835: Delta = 69'sb111111111111111111111111111111111111111111000000000000100000000000000;
		30026: Delta = 69'sb000000000000000000000000000000000000000000111111111111100000000000000;
		38928: Delta = 69'sb111111111111111111111111111111111111111110111111111111100000000000000;
		7482: Delta = 69'sb000000000000000000000000000000000000000010000000000000100000000000000;
		25286: Delta = 69'sb111111111111111111111111111111111111111110000000000000100000000000000;
		25575: Delta = 69'sb000000000000000000000000000000000000000001111111111111100000000000000;
		43379: Delta = 69'sb111111111111111111111111111111111111111101111111111111100000000000000;
		49441: Delta = 69'sb000000000000000000000000000000000000000100000000000000100000000000000;
		34188: Delta = 69'sb111111111111111111111111111111111111111100000000000000100000000000000;
		16673: Delta = 69'sb000000000000000000000000000000000000000011111111111111100000000000000;
		1420: Delta = 69'sb111111111111111111111111111111111111111011111111111111100000000000000;
		31637: Delta = 69'sb000000000000000000000000000000000000001000000000000000100000000000000;
		1131: Delta = 69'sb111111111111111111111111111111111111111000000000000000100000000000000;
		49730: Delta = 69'sb000000000000000000000000000000000000000111111111111111100000000000000;
		19224: Delta = 69'sb111111111111111111111111111111111111110111111111111111100000000000000;
		46890: Delta = 69'sb000000000000000000000000000000000000010000000000000000100000000000000;
		36739: Delta = 69'sb111111111111111111111111111111111111110000000000000000100000000000000;
		14122: Delta = 69'sb000000000000000000000000000000000000001111111111111111100000000000000;
		3971: Delta = 69'sb111111111111111111111111111111111111101111111111111111100000000000000;
		26535: Delta = 69'sb000000000000000000000000000000000000100000000000000000100000000000000;
		6233: Delta = 69'sb111111111111111111111111111111111111100000000000000000100000000000000;
		44628: Delta = 69'sb000000000000000000000000000000000000011111111111111111100000000000000;
		24326: Delta = 69'sb111111111111111111111111111111111111011111111111111111100000000000000;
		36686: Delta = 69'sb000000000000000000000000000000000001000000000000000000100000000000000;
		46943: Delta = 69'sb111111111111111111111111111111111111000000000000000000100000000000000;
		3918: Delta = 69'sb000000000000000000000000000000000000111111111111111111100000000000000;
		14175: Delta = 69'sb111111111111111111111111111111111110111111111111111111100000000000000;
		6127: Delta = 69'sb000000000000000000000000000000000010000000000000000000100000000000000;
		26641: Delta = 69'sb111111111111111111111111111111111110000000000000000000100000000000000;
		24220: Delta = 69'sb000000000000000000000000000000000001111111111111111111100000000000000;
		44734: Delta = 69'sb111111111111111111111111111111111101111111111111111111100000000000000;
		46731: Delta = 69'sb000000000000000000000000000000000100000000000000000000100000000000000;
		36898: Delta = 69'sb111111111111111111111111111111111100000000000000000000100000000000000;
		13963: Delta = 69'sb000000000000000000000000000000000011111111111111111111100000000000000;
		4130: Delta = 69'sb111111111111111111111111111111111011111111111111111111100000000000000;
		26217: Delta = 69'sb000000000000000000000000000000001000000000000000000000100000000000000;
		6551: Delta = 69'sb111111111111111111111111111111111000000000000000000000100000000000000;
		44310: Delta = 69'sb000000000000000000000000000000000111111111111111111111100000000000000;
		24644: Delta = 69'sb111111111111111111111111111111110111111111111111111111100000000000000;
		36050: Delta = 69'sb000000000000000000000000000000010000000000000000000000100000000000000;
		47579: Delta = 69'sb111111111111111111111111111111110000000000000000000000100000000000000;
		3282: Delta = 69'sb000000000000000000000000000000001111111111111111111111100000000000000;
		14811: Delta = 69'sb111111111111111111111111111111101111111111111111111111100000000000000;
		4855: Delta = 69'sb000000000000000000000000000000100000000000000000000000100000000000000;
		27913: Delta = 69'sb111111111111111111111111111111100000000000000000000000100000000000000;
		22948: Delta = 69'sb000000000000000000000000000000011111111111111111111111100000000000000;
		46006: Delta = 69'sb111111111111111111111111111111011111111111111111111111100000000000000;
		44187: Delta = 69'sb000000000000000000000000000001000000000000000000000000100000000000000;
		39442: Delta = 69'sb111111111111111111111111111111000000000000000000000000100000000000000;
		11419: Delta = 69'sb000000000000000000000000000000111111111111111111111111100000000000000;
		6674: Delta = 69'sb111111111111111111111111111110111111111111111111111111100000000000000;
		21129: Delta = 69'sb000000000000000000000000000010000000000000000000000000100000000000000;
		11639: Delta = 69'sb111111111111111111111111111110000000000000000000000000100000000000000;
		39222: Delta = 69'sb000000000000000000000000000001111111111111111111111111100000000000000;
		29732: Delta = 69'sb111111111111111111111111111101111111111111111111111111100000000000000;
		25874: Delta = 69'sb000000000000000000000000000100000000000000000000000000100000000000000;
		6894: Delta = 69'sb111111111111111111111111111100000000000000000000000000100000000000000;
		43967: Delta = 69'sb000000000000000000000000000011111111111111111111111111100000000000000;
		24987: Delta = 69'sb111111111111111111111111111011111111111111111111111111100000000000000;
		35364: Delta = 69'sb000000000000000000000000001000000000000000000000000000100000000000000;
		48265: Delta = 69'sb111111111111111111111111111000000000000000000000000000100000000000000;
		2596: Delta = 69'sb000000000000000000000000000111111111111111111111111111100000000000000;
		15497: Delta = 69'sb111111111111111111111111110111111111111111111111111111100000000000000;
		3483: Delta = 69'sb000000000000000000000000010000000000000000000000000000100000000000000;
		29285: Delta = 69'sb111111111111111111111111110000000000000000000000000000100000000000000;
		21576: Delta = 69'sb000000000000000000000000001111111111111111111111111111100000000000000;
		47378: Delta = 69'sb111111111111111111111111101111111111111111111111111111100000000000000;
		41443: Delta = 69'sb000000000000000000000000100000000000000000000000000000100000000000000;
		42186: Delta = 69'sb111111111111111111111111100000000000000000000000000000100000000000000;
		8675: Delta = 69'sb000000000000000000000000011111111111111111111111111111100000000000000;
		9418: Delta = 69'sb111111111111111111111111011111111111111111111111111111100000000000000;
		15641: Delta = 69'sb000000000000000000000001000000000000000000000000000000100000000000000;
		17127: Delta = 69'sb111111111111111111111111000000000000000000000000000000100000000000000;
		33734: Delta = 69'sb000000000000000000000000111111111111111111111111111111100000000000000;
		35220: Delta = 69'sb111111111111111111111110111111111111111111111111111111100000000000000;
		14898: Delta = 69'sb000000000000000000000010000000000000000000000000000000100000000000000;
		17870: Delta = 69'sb111111111111111111111110000000000000000000000000000000100000000000000;
		32991: Delta = 69'sb000000000000000000000001111111111111111111111111111111100000000000000;
		35963: Delta = 69'sb111111111111111111111101111111111111111111111111111111100000000000000;
		13412: Delta = 69'sb000000000000000000000100000000000000000000000000000000100000000000000;
		19356: Delta = 69'sb111111111111111111111100000000000000000000000000000000100000000000000;
		31505: Delta = 69'sb000000000000000000000011111111111111111111111111111111100000000000000;
		37449: Delta = 69'sb111111111111111111111011111111111111111111111111111111100000000000000;
		10440: Delta = 69'sb000000000000000000001000000000000000000000000000000000100000000000000;
		22328: Delta = 69'sb111111111111111111111000000000000000000000000000000000100000000000000;
		28533: Delta = 69'sb000000000000000000000111111111111111111111111111111111100000000000000;
		40421: Delta = 69'sb111111111111111111110111111111111111111111111111111111100000000000000;
		4496: Delta = 69'sb000000000000000000010000000000000000000000000000000000100000000000000;
		28272: Delta = 69'sb111111111111111111110000000000000000000000000000000000100000000000000;
		22589: Delta = 69'sb000000000000000000001111111111111111111111111111111111100000000000000;
		46365: Delta = 69'sb111111111111111111101111111111111111111111111111111111100000000000000;
		43469: Delta = 69'sb000000000000000000100000000000000000000000000000000000100000000000000;
		40160: Delta = 69'sb111111111111111111100000000000000000000000000000000000100000000000000;
		10701: Delta = 69'sb000000000000000000011111111111111111111111111111111111100000000000000;
		7392: Delta = 69'sb111111111111111111011111111111111111111111111111111111100000000000000;
		19693: Delta = 69'sb000000000000000001000000000000000000000000000000000000100000000000000;
		13075: Delta = 69'sb111111111111111111000000000000000000000000000000000000100000000000000;
		37786: Delta = 69'sb000000000000000000111111111111111111111111111111111111100000000000000;
		31168: Delta = 69'sb111111111111111110111111111111111111111111111111111111100000000000000;
		23002: Delta = 69'sb000000000000000010000000000000000000000000000000000000100000000000000;
		9766: Delta = 69'sb111111111111111110000000000000000000000000000000000000100000000000000;
		41095: Delta = 69'sb000000000000000001111111111111111111111111111111111111100000000000000;
		27859: Delta = 69'sb111111111111111101111111111111111111111111111111111111100000000000000;
		29620: Delta = 69'sb000000000000000100000000000000000000000000000000000000100000000000000;
		3148: Delta = 69'sb111111111111111100000000000000000000000000000000000000100000000000000;
		47713: Delta = 69'sb000000000000000011111111111111111111111111111111111111100000000000000;
		21241: Delta = 69'sb111111111111111011111111111111111111111111111111111111100000000000000;
		42856: Delta = 69'sb000000000000001000000000000000000000000000000000000000100000000000000;
		40773: Delta = 69'sb111111111111111000000000000000000000000000000000000000100000000000000;
		10088: Delta = 69'sb000000000000000111111111111111111111111111111111111111100000000000000;
		8005: Delta = 69'sb111111111111110111111111111111111111111111111111111111100000000000000;
		18467: Delta = 69'sb000000000000010000000000000000000000000000000000000000100000000000000;
		14301: Delta = 69'sb111111111111110000000000000000000000000000000000000000100000000000000;
		36560: Delta = 69'sb000000000000001111111111111111111111111111111111111111100000000000000;
		32394: Delta = 69'sb111111111111101111111111111111111111111111111111111111100000000000000;
		20550: Delta = 69'sb000000000000100000000000000000000000000000000000000000100000000000000;
		12218: Delta = 69'sb111111111111100000000000000000000000000000000000000000100000000000000;
		38643: Delta = 69'sb000000000000011111111111111111111111111111111111111111100000000000000;
		30311: Delta = 69'sb111111111111011111111111111111111111111111111111111111100000000000000;
		24716: Delta = 69'sb000000000001000000000000000000000000000000000000000000100000000000000;
		8052: Delta = 69'sb111111111111000000000000000000000000000000000000000000100000000000000;
		42809: Delta = 69'sb000000000000111111111111111111111111111111111111111111100000000000000;
		26145: Delta = 69'sb111111111110111111111111111111111111111111111111111111100000000000000;
		33048: Delta = 69'sb000000000010000000000000000000000000000000000000000000100000000000000;
		50581: Delta = 69'sb111111111110000000000000000000000000000000000000000000100000000000000;
		280: Delta = 69'sb000000000001111111111111111111111111111111111111111111100000000000000;
		17813: Delta = 69'sb111111111101111111111111111111111111111111111111111111100000000000000;
		49712: Delta = 69'sb000000000100000000000000000000000000000000000000000000100000000000000;
		33917: Delta = 69'sb111111111100000000000000000000000000000000000000000000100000000000000;
		16944: Delta = 69'sb000000000011111111111111111111111111111111111111111111100000000000000;
		1149: Delta = 69'sb111111111011111111111111111111111111111111111111111111100000000000000;
		32179: Delta = 69'sb000000001000000000000000000000000000000000000000000000100000000000000;
		589: Delta = 69'sb111111111000000000000000000000000000000000000000000000100000000000000;
		50272: Delta = 69'sb000000000111111111111111111111111111111111111111111111100000000000000;
		18682: Delta = 69'sb111111110111111111111111111111111111111111111111111111100000000000000;
		47974: Delta = 69'sb000000010000000000000000000000000000000000000000000000100000000000000;
		35655: Delta = 69'sb111111110000000000000000000000000000000000000000000000100000000000000;
		15206: Delta = 69'sb000000001111111111111111111111111111111111111111111111100000000000000;
		2887: Delta = 69'sb111111101111111111111111111111111111111111111111111111100000000000000;
		28703: Delta = 69'sb000000100000000000000000000000000000000000000000000000100000000000000;
		4065: Delta = 69'sb111111100000000000000000000000000000000000000000000000100000000000000;
		46796: Delta = 69'sb000000011111111111111111111111111111111111111111111111100000000000000;
		22158: Delta = 69'sb111111011111111111111111111111111111111111111111111111100000000000000;
		41022: Delta = 69'sb000001000000000000000000000000000000000000000000000000100000000000000;
		42607: Delta = 69'sb111111000000000000000000000000000000000000000000000000100000000000000;
		8254: Delta = 69'sb000000111111111111111111111111111111111111111111111111100000000000000;
		9839: Delta = 69'sb111110111111111111111111111111111111111111111111111111100000000000000;
		14799: Delta = 69'sb000010000000000000000000000000000000000000000000000000100000000000000;
		17969: Delta = 69'sb111110000000000000000000000000000000000000000000000000100000000000000;
		32892: Delta = 69'sb000001111111111111111111111111111111111111111111111111100000000000000;
		36062: Delta = 69'sb111101111111111111111111111111111111111111111111111111100000000000000;
		13214: Delta = 69'sb000100000000000000000000000000000000000000000000000000100000000000000;
		19554: Delta = 69'sb111100000000000000000000000000000000000000000000000000100000000000000;
		31307: Delta = 69'sb000011111111111111111111111111111111111111111111111111100000000000000;
		37647: Delta = 69'sb111011111111111111111111111111111111111111111111111111100000000000000;
		10044: Delta = 69'sb001000000000000000000000000000000000000000000000000000100000000000000;
		22724: Delta = 69'sb111000000000000000000000000000000000000000000000000000100000000000000;
		28137: Delta = 69'sb000111111111111111111111111111111111111111111111111111100000000000000;
		40817: Delta = 69'sb110111111111111111111111111111111111111111111111111111100000000000000;
		3704: Delta = 69'sb010000000000000000000000000000000000000000000000000000100000000000000;
		29064: Delta = 69'sb110000000000000000000000000000000000000000000000000000100000000000000;
		21797: Delta = 69'sb001111111111111111111111111111111111111111111111111111100000000000000;
		47157: Delta = 69'sb101111111111111111111111111111111111111111111111111111100000000000000;
		47443: Delta = 69'sb000000000000000000000000000000000000000000000000000011000000000000000;
		3418: Delta = 69'sb111111111111111111111111111111111111111111111111111101000000000000000;
		11257: Delta = 69'sb000000000000000000000000000000000000000000000000000101000000000000000;
		39604: Delta = 69'sb111111111111111111111111111111111111111111111111111011000000000000000;
		40607: Delta = 69'sb000000000000000000000000000000000000000000000000001001000000000000000;
		24929: Delta = 69'sb111111111111111111111111111111111111111111111111111001000000000000000;
		25932: Delta = 69'sb000000000000000000000000000000000000000000000000000111000000000000000;
		10254: Delta = 69'sb111111111111111111111111111111111111111111111111110111000000000000000;
		48446: Delta = 69'sb000000000000000000000000000000000000000000000000010001000000000000000;
		17090: Delta = 69'sb111111111111111111111111111111111111111111111111110001000000000000000;
		33771: Delta = 69'sb000000000000000000000000000000000000000000000000001111000000000000000;
		2415: Delta = 69'sb111111111111111111111111111111111111111111111111101111000000000000000;
		13263: Delta = 69'sb000000000000000000000000000000000000000000000000100001000000000000000;
		1412: Delta = 69'sb111111111111111111111111111111111111111111111111100001000000000000000;
		49449: Delta = 69'sb000000000000000000000000000000000000000000000000011111000000000000000;
		37598: Delta = 69'sb111111111111111111111111111111111111111111111111011111000000000000000;
		44619: Delta = 69'sb000000000000000000000000000000000000000000000001000001000000000000000;
		20917: Delta = 69'sb111111111111111111111111111111111111111111111111000001000000000000000;
		29944: Delta = 69'sb000000000000000000000000000000000000000000000000111111000000000000000;
		6242: Delta = 69'sb111111111111111111111111111111111111111111111110111111000000000000000;
		5609: Delta = 69'sb000000000000000000000000000000000000000000000010000001000000000000000;
		9066: Delta = 69'sb111111111111111111111111111111111111111111111110000001000000000000000;
		41795: Delta = 69'sb000000000000000000000000000000000000000000000001111111000000000000000;
		45252: Delta = 69'sb111111111111111111111111111111111111111111111101111111000000000000000;
		29311: Delta = 69'sb000000000000000000000000000000000000000000000100000001000000000000000;
		36225: Delta = 69'sb111111111111111111111111111111111111111111111100000001000000000000000;
		14636: Delta = 69'sb000000000000000000000000000000000000000000000011111111000000000000000;
		21550: Delta = 69'sb111111111111111111111111111111111111111111111011111111000000000000000;
		25854: Delta = 69'sb000000000000000000000000000000000000000000001000000001000000000000000;
		39682: Delta = 69'sb111111111111111111111111111111111111111111111000000001000000000000000;
		11179: Delta = 69'sb000000000000000000000000000000000000000000000111111111000000000000000;
		25007: Delta = 69'sb111111111111111111111111111111111111111111110111111111000000000000000;
		18940: Delta = 69'sb000000000000000000000000000000000000000000010000000001000000000000000;
		46596: Delta = 69'sb111111111111111111111111111111111111111111110000000001000000000000000;
		4265: Delta = 69'sb000000000000000000000000000000000000000000001111111111000000000000000;
		31921: Delta = 69'sb111111111111111111111111111111111111111111101111111111000000000000000;
		5112: Delta = 69'sb000000000000000000000000000000000000000000100000000001000000000000000;
		9563: Delta = 69'sb111111111111111111111111111111111111111111100000000001000000000000000;
		41298: Delta = 69'sb000000000000000000000000000000000000000000011111111111000000000000000;
		45749: Delta = 69'sb111111111111111111111111111111111111111111011111111111000000000000000;
		28317: Delta = 69'sb000000000000000000000000000000000000000001000000000001000000000000000;
		37219: Delta = 69'sb111111111111111111111111111111111111111111000000000001000000000000000;
		13642: Delta = 69'sb000000000000000000000000000000000000000000111111111111000000000000000;
		22544: Delta = 69'sb111111111111111111111111111111111111111110111111111111000000000000000;
		23866: Delta = 69'sb000000000000000000000000000000000000000010000000000001000000000000000;
		41670: Delta = 69'sb111111111111111111111111111111111111111110000000000001000000000000000;
		9191: Delta = 69'sb000000000000000000000000000000000000000001111111111111000000000000000;
		26995: Delta = 69'sb111111111111111111111111111111111111111101111111111111000000000000000;
		14964: Delta = 69'sb000000000000000000000000000000000000000100000000000001000000000000000;
		50572: Delta = 69'sb111111111111111111111111111111111111111100000000000001000000000000000;
		289: Delta = 69'sb000000000000000000000000000000000000000011111111111111000000000000000;
		35897: Delta = 69'sb111111111111111111111111111111111111111011111111111111000000000000000;
		48021: Delta = 69'sb000000000000000000000000000000000000001000000000000001000000000000000;
		17515: Delta = 69'sb111111111111111111111111111111111111111000000000000001000000000000000;
		33346: Delta = 69'sb000000000000000000000000000000000000000111111111111111000000000000000;
		2840: Delta = 69'sb111111111111111111111111111111111111110111111111111111000000000000000;
		12413: Delta = 69'sb000000000000000000000000000000000000010000000000000001000000000000000;
		2262: Delta = 69'sb111111111111111111111111111111111111110000000000000001000000000000000;
		48599: Delta = 69'sb000000000000000000000000000000000000001111111111111111000000000000000;
		38448: Delta = 69'sb111111111111111111111111111111111111101111111111111111000000000000000;
		42919: Delta = 69'sb000000000000000000000000000000000000100000000000000001000000000000000;
		22617: Delta = 69'sb111111111111111111111111111111111111100000000000000001000000000000000;
		28244: Delta = 69'sb000000000000000000000000000000000000011111111111111111000000000000000;
		7942: Delta = 69'sb111111111111111111111111111111111111011111111111111111000000000000000;
		2209: Delta = 69'sb000000000000000000000000000000000001000000000000000001000000000000000;
		12466: Delta = 69'sb111111111111111111111111111111111111000000000000000001000000000000000;
		38395: Delta = 69'sb000000000000000000000000000000000000111111111111111111000000000000000;
		48652: Delta = 69'sb111111111111111111111111111111111110111111111111111111000000000000000;
		22511: Delta = 69'sb000000000000000000000000000000000010000000000000000001000000000000000;
		43025: Delta = 69'sb111111111111111111111111111111111110000000000000000001000000000000000;
		7836: Delta = 69'sb000000000000000000000000000000000001111111111111111111000000000000000;
		28350: Delta = 69'sb111111111111111111111111111111111101111111111111111111000000000000000;
		12254: Delta = 69'sb000000000000000000000000000000000100000000000000000001000000000000000;
		2421: Delta = 69'sb111111111111111111111111111111111100000000000000000001000000000000000;
		48440: Delta = 69'sb000000000000000000000000000000000011111111111111111111000000000000000;
		38607: Delta = 69'sb111111111111111111111111111111111011111111111111111111000000000000000;
		42601: Delta = 69'sb000000000000000000000000000000001000000000000000000001000000000000000;
		22935: Delta = 69'sb111111111111111111111111111111111000000000000000000001000000000000000;
		27926: Delta = 69'sb000000000000000000000000000000000111111111111111111111000000000000000;
		8260: Delta = 69'sb111111111111111111111111111111110111111111111111111111000000000000000;
		1573: Delta = 69'sb000000000000000000000000000000010000000000000000000001000000000000000;
		13102: Delta = 69'sb111111111111111111111111111111110000000000000000000001000000000000000;
		37759: Delta = 69'sb000000000000000000000000000000001111111111111111111111000000000000000;
		49288: Delta = 69'sb111111111111111111111111111111101111111111111111111111000000000000000;
		21239: Delta = 69'sb000000000000000000000000000000100000000000000000000001000000000000000;
		44297: Delta = 69'sb111111111111111111111111111111100000000000000000000001000000000000000;
		6564: Delta = 69'sb000000000000000000000000000000011111111111111111111111000000000000000;
		29622: Delta = 69'sb111111111111111111111111111111011111111111111111111111000000000000000;
		9710: Delta = 69'sb000000000000000000000000000001000000000000000000000001000000000000000;
		4965: Delta = 69'sb111111111111111111111111111111000000000000000000000001000000000000000;
		45896: Delta = 69'sb000000000000000000000000000000111111111111111111111111000000000000000;
		41151: Delta = 69'sb111111111111111111111111111110111111111111111111111111000000000000000;
		37513: Delta = 69'sb000000000000000000000000000010000000000000000000000001000000000000000;
		28023: Delta = 69'sb111111111111111111111111111110000000000000000000000001000000000000000;
		22838: Delta = 69'sb000000000000000000000000000001111111111111111111111111000000000000000;
		13348: Delta = 69'sb111111111111111111111111111101111111111111111111111111000000000000000;
		42258: Delta = 69'sb000000000000000000000000000100000000000000000000000001000000000000000;
		23278: Delta = 69'sb111111111111111111111111111100000000000000000000000001000000000000000;
		27583: Delta = 69'sb000000000000000000000000000011111111111111111111111111000000000000000;
		8603: Delta = 69'sb111111111111111111111111111011111111111111111111111111000000000000000;
		887: Delta = 69'sb000000000000000000000000001000000000000000000000000001000000000000000;
		13788: Delta = 69'sb111111111111111111111111111000000000000000000000000001000000000000000;
		37073: Delta = 69'sb000000000000000000000000000111111111111111111111111111000000000000000;
		49974: Delta = 69'sb111111111111111111111111110111111111111111111111111111000000000000000;
		19867: Delta = 69'sb000000000000000000000000010000000000000000000000000001000000000000000;
		45669: Delta = 69'sb111111111111111111111111110000000000000000000000000001000000000000000;
		5192: Delta = 69'sb000000000000000000000000001111111111111111111111111111000000000000000;
		30994: Delta = 69'sb111111111111111111111111101111111111111111111111111111000000000000000;
		6966: Delta = 69'sb000000000000000000000000100000000000000000000000000001000000000000000;
		7709: Delta = 69'sb111111111111111111111111100000000000000000000000000001000000000000000;
		43152: Delta = 69'sb000000000000000000000000011111111111111111111111111111000000000000000;
		43895: Delta = 69'sb111111111111111111111111011111111111111111111111111111000000000000000;
		32025: Delta = 69'sb000000000000000000000001000000000000000000000000000001000000000000000;
		33511: Delta = 69'sb111111111111111111111111000000000000000000000000000001000000000000000;
		17350: Delta = 69'sb000000000000000000000000111111111111111111111111111111000000000000000;
		18836: Delta = 69'sb111111111111111111111110111111111111111111111111111111000000000000000;
		31282: Delta = 69'sb000000000000000000000010000000000000000000000000000001000000000000000;
		34254: Delta = 69'sb111111111111111111111110000000000000000000000000000001000000000000000;
		16607: Delta = 69'sb000000000000000000000001111111111111111111111111111111000000000000000;
		19579: Delta = 69'sb111111111111111111111101111111111111111111111111111111000000000000000;
		29796: Delta = 69'sb000000000000000000000100000000000000000000000000000001000000000000000;
		35740: Delta = 69'sb111111111111111111111100000000000000000000000000000001000000000000000;
		15121: Delta = 69'sb000000000000000000000011111111111111111111111111111111000000000000000;
		21065: Delta = 69'sb111111111111111111111011111111111111111111111111111111000000000000000;
		26824: Delta = 69'sb000000000000000000001000000000000000000000000000000001000000000000000;
		38712: Delta = 69'sb111111111111111111111000000000000000000000000000000001000000000000000;
		12149: Delta = 69'sb000000000000000000000111111111111111111111111111111111000000000000000;
		24037: Delta = 69'sb111111111111111111110111111111111111111111111111111111000000000000000;
		20880: Delta = 69'sb000000000000000000010000000000000000000000000000000001000000000000000;
		44656: Delta = 69'sb111111111111111111110000000000000000000000000000000001000000000000000;
		6205: Delta = 69'sb000000000000000000001111111111111111111111111111111111000000000000000;
		29981: Delta = 69'sb111111111111111111101111111111111111111111111111111111000000000000000;
		8992: Delta = 69'sb000000000000000000100000000000000000000000000000000001000000000000000;
		5683: Delta = 69'sb111111111111111111100000000000000000000000000000000001000000000000000;
		45178: Delta = 69'sb000000000000000000011111111111111111111111111111111111000000000000000;
		41869: Delta = 69'sb111111111111111111011111111111111111111111111111111111000000000000000;
		36077: Delta = 69'sb000000000000000001000000000000000000000000000000000001000000000000000;
		29459: Delta = 69'sb111111111111111111000000000000000000000000000000000001000000000000000;
		21402: Delta = 69'sb000000000000000000111111111111111111111111111111111111000000000000000;
		14784: Delta = 69'sb111111111111111110111111111111111111111111111111111111000000000000000;
		39386: Delta = 69'sb000000000000000010000000000000000000000000000000000001000000000000000;
		26150: Delta = 69'sb111111111111111110000000000000000000000000000000000001000000000000000;
		24711: Delta = 69'sb000000000000000001111111111111111111111111111111111111000000000000000;
		11475: Delta = 69'sb111111111111111101111111111111111111111111111111111111000000000000000;
		46004: Delta = 69'sb000000000000000100000000000000000000000000000000000001000000000000000;
		19532: Delta = 69'sb111111111111111100000000000000000000000000000000000001000000000000000;
		31329: Delta = 69'sb000000000000000011111111111111111111111111111111111111000000000000000;
		4857: Delta = 69'sb111111111111111011111111111111111111111111111111111111000000000000000;
		8379: Delta = 69'sb000000000000001000000000000000000000000000000000000001000000000000000;
		6296: Delta = 69'sb111111111111111000000000000000000000000000000000000001000000000000000;
		44565: Delta = 69'sb000000000000000111111111111111111111111111111111111111000000000000000;
		42482: Delta = 69'sb111111111111110111111111111111111111111111111111111111000000000000000;
		34851: Delta = 69'sb000000000000010000000000000000000000000000000000000001000000000000000;
		30685: Delta = 69'sb111111111111110000000000000000000000000000000000000001000000000000000;
		20176: Delta = 69'sb000000000000001111111111111111111111111111111111111111000000000000000;
		16010: Delta = 69'sb111111111111101111111111111111111111111111111111111111000000000000000;
		36934: Delta = 69'sb000000000000100000000000000000000000000000000000000001000000000000000;
		28602: Delta = 69'sb111111111111100000000000000000000000000000000000000001000000000000000;
		22259: Delta = 69'sb000000000000011111111111111111111111111111111111111111000000000000000;
		13927: Delta = 69'sb111111111111011111111111111111111111111111111111111111000000000000000;
		41100: Delta = 69'sb000000000001000000000000000000000000000000000000000001000000000000000;
		24436: Delta = 69'sb111111111111000000000000000000000000000000000000000001000000000000000;
		26425: Delta = 69'sb000000000000111111111111111111111111111111111111111111000000000000000;
		9761: Delta = 69'sb111111111110111111111111111111111111111111111111111111000000000000000;
		49432: Delta = 69'sb000000000010000000000000000000000000000000000000000001000000000000000;
		16104: Delta = 69'sb111111111110000000000000000000000000000000000000000001000000000000000;
		34757: Delta = 69'sb000000000001111111111111111111111111111111111111111111000000000000000;
		1429: Delta = 69'sb111111111101111111111111111111111111111111111111111111000000000000000;
		15235: Delta = 69'sb000000000100000000000000000000000000000000000000000001000000000000000;
		50301: Delta = 69'sb111111111100000000000000000000000000000000000000000001000000000000000;
		560: Delta = 69'sb000000000011111111111111111111111111111111111111111111000000000000000;
		35626: Delta = 69'sb111111111011111111111111111111111111111111111111111111000000000000000;
		48563: Delta = 69'sb000000001000000000000000000000000000000000000000000001000000000000000;
		16973: Delta = 69'sb111111111000000000000000000000000000000000000000000001000000000000000;
		33888: Delta = 69'sb000000000111111111111111111111111111111111111111111111000000000000000;
		2298: Delta = 69'sb111111110111111111111111111111111111111111111111111111000000000000000;
		13497: Delta = 69'sb000000010000000000000000000000000000000000000000000001000000000000000;
		1178: Delta = 69'sb111111110000000000000000000000000000000000000000000001000000000000000;
		49683: Delta = 69'sb000000001111111111111111111111111111111111111111111111000000000000000;
		37364: Delta = 69'sb111111101111111111111111111111111111111111111111111111000000000000000;
		45087: Delta = 69'sb000000100000000000000000000000000000000000000000000001000000000000000;
		20449: Delta = 69'sb111111100000000000000000000000000000000000000000000001000000000000000;
		30412: Delta = 69'sb000000011111111111111111111111111111111111111111111111000000000000000;
		5774: Delta = 69'sb111111011111111111111111111111111111111111111111111111000000000000000;
		6545: Delta = 69'sb000001000000000000000000000000000000000000000000000001000000000000000;
		8130: Delta = 69'sb111111000000000000000000000000000000000000000000000001000000000000000;
		42731: Delta = 69'sb000000111111111111111111111111111111111111111111111111000000000000000;
		44316: Delta = 69'sb111110111111111111111111111111111111111111111111111111000000000000000;
		31183: Delta = 69'sb000010000000000000000000000000000000000000000000000001000000000000000;
		34353: Delta = 69'sb111110000000000000000000000000000000000000000000000001000000000000000;
		16508: Delta = 69'sb000001111111111111111111111111111111111111111111111111000000000000000;
		19678: Delta = 69'sb111101111111111111111111111111111111111111111111111111000000000000000;
		29598: Delta = 69'sb000100000000000000000000000000000000000000000000000001000000000000000;
		35938: Delta = 69'sb111100000000000000000000000000000000000000000000000001000000000000000;
		14923: Delta = 69'sb000011111111111111111111111111111111111111111111111111000000000000000;
		21263: Delta = 69'sb111011111111111111111111111111111111111111111111111111000000000000000;
		26428: Delta = 69'sb001000000000000000000000000000000000000000000000000001000000000000000;
		39108: Delta = 69'sb111000000000000000000000000000000000000000000000000001000000000000000;
		11753: Delta = 69'sb000111111111111111111111111111111111111111111111111111000000000000000;
		24433: Delta = 69'sb110111111111111111111111111111111111111111111111111111000000000000000;
		20088: Delta = 69'sb010000000000000000000000000000000000000000000000000001000000000000000;
		45448: Delta = 69'sb110000000000000000000000000000000000000000000000000001000000000000000;
		5413: Delta = 69'sb001111111111111111111111111111111111111111111111111111000000000000000;
		30773: Delta = 69'sb101111111111111111111111111111111111111111111111111111000000000000000;
		44025: Delta = 69'sb000000000000000000000000000000000000000000000000000110000000000000000;
		6836: Delta = 69'sb111111111111111111111111111111111111111111111111111010000000000000000;
		22514: Delta = 69'sb000000000000000000000000000000000000000000000000001010000000000000000;
		28347: Delta = 69'sb111111111111111111111111111111111111111111111111110110000000000000000;
		30353: Delta = 69'sb000000000000000000000000000000000000000000000000010010000000000000000;
		49858: Delta = 69'sb111111111111111111111111111111111111111111111111110010000000000000000;
		1003: Delta = 69'sb000000000000000000000000000000000000000000000000001110000000000000000;
		20508: Delta = 69'sb111111111111111111111111111111111111111111111111101110000000000000000;
		46031: Delta = 69'sb000000000000000000000000000000000000000000000000100010000000000000000;
		34180: Delta = 69'sb111111111111111111111111111111111111111111111111100010000000000000000;
		16681: Delta = 69'sb000000000000000000000000000000000000000000000000011110000000000000000;
		4830: Delta = 69'sb111111111111111111111111111111111111111111111111011110000000000000000;
		26526: Delta = 69'sb000000000000000000000000000000000000000000000001000010000000000000000;
		2824: Delta = 69'sb111111111111111111111111111111111111111111111111000010000000000000000;
		48037: Delta = 69'sb000000000000000000000000000000000000000000000000111110000000000000000;
		24335: Delta = 69'sb111111111111111111111111111111111111111111111110111110000000000000000;
		38377: Delta = 69'sb000000000000000000000000000000000000000000000010000010000000000000000;
		41834: Delta = 69'sb111111111111111111111111111111111111111111111110000010000000000000000;
		9027: Delta = 69'sb000000000000000000000000000000000000000000000001111110000000000000000;
		12484: Delta = 69'sb111111111111111111111111111111111111111111111101111110000000000000000;
		11218: Delta = 69'sb000000000000000000000000000000000000000000000100000010000000000000000;
		18132: Delta = 69'sb111111111111111111111111111111111111111111111100000010000000000000000;
		32729: Delta = 69'sb000000000000000000000000000000000000000000000011111110000000000000000;
		39643: Delta = 69'sb111111111111111111111111111111111111111111111011111110000000000000000;
		7761: Delta = 69'sb000000000000000000000000000000000000000000001000000010000000000000000;
		21589: Delta = 69'sb111111111111111111111111111111111111111111111000000010000000000000000;
		29272: Delta = 69'sb000000000000000000000000000000000000000000000111111110000000000000000;
		43100: Delta = 69'sb111111111111111111111111111111111111111111110111111110000000000000000;
		847: Delta = 69'sb000000000000000000000000000000000000000000010000000010000000000000000;
		28503: Delta = 69'sb111111111111111111111111111111111111111111110000000010000000000000000;
		22358: Delta = 69'sb000000000000000000000000000000000000000000001111111110000000000000000;
		50014: Delta = 69'sb111111111111111111111111111111111111111111101111111110000000000000000;
		37880: Delta = 69'sb000000000000000000000000000000000000000000100000000010000000000000000;
		42331: Delta = 69'sb111111111111111111111111111111111111111111100000000010000000000000000;
		8530: Delta = 69'sb000000000000000000000000000000000000000000011111111110000000000000000;
		12981: Delta = 69'sb111111111111111111111111111111111111111111011111111110000000000000000;
		10224: Delta = 69'sb000000000000000000000000000000000000000001000000000010000000000000000;
		19126: Delta = 69'sb111111111111111111111111111111111111111111000000000010000000000000000;
		31735: Delta = 69'sb000000000000000000000000000000000000000000111111111110000000000000000;
		40637: Delta = 69'sb111111111111111111111111111111111111111110111111111110000000000000000;
		5773: Delta = 69'sb000000000000000000000000000000000000000010000000000010000000000000000;
		23577: Delta = 69'sb111111111111111111111111111111111111111110000000000010000000000000000;
		27284: Delta = 69'sb000000000000000000000000000000000000000001111111111110000000000000000;
		45088: Delta = 69'sb111111111111111111111111111111111111111101111111111110000000000000000;
		47732: Delta = 69'sb000000000000000000000000000000000000000100000000000010000000000000000;
		32479: Delta = 69'sb111111111111111111111111111111111111111100000000000010000000000000000;
		18382: Delta = 69'sb000000000000000000000000000000000000000011111111111110000000000000000;
		3129: Delta = 69'sb111111111111111111111111111111111111111011111111111110000000000000000;
		29928: Delta = 69'sb000000000000000000000000000000000000001000000000000010000000000000000;
		50283: Delta = 69'sb111111111111111111111111111111111111111000000000000010000000000000000;
		578: Delta = 69'sb000000000000000000000000000000000000000111111111111110000000000000000;
		20933: Delta = 69'sb111111111111111111111111111111111111110111111111111110000000000000000;
		45181: Delta = 69'sb000000000000000000000000000000000000010000000000000010000000000000000;
		35030: Delta = 69'sb111111111111111111111111111111111111110000000000000010000000000000000;
		15831: Delta = 69'sb000000000000000000000000000000000000001111111111111110000000000000000;
		5680: Delta = 69'sb111111111111111111111111111111111111101111111111111110000000000000000;
		24826: Delta = 69'sb000000000000000000000000000000000000100000000000000010000000000000000;
		4524: Delta = 69'sb111111111111111111111111111111111111100000000000000010000000000000000;
		46337: Delta = 69'sb000000000000000000000000000000000000011111111111111110000000000000000;
		26035: Delta = 69'sb111111111111111111111111111111111111011111111111111110000000000000000;
		34977: Delta = 69'sb000000000000000000000000000000000001000000000000000010000000000000000;
		45234: Delta = 69'sb111111111111111111111111111111111111000000000000000010000000000000000;
		5627: Delta = 69'sb000000000000000000000000000000000000111111111111111110000000000000000;
		15884: Delta = 69'sb111111111111111111111111111111111110111111111111111110000000000000000;
		4418: Delta = 69'sb000000000000000000000000000000000010000000000000000010000000000000000;
		24932: Delta = 69'sb111111111111111111111111111111111110000000000000000010000000000000000;
		25929: Delta = 69'sb000000000000000000000000000000000001111111111111111110000000000000000;
		46443: Delta = 69'sb111111111111111111111111111111111101111111111111111110000000000000000;
		45022: Delta = 69'sb000000000000000000000000000000000100000000000000000010000000000000000;
		35189: Delta = 69'sb111111111111111111111111111111111100000000000000000010000000000000000;
		15672: Delta = 69'sb000000000000000000000000000000000011111111111111111110000000000000000;
		5839: Delta = 69'sb111111111111111111111111111111111011111111111111111110000000000000000;
		24508: Delta = 69'sb000000000000000000000000000000001000000000000000000010000000000000000;
		4842: Delta = 69'sb111111111111111111111111111111111000000000000000000010000000000000000;
		46019: Delta = 69'sb000000000000000000000000000000000111111111111111111110000000000000000;
		26353: Delta = 69'sb111111111111111111111111111111110111111111111111111110000000000000000;
		34341: Delta = 69'sb000000000000000000000000000000010000000000000000000010000000000000000;
		45870: Delta = 69'sb111111111111111111111111111111110000000000000000000010000000000000000;
		4991: Delta = 69'sb000000000000000000000000000000001111111111111111111110000000000000000;
		16520: Delta = 69'sb111111111111111111111111111111101111111111111111111110000000000000000;
		3146: Delta = 69'sb000000000000000000000000000000100000000000000000000010000000000000000;
		26204: Delta = 69'sb111111111111111111111111111111100000000000000000000010000000000000000;
		24657: Delta = 69'sb000000000000000000000000000000011111111111111111111110000000000000000;
		47715: Delta = 69'sb111111111111111111111111111111011111111111111111111110000000000000000;
		42478: Delta = 69'sb000000000000000000000000000001000000000000000000000010000000000000000;
		37733: Delta = 69'sb111111111111111111111111111111000000000000000000000010000000000000000;
		13128: Delta = 69'sb000000000000000000000000000000111111111111111111111110000000000000000;
		8383: Delta = 69'sb111111111111111111111111111110111111111111111111111110000000000000000;
		19420: Delta = 69'sb000000000000000000000000000010000000000000000000000010000000000000000;
		9930: Delta = 69'sb111111111111111111111111111110000000000000000000000010000000000000000;
		40931: Delta = 69'sb000000000000000000000000000001111111111111111111111110000000000000000;
		31441: Delta = 69'sb111111111111111111111111111101111111111111111111111110000000000000000;
		24165: Delta = 69'sb000000000000000000000000000100000000000000000000000010000000000000000;
		5185: Delta = 69'sb111111111111111111111111111100000000000000000000000010000000000000000;
		45676: Delta = 69'sb000000000000000000000000000011111111111111111111111110000000000000000;
		26696: Delta = 69'sb111111111111111111111111111011111111111111111111111110000000000000000;
		33655: Delta = 69'sb000000000000000000000000001000000000000000000000000010000000000000000;
		46556: Delta = 69'sb111111111111111111111111111000000000000000000000000010000000000000000;
		4305: Delta = 69'sb000000000000000000000000000111111111111111111111111110000000000000000;
		17206: Delta = 69'sb111111111111111111111111110111111111111111111111111110000000000000000;
		1774: Delta = 69'sb000000000000000000000000010000000000000000000000000010000000000000000;
		27576: Delta = 69'sb111111111111111111111111110000000000000000000000000010000000000000000;
		23285: Delta = 69'sb000000000000000000000000001111111111111111111111111110000000000000000;
		49087: Delta = 69'sb111111111111111111111111101111111111111111111111111110000000000000000;
		39734: Delta = 69'sb000000000000000000000000100000000000000000000000000010000000000000000;
		40477: Delta = 69'sb111111111111111111111111100000000000000000000000000010000000000000000;
		10384: Delta = 69'sb000000000000000000000000011111111111111111111111111110000000000000000;
		11127: Delta = 69'sb111111111111111111111111011111111111111111111111111110000000000000000;
		13932: Delta = 69'sb000000000000000000000001000000000000000000000000000010000000000000000;
		15418: Delta = 69'sb111111111111111111111111000000000000000000000000000010000000000000000;
		35443: Delta = 69'sb000000000000000000000000111111111111111111111111111110000000000000000;
		36929: Delta = 69'sb111111111111111111111110111111111111111111111111111110000000000000000;
		13189: Delta = 69'sb000000000000000000000010000000000000000000000000000010000000000000000;
		16161: Delta = 69'sb111111111111111111111110000000000000000000000000000010000000000000000;
		34700: Delta = 69'sb000000000000000000000001111111111111111111111111111110000000000000000;
		37672: Delta = 69'sb111111111111111111111101111111111111111111111111111110000000000000000;
		11703: Delta = 69'sb000000000000000000000100000000000000000000000000000010000000000000000;
		17647: Delta = 69'sb111111111111111111111100000000000000000000000000000010000000000000000;
		33214: Delta = 69'sb000000000000000000000011111111111111111111111111111110000000000000000;
		39158: Delta = 69'sb111111111111111111111011111111111111111111111111111110000000000000000;
		8731: Delta = 69'sb000000000000000000001000000000000000000000000000000010000000000000000;
		20619: Delta = 69'sb111111111111111111111000000000000000000000000000000010000000000000000;
		30242: Delta = 69'sb000000000000000000000111111111111111111111111111111110000000000000000;
		42130: Delta = 69'sb111111111111111111110111111111111111111111111111111110000000000000000;
		2787: Delta = 69'sb000000000000000000010000000000000000000000000000000010000000000000000;
		26563: Delta = 69'sb111111111111111111110000000000000000000000000000000010000000000000000;
		24298: Delta = 69'sb000000000000000000001111111111111111111111111111111110000000000000000;
		48074: Delta = 69'sb111111111111111111101111111111111111111111111111111110000000000000000;
		41760: Delta = 69'sb000000000000000000100000000000000000000000000000000010000000000000000;
		38451: Delta = 69'sb111111111111111111100000000000000000000000000000000010000000000000000;
		12410: Delta = 69'sb000000000000000000011111111111111111111111111111111110000000000000000;
		9101: Delta = 69'sb111111111111111111011111111111111111111111111111111110000000000000000;
		17984: Delta = 69'sb000000000000000001000000000000000000000000000000000010000000000000000;
		11366: Delta = 69'sb111111111111111111000000000000000000000000000000000010000000000000000;
		39495: Delta = 69'sb000000000000000000111111111111111111111111111111111110000000000000000;
		32877: Delta = 69'sb111111111111111110111111111111111111111111111111111110000000000000000;
		21293: Delta = 69'sb000000000000000010000000000000000000000000000000000010000000000000000;
		8057: Delta = 69'sb111111111111111110000000000000000000000000000000000010000000000000000;
		42804: Delta = 69'sb000000000000000001111111111111111111111111111111111110000000000000000;
		29568: Delta = 69'sb111111111111111101111111111111111111111111111111111110000000000000000;
		27911: Delta = 69'sb000000000000000100000000000000000000000000000000000010000000000000000;
		1439: Delta = 69'sb111111111111111100000000000000000000000000000000000010000000000000000;
		49422: Delta = 69'sb000000000000000011111111111111111111111111111111111110000000000000000;
		22950: Delta = 69'sb111111111111111011111111111111111111111111111111111110000000000000000;
		41147: Delta = 69'sb000000000000001000000000000000000000000000000000000010000000000000000;
		39064: Delta = 69'sb111111111111111000000000000000000000000000000000000010000000000000000;
		11797: Delta = 69'sb000000000000000111111111111111111111111111111111111110000000000000000;
		9714: Delta = 69'sb111111111111110111111111111111111111111111111111111110000000000000000;
		16758: Delta = 69'sb000000000000010000000000000000000000000000000000000010000000000000000;
		12592: Delta = 69'sb111111111111110000000000000000000000000000000000000010000000000000000;
		38269: Delta = 69'sb000000000000001111111111111111111111111111111111111110000000000000000;
		34103: Delta = 69'sb111111111111101111111111111111111111111111111111111110000000000000000;
		18841: Delta = 69'sb000000000000100000000000000000000000000000000000000010000000000000000;
		10509: Delta = 69'sb111111111111100000000000000000000000000000000000000010000000000000000;
		40352: Delta = 69'sb000000000000011111111111111111111111111111111111111110000000000000000;
		32020: Delta = 69'sb111111111111011111111111111111111111111111111111111110000000000000000;
		23007: Delta = 69'sb000000000001000000000000000000000000000000000000000010000000000000000;
		6343: Delta = 69'sb111111111111000000000000000000000000000000000000000010000000000000000;
		44518: Delta = 69'sb000000000000111111111111111111111111111111111111111110000000000000000;
		27854: Delta = 69'sb111111111110111111111111111111111111111111111111111110000000000000000;
		31339: Delta = 69'sb000000000010000000000000000000000000000000000000000010000000000000000;
		48872: Delta = 69'sb111111111110000000000000000000000000000000000000000010000000000000000;
		1989: Delta = 69'sb000000000001111111111111111111111111111111111111111110000000000000000;
		19522: Delta = 69'sb111111111101111111111111111111111111111111111111111110000000000000000;
		48003: Delta = 69'sb000000000100000000000000000000000000000000000000000010000000000000000;
		32208: Delta = 69'sb111111111100000000000000000000000000000000000000000010000000000000000;
		18653: Delta = 69'sb000000000011111111111111111111111111111111111111111110000000000000000;
		2858: Delta = 69'sb111111111011111111111111111111111111111111111111111110000000000000000;
		30470: Delta = 69'sb000000001000000000000000000000000000000000000000000010000000000000000;
		49741: Delta = 69'sb111111111000000000000000000000000000000000000000000010000000000000000;
		1120: Delta = 69'sb000000000111111111111111111111111111111111111111111110000000000000000;
		20391: Delta = 69'sb111111110111111111111111111111111111111111111111111110000000000000000;
		46265: Delta = 69'sb000000010000000000000000000000000000000000000000000010000000000000000;
		33946: Delta = 69'sb111111110000000000000000000000000000000000000000000010000000000000000;
		16915: Delta = 69'sb000000001111111111111111111111111111111111111111111110000000000000000;
		4596: Delta = 69'sb111111101111111111111111111111111111111111111111111110000000000000000;
		26994: Delta = 69'sb000000100000000000000000000000000000000000000000000010000000000000000;
		2356: Delta = 69'sb111111100000000000000000000000000000000000000000000010000000000000000;
		48505: Delta = 69'sb000000011111111111111111111111111111111111111111111110000000000000000;
		23867: Delta = 69'sb111111011111111111111111111111111111111111111111111110000000000000000;
		39313: Delta = 69'sb000001000000000000000000000000000000000000000000000010000000000000000;
		40898: Delta = 69'sb111111000000000000000000000000000000000000000000000010000000000000000;
		9963: Delta = 69'sb000000111111111111111111111111111111111111111111111110000000000000000;
		11548: Delta = 69'sb111110111111111111111111111111111111111111111111111110000000000000000;
		13090: Delta = 69'sb000010000000000000000000000000000000000000000000000010000000000000000;
		16260: Delta = 69'sb111110000000000000000000000000000000000000000000000010000000000000000;
		34601: Delta = 69'sb000001111111111111111111111111111111111111111111111110000000000000000;
		37771: Delta = 69'sb111101111111111111111111111111111111111111111111111110000000000000000;
		11505: Delta = 69'sb000100000000000000000000000000000000000000000000000010000000000000000;
		17845: Delta = 69'sb111100000000000000000000000000000000000000000000000010000000000000000;
		33016: Delta = 69'sb000011111111111111111111111111111111111111111111111110000000000000000;
		39356: Delta = 69'sb111011111111111111111111111111111111111111111111111110000000000000000;
		8335: Delta = 69'sb001000000000000000000000000000000000000000000000000010000000000000000;
		21015: Delta = 69'sb111000000000000000000000000000000000000000000000000010000000000000000;
		29846: Delta = 69'sb000111111111111111111111111111111111111111111111111110000000000000000;
		42526: Delta = 69'sb110111111111111111111111111111111111111111111111111110000000000000000;
		1995: Delta = 69'sb010000000000000000000000000000000000000000000000000010000000000000000;
		27355: Delta = 69'sb110000000000000000000000000000000000000000000000000010000000000000000;
		23506: Delta = 69'sb001111111111111111111111111111111111111111111111111110000000000000000;
		48866: Delta = 69'sb101111111111111111111111111111111111111111111111111110000000000000000;
		37189: Delta = 69'sb000000000000000000000000000000000000000000000000001100000000000000000;
		13672: Delta = 69'sb111111111111111111111111111111111111111111111111110100000000000000000;
		45028: Delta = 69'sb000000000000000000000000000000000000000000000000010100000000000000000;
		5833: Delta = 69'sb111111111111111111111111111111111111111111111111101100000000000000000;
		9845: Delta = 69'sb000000000000000000000000000000000000000000000000100100000000000000000;
		48855: Delta = 69'sb111111111111111111111111111111111111111111111111100100000000000000000;
		2006: Delta = 69'sb000000000000000000000000000000000000000000000000011100000000000000000;
		41016: Delta = 69'sb111111111111111111111111111111111111111111111111011100000000000000000;
		41201: Delta = 69'sb000000000000000000000000000000000000000000000001000100000000000000000;
		17499: Delta = 69'sb111111111111111111111111111111111111111111111111000100000000000000000;
		33362: Delta = 69'sb000000000000000000000000000000000000000000000000111100000000000000000;
		9660: Delta = 69'sb111111111111111111111111111111111111111111111110111100000000000000000;
		2191: Delta = 69'sb000000000000000000000000000000000000000000000010000100000000000000000;
		5648: Delta = 69'sb111111111111111111111111111111111111111111111110000100000000000000000;
		45213: Delta = 69'sb000000000000000000000000000000000000000000000001111100000000000000000;
		48670: Delta = 69'sb111111111111111111111111111111111111111111111101111100000000000000000;
		25893: Delta = 69'sb000000000000000000000000000000000000000000000100000100000000000000000;
		32807: Delta = 69'sb111111111111111111111111111111111111111111111100000100000000000000000;
		18054: Delta = 69'sb000000000000000000000000000000000000000000000011111100000000000000000;
		24968: Delta = 69'sb111111111111111111111111111111111111111111111011111100000000000000000;
		22436: Delta = 69'sb000000000000000000000000000000000000000000001000000100000000000000000;
		36264: Delta = 69'sb111111111111111111111111111111111111111111111000000100000000000000000;
		14597: Delta = 69'sb000000000000000000000000000000000000000000000111111100000000000000000;
		28425: Delta = 69'sb111111111111111111111111111111111111111111110111111100000000000000000;
		15522: Delta = 69'sb000000000000000000000000000000000000000000010000000100000000000000000;
		43178: Delta = 69'sb111111111111111111111111111111111111111111110000000100000000000000000;
		7683: Delta = 69'sb000000000000000000000000000000000000000000001111111100000000000000000;
		35339: Delta = 69'sb111111111111111111111111111111111111111111101111111100000000000000000;
		1694: Delta = 69'sb000000000000000000000000000000000000000000100000000100000000000000000;
		6145: Delta = 69'sb111111111111111111111111111111111111111111100000000100000000000000000;
		44716: Delta = 69'sb000000000000000000000000000000000000000000011111111100000000000000000;
		49167: Delta = 69'sb111111111111111111111111111111111111111111011111111100000000000000000;
		24899: Delta = 69'sb000000000000000000000000000000000000000001000000000100000000000000000;
		33801: Delta = 69'sb111111111111111111111111111111111111111111000000000100000000000000000;
		17060: Delta = 69'sb000000000000000000000000000000000000000000111111111100000000000000000;
		25962: Delta = 69'sb111111111111111111111111111111111111111110111111111100000000000000000;
		20448: Delta = 69'sb000000000000000000000000000000000000000010000000000100000000000000000;
		38252: Delta = 69'sb111111111111111111111111111111111111111110000000000100000000000000000;
		12609: Delta = 69'sb000000000000000000000000000000000000000001111111111100000000000000000;
		30413: Delta = 69'sb111111111111111111111111111111111111111101111111111100000000000000000;
		11546: Delta = 69'sb000000000000000000000000000000000000000100000000000100000000000000000;
		47154: Delta = 69'sb111111111111111111111111111111111111111100000000000100000000000000000;
		3707: Delta = 69'sb000000000000000000000000000000000000000011111111111100000000000000000;
		39315: Delta = 69'sb111111111111111111111111111111111111111011111111111100000000000000000;
		44603: Delta = 69'sb000000000000000000000000000000000000001000000000000100000000000000000;
		14097: Delta = 69'sb111111111111111111111111111111111111111000000000000100000000000000000;
		36764: Delta = 69'sb000000000000000000000000000000000000000111111111111100000000000000000;
		6258: Delta = 69'sb111111111111111111111111111111111111110111111111111100000000000000000;
		8995: Delta = 69'sb000000000000000000000000000000000000010000000000000100000000000000000;
		49705: Delta = 69'sb111111111111111111111111111111111111110000000000000100000000000000000;
		1156: Delta = 69'sb000000000000000000000000000000000000001111111111111100000000000000000;
		41866: Delta = 69'sb111111111111111111111111111111111111101111111111111100000000000000000;
		39501: Delta = 69'sb000000000000000000000000000000000000100000000000000100000000000000000;
		19199: Delta = 69'sb111111111111111111111111111111111111100000000000000100000000000000000;
		31662: Delta = 69'sb000000000000000000000000000000000000011111111111111100000000000000000;
		11360: Delta = 69'sb111111111111111111111111111111111111011111111111111100000000000000000;
		49652: Delta = 69'sb000000000000000000000000000000000001000000000000000100000000000000000;
		9048: Delta = 69'sb111111111111111111111111111111111111000000000000000100000000000000000;
		41813: Delta = 69'sb000000000000000000000000000000000000111111111111111100000000000000000;
		1209: Delta = 69'sb111111111111111111111111111111111110111111111111111100000000000000000;
		19093: Delta = 69'sb000000000000000000000000000000000010000000000000000100000000000000000;
		39607: Delta = 69'sb111111111111111111111111111111111110000000000000000100000000000000000;
		11254: Delta = 69'sb000000000000000000000000000000000001111111111111111100000000000000000;
		31768: Delta = 69'sb111111111111111111111111111111111101111111111111111100000000000000000;
		8836: Delta = 69'sb000000000000000000000000000000000100000000000000000100000000000000000;
		49864: Delta = 69'sb111111111111111111111111111111111100000000000000000100000000000000000;
		997: Delta = 69'sb000000000000000000000000000000000011111111111111111100000000000000000;
		42025: Delta = 69'sb111111111111111111111111111111111011111111111111111100000000000000000;
		39183: Delta = 69'sb000000000000000000000000000000001000000000000000000100000000000000000;
		19517: Delta = 69'sb111111111111111111111111111111111000000000000000000100000000000000000;
		31344: Delta = 69'sb000000000000000000000000000000000111111111111111111100000000000000000;
		11678: Delta = 69'sb111111111111111111111111111111110111111111111111111100000000000000000;
		49016: Delta = 69'sb000000000000000000000000000000010000000000000000000100000000000000000;
		9684: Delta = 69'sb111111111111111111111111111111110000000000000000000100000000000000000;
		41177: Delta = 69'sb000000000000000000000000000000001111111111111111111100000000000000000;
		1845: Delta = 69'sb111111111111111111111111111111101111111111111111111100000000000000000;
		17821: Delta = 69'sb000000000000000000000000000000100000000000000000000100000000000000000;
		40879: Delta = 69'sb111111111111111111111111111111100000000000000000000100000000000000000;
		9982: Delta = 69'sb000000000000000000000000000000011111111111111111111100000000000000000;
		33040: Delta = 69'sb111111111111111111111111111111011111111111111111111100000000000000000;
		6292: Delta = 69'sb000000000000000000000000000001000000000000000000000100000000000000000;
		1547: Delta = 69'sb111111111111111111111111111111000000000000000000000100000000000000000;
		49314: Delta = 69'sb000000000000000000000000000000111111111111111111111100000000000000000;
		44569: Delta = 69'sb111111111111111111111111111110111111111111111111111100000000000000000;
		34095: Delta = 69'sb000000000000000000000000000010000000000000000000000100000000000000000;
		24605: Delta = 69'sb111111111111111111111111111110000000000000000000000100000000000000000;
		26256: Delta = 69'sb000000000000000000000000000001111111111111111111111100000000000000000;
		16766: Delta = 69'sb111111111111111111111111111101111111111111111111111100000000000000000;
		38840: Delta = 69'sb000000000000000000000000000100000000000000000000000100000000000000000;
		19860: Delta = 69'sb111111111111111111111111111100000000000000000000000100000000000000000;
		31001: Delta = 69'sb000000000000000000000000000011111111111111111111111100000000000000000;
		12021: Delta = 69'sb111111111111111111111111111011111111111111111111111100000000000000000;
		48330: Delta = 69'sb000000000000000000000000001000000000000000000000000100000000000000000;
		10370: Delta = 69'sb111111111111111111111111111000000000000000000000000100000000000000000;
		40491: Delta = 69'sb000000000000000000000000000111111111111111111111111100000000000000000;
		2531: Delta = 69'sb111111111111111111111111110111111111111111111111111100000000000000000;
		16449: Delta = 69'sb000000000000000000000000010000000000000000000000000100000000000000000;
		42251: Delta = 69'sb111111111111111111111111110000000000000000000000000100000000000000000;
		8610: Delta = 69'sb000000000000000000000000001111111111111111111111111100000000000000000;
		34412: Delta = 69'sb111111111111111111111111101111111111111111111111111100000000000000000;
		3548: Delta = 69'sb000000000000000000000000100000000000000000000000000100000000000000000;
		4291: Delta = 69'sb111111111111111111111111100000000000000000000000000100000000000000000;
		46570: Delta = 69'sb000000000000000000000000011111111111111111111111111100000000000000000;
		47313: Delta = 69'sb111111111111111111111111011111111111111111111111111100000000000000000;
		28607: Delta = 69'sb000000000000000000000001000000000000000000000000000100000000000000000;
		30093: Delta = 69'sb111111111111111111111111000000000000000000000000000100000000000000000;
		20768: Delta = 69'sb000000000000000000000000111111111111111111111111111100000000000000000;
		22254: Delta = 69'sb111111111111111111111110111111111111111111111111111100000000000000000;
		27864: Delta = 69'sb000000000000000000000010000000000000000000000000000100000000000000000;
		30836: Delta = 69'sb111111111111111111111110000000000000000000000000000100000000000000000;
		20025: Delta = 69'sb000000000000000000000001111111111111111111111111111100000000000000000;
		22997: Delta = 69'sb111111111111111111111101111111111111111111111111111100000000000000000;
		26378: Delta = 69'sb000000000000000000000100000000000000000000000000000100000000000000000;
		32322: Delta = 69'sb111111111111111111111100000000000000000000000000000100000000000000000;
		18539: Delta = 69'sb000000000000000000000011111111111111111111111111111100000000000000000;
		24483: Delta = 69'sb111111111111111111111011111111111111111111111111111100000000000000000;
		23406: Delta = 69'sb000000000000000000001000000000000000000000000000000100000000000000000;
		35294: Delta = 69'sb111111111111111111111000000000000000000000000000000100000000000000000;
		15567: Delta = 69'sb000000000000000000000111111111111111111111111111111100000000000000000;
		27455: Delta = 69'sb111111111111111111110111111111111111111111111111111100000000000000000;
		17462: Delta = 69'sb000000000000000000010000000000000000000000000000000100000000000000000;
		41238: Delta = 69'sb111111111111111111110000000000000000000000000000000100000000000000000;
		9623: Delta = 69'sb000000000000000000001111111111111111111111111111111100000000000000000;
		33399: Delta = 69'sb111111111111111111101111111111111111111111111111111100000000000000000;
		5574: Delta = 69'sb000000000000000000100000000000000000000000000000000100000000000000000;
		2265: Delta = 69'sb111111111111111111100000000000000000000000000000000100000000000000000;
		48596: Delta = 69'sb000000000000000000011111111111111111111111111111111100000000000000000;
		45287: Delta = 69'sb111111111111111111011111111111111111111111111111111100000000000000000;
		32659: Delta = 69'sb000000000000000001000000000000000000000000000000000100000000000000000;
		26041: Delta = 69'sb111111111111111111000000000000000000000000000000000100000000000000000;
		24820: Delta = 69'sb000000000000000000111111111111111111111111111111111100000000000000000;
		18202: Delta = 69'sb111111111111111110111111111111111111111111111111111100000000000000000;
		35968: Delta = 69'sb000000000000000010000000000000000000000000000000000100000000000000000;
		22732: Delta = 69'sb111111111111111110000000000000000000000000000000000100000000000000000;
		28129: Delta = 69'sb000000000000000001111111111111111111111111111111111100000000000000000;
		14893: Delta = 69'sb111111111111111101111111111111111111111111111111111100000000000000000;
		42586: Delta = 69'sb000000000000000100000000000000000000000000000000000100000000000000000;
		16114: Delta = 69'sb111111111111111100000000000000000000000000000000000100000000000000000;
		34747: Delta = 69'sb000000000000000011111111111111111111111111111111111100000000000000000;
		8275: Delta = 69'sb111111111111111011111111111111111111111111111111111100000000000000000;
		4961: Delta = 69'sb000000000000001000000000000000000000000000000000000100000000000000000;
		2878: Delta = 69'sb111111111111111000000000000000000000000000000000000100000000000000000;
		47983: Delta = 69'sb000000000000000111111111111111111111111111111111111100000000000000000;
		45900: Delta = 69'sb111111111111110111111111111111111111111111111111111100000000000000000;
		31433: Delta = 69'sb000000000000010000000000000000000000000000000000000100000000000000000;
		27267: Delta = 69'sb111111111111110000000000000000000000000000000000000100000000000000000;
		23594: Delta = 69'sb000000000000001111111111111111111111111111111111111100000000000000000;
		19428: Delta = 69'sb111111111111101111111111111111111111111111111111111100000000000000000;
		33516: Delta = 69'sb000000000000100000000000000000000000000000000000000100000000000000000;
		25184: Delta = 69'sb111111111111100000000000000000000000000000000000000100000000000000000;
		25677: Delta = 69'sb000000000000011111111111111111111111111111111111111100000000000000000;
		17345: Delta = 69'sb111111111111011111111111111111111111111111111111111100000000000000000;
		37682: Delta = 69'sb000000000001000000000000000000000000000000000000000100000000000000000;
		21018: Delta = 69'sb111111111111000000000000000000000000000000000000000100000000000000000;
		29843: Delta = 69'sb000000000000111111111111111111111111111111111111111100000000000000000;
		13179: Delta = 69'sb111111111110111111111111111111111111111111111111111100000000000000000;
		46014: Delta = 69'sb000000000010000000000000000000000000000000000000000100000000000000000;
		12686: Delta = 69'sb111111111110000000000000000000000000000000000000000100000000000000000;
		38175: Delta = 69'sb000000000001111111111111111111111111111111111111111100000000000000000;
		4847: Delta = 69'sb111111111101111111111111111111111111111111111111111100000000000000000;
		11817: Delta = 69'sb000000000100000000000000000000000000000000000000000100000000000000000;
		46883: Delta = 69'sb111111111100000000000000000000000000000000000000000100000000000000000;
		3978: Delta = 69'sb000000000011111111111111111111111111111111111111111100000000000000000;
		39044: Delta = 69'sb111111111011111111111111111111111111111111111111111100000000000000000;
		45145: Delta = 69'sb000000001000000000000000000000000000000000000000000100000000000000000;
		13555: Delta = 69'sb111111111000000000000000000000000000000000000000000100000000000000000;
		37306: Delta = 69'sb000000000111111111111111111111111111111111111111111100000000000000000;
		5716: Delta = 69'sb111111110111111111111111111111111111111111111111111100000000000000000;
		10079: Delta = 69'sb000000010000000000000000000000000000000000000000000100000000000000000;
		48621: Delta = 69'sb111111110000000000000000000000000000000000000000000100000000000000000;
		2240: Delta = 69'sb000000001111111111111111111111111111111111111111111100000000000000000;
		40782: Delta = 69'sb111111101111111111111111111111111111111111111111111100000000000000000;
		41669: Delta = 69'sb000000100000000000000000000000000000000000000000000100000000000000000;
		17031: Delta = 69'sb111111100000000000000000000000000000000000000000000100000000000000000;
		33830: Delta = 69'sb000000011111111111111111111111111111111111111111111100000000000000000;
		9192: Delta = 69'sb111111011111111111111111111111111111111111111111111100000000000000000;
		3127: Delta = 69'sb000001000000000000000000000000000000000000000000000100000000000000000;
		4712: Delta = 69'sb111111000000000000000000000000000000000000000000000100000000000000000;
		46149: Delta = 69'sb000000111111111111111111111111111111111111111111111100000000000000000;
		47734: Delta = 69'sb111110111111111111111111111111111111111111111111111100000000000000000;
		27765: Delta = 69'sb000010000000000000000000000000000000000000000000000100000000000000000;
		30935: Delta = 69'sb111110000000000000000000000000000000000000000000000100000000000000000;
		19926: Delta = 69'sb000001111111111111111111111111111111111111111111111100000000000000000;
		23096: Delta = 69'sb111101111111111111111111111111111111111111111111111100000000000000000;
		26180: Delta = 69'sb000100000000000000000000000000000000000000000000000100000000000000000;
		32520: Delta = 69'sb111100000000000000000000000000000000000000000000000100000000000000000;
		18341: Delta = 69'sb000011111111111111111111111111111111111111111111111100000000000000000;
		24681: Delta = 69'sb111011111111111111111111111111111111111111111111111100000000000000000;
		23010: Delta = 69'sb001000000000000000000000000000000000000000000000000100000000000000000;
		35690: Delta = 69'sb111000000000000000000000000000000000000000000000000100000000000000000;
		15171: Delta = 69'sb000111111111111111111111111111111111111111111111111100000000000000000;
		27851: Delta = 69'sb110111111111111111111111111111111111111111111111111100000000000000000;
		16670: Delta = 69'sb010000000000000000000000000000000000000000000000000100000000000000000;
		42030: Delta = 69'sb110000000000000000000000000000000000000000000000000100000000000000000;
		8831: Delta = 69'sb001111111111111111111111111111111111111111111111111100000000000000000;
		34191: Delta = 69'sb101111111111111111111111111111111111111111111111111100000000000000000;
		23517: Delta = 69'sb000000000000000000000000000000000000000000000000011000000000000000000;
		27344: Delta = 69'sb111111111111111111111111111111111111111111111111101000000000000000000;
		39195: Delta = 69'sb000000000000000000000000000000000000000000000000101000000000000000000;
		11666: Delta = 69'sb111111111111111111111111111111111111111111111111011000000000000000000;
		19690: Delta = 69'sb000000000000000000000000000000000000000000000001001000000000000000000;
		46849: Delta = 69'sb111111111111111111111111111111111111111111111111001000000000000000000;
		4012: Delta = 69'sb000000000000000000000000000000000000000000000000111000000000000000000;
		31171: Delta = 69'sb111111111111111111111111111111111111111111111110111000000000000000000;
		31541: Delta = 69'sb000000000000000000000000000000000000000000000010001000000000000000000;
		34998: Delta = 69'sb111111111111111111111111111111111111111111111110001000000000000000000;
		15863: Delta = 69'sb000000000000000000000000000000000000000000000001111000000000000000000;
		19320: Delta = 69'sb111111111111111111111111111111111111111111111101111000000000000000000;
		4382: Delta = 69'sb000000000000000000000000000000000000000000000100001000000000000000000;
		11296: Delta = 69'sb111111111111111111111111111111111111111111111100001000000000000000000;
		39565: Delta = 69'sb000000000000000000000000000000000000000000000011111000000000000000000;
		46479: Delta = 69'sb111111111111111111111111111111111111111111111011111000000000000000000;
		925: Delta = 69'sb000000000000000000000000000000000000000000001000001000000000000000000;
		14753: Delta = 69'sb111111111111111111111111111111111111111111111000001000000000000000000;
		36108: Delta = 69'sb000000000000000000000000000000000000000000000111111000000000000000000;
		49936: Delta = 69'sb111111111111111111111111111111111111111111110111111000000000000000000;
		44872: Delta = 69'sb000000000000000000000000000000000000000000010000001000000000000000000;
		21667: Delta = 69'sb111111111111111111111111111111111111111111110000001000000000000000000;
		29194: Delta = 69'sb000000000000000000000000000000000000000000001111111000000000000000000;
		5989: Delta = 69'sb111111111111111111111111111111111111111111101111111000000000000000000;
		31044: Delta = 69'sb000000000000000000000000000000000000000000100000001000000000000000000;
		35495: Delta = 69'sb111111111111111111111111111111111111111111100000001000000000000000000;
		15366: Delta = 69'sb000000000000000000000000000000000000000000011111111000000000000000000;
		19817: Delta = 69'sb111111111111111111111111111111111111111111011111111000000000000000000;
		3388: Delta = 69'sb000000000000000000000000000000000000000001000000001000000000000000000;
		12290: Delta = 69'sb111111111111111111111111111111111111111111000000001000000000000000000;
		38571: Delta = 69'sb000000000000000000000000000000000000000000111111111000000000000000000;
		47473: Delta = 69'sb111111111111111111111111111111111111111110111111111000000000000000000;
		49798: Delta = 69'sb000000000000000000000000000000000000000010000000001000000000000000000;
		16741: Delta = 69'sb111111111111111111111111111111111111111110000000001000000000000000000;
		34120: Delta = 69'sb000000000000000000000000000000000000000001111111111000000000000000000;
		1063: Delta = 69'sb111111111111111111111111111111111111111101111111111000000000000000000;
		40896: Delta = 69'sb000000000000000000000000000000000000000100000000001000000000000000000;
		25643: Delta = 69'sb111111111111111111111111111111111111111100000000001000000000000000000;
		25218: Delta = 69'sb000000000000000000000000000000000000000011111111111000000000000000000;
		9965: Delta = 69'sb111111111111111111111111111111111111111011111111111000000000000000000;
		23092: Delta = 69'sb000000000000000000000000000000000000001000000000001000000000000000000;
		43447: Delta = 69'sb111111111111111111111111111111111111111000000000001000000000000000000;
		7414: Delta = 69'sb000000000000000000000000000000000000000111111111111000000000000000000;
		27769: Delta = 69'sb111111111111111111111111111111111111110111111111111000000000000000000;
		38345: Delta = 69'sb000000000000000000000000000000000000010000000000001000000000000000000;
		28194: Delta = 69'sb111111111111111111111111111111111111110000000000001000000000000000000;
		22667: Delta = 69'sb000000000000000000000000000000000000001111111111111000000000000000000;
		12516: Delta = 69'sb111111111111111111111111111111111111101111111111111000000000000000000;
		17990: Delta = 69'sb000000000000000000000000000000000000100000000000001000000000000000000;
		48549: Delta = 69'sb111111111111111111111111111111111111100000000000001000000000000000000;
		2312: Delta = 69'sb000000000000000000000000000000000000011111111111111000000000000000000;
		32871: Delta = 69'sb111111111111111111111111111111111111011111111111111000000000000000000;
		28141: Delta = 69'sb000000000000000000000000000000000001000000000000001000000000000000000;
		38398: Delta = 69'sb111111111111111111111111111111111111000000000000001000000000000000000;
		12463: Delta = 69'sb000000000000000000000000000000000000111111111111111000000000000000000;
		22720: Delta = 69'sb111111111111111111111111111111111110111111111111111000000000000000000;
		48443: Delta = 69'sb000000000000000000000000000000000010000000000000001000000000000000000;
		18096: Delta = 69'sb111111111111111111111111111111111110000000000000001000000000000000000;
		32765: Delta = 69'sb000000000000000000000000000000000001111111111111111000000000000000000;
		2418: Delta = 69'sb111111111111111111111111111111111101111111111111111000000000000000000;
		38186: Delta = 69'sb000000000000000000000000000000000100000000000000001000000000000000000;
		28353: Delta = 69'sb111111111111111111111111111111111100000000000000001000000000000000000;
		22508: Delta = 69'sb000000000000000000000000000000000011111111111111111000000000000000000;
		12675: Delta = 69'sb111111111111111111111111111111111011111111111111111000000000000000000;
		17672: Delta = 69'sb000000000000000000000000000000001000000000000000001000000000000000000;
		48867: Delta = 69'sb111111111111111111111111111111111000000000000000001000000000000000000;
		1994: Delta = 69'sb000000000000000000000000000000000111111111111111111000000000000000000;
		33189: Delta = 69'sb111111111111111111111111111111110111111111111111111000000000000000000;
		27505: Delta = 69'sb000000000000000000000000000000010000000000000000001000000000000000000;
		39034: Delta = 69'sb111111111111111111111111111111110000000000000000001000000000000000000;
		11827: Delta = 69'sb000000000000000000000000000000001111111111111111111000000000000000000;
		23356: Delta = 69'sb111111111111111111111111111111101111111111111111111000000000000000000;
		47171: Delta = 69'sb000000000000000000000000000000100000000000000000001000000000000000000;
		19368: Delta = 69'sb111111111111111111111111111111100000000000000000001000000000000000000;
		31493: Delta = 69'sb000000000000000000000000000000011111111111111111111000000000000000000;
		3690: Delta = 69'sb111111111111111111111111111111011111111111111111111000000000000000000;
		35642: Delta = 69'sb000000000000000000000000000001000000000000000000001000000000000000000;
		30897: Delta = 69'sb111111111111111111111111111111000000000000000000001000000000000000000;
		19964: Delta = 69'sb000000000000000000000000000000111111111111111111111000000000000000000;
		15219: Delta = 69'sb111111111111111111111111111110111111111111111111111000000000000000000;
		12584: Delta = 69'sb000000000000000000000000000010000000000000000000001000000000000000000;
		3094: Delta = 69'sb111111111111111111111111111110000000000000000000001000000000000000000;
		47767: Delta = 69'sb000000000000000000000000000001111111111111111111111000000000000000000;
		38277: Delta = 69'sb111111111111111111111111111101111111111111111111111000000000000000000;
		17329: Delta = 69'sb000000000000000000000000000100000000000000000000001000000000000000000;
		49210: Delta = 69'sb111111111111111111111111111100000000000000000000001000000000000000000;
		1651: Delta = 69'sb000000000000000000000000000011111111111111111111111000000000000000000;
		33532: Delta = 69'sb111111111111111111111111111011111111111111111111111000000000000000000;
		26819: Delta = 69'sb000000000000000000000000001000000000000000000000001000000000000000000;
		39720: Delta = 69'sb111111111111111111111111111000000000000000000000001000000000000000000;
		11141: Delta = 69'sb000000000000000000000000000111111111111111111111111000000000000000000;
		24042: Delta = 69'sb111111111111111111111111110111111111111111111111111000000000000000000;
		45799: Delta = 69'sb000000000000000000000000010000000000000000000000001000000000000000000;
		20740: Delta = 69'sb111111111111111111111111110000000000000000000000001000000000000000000;
		30121: Delta = 69'sb000000000000000000000000001111111111111111111111111000000000000000000;
		5062: Delta = 69'sb111111111111111111111111101111111111111111111111111000000000000000000;
		32898: Delta = 69'sb000000000000000000000000100000000000000000000000001000000000000000000;
		33641: Delta = 69'sb111111111111111111111111100000000000000000000000001000000000000000000;
		17220: Delta = 69'sb000000000000000000000000011111111111111111111111111000000000000000000;
		17963: Delta = 69'sb111111111111111111111111011111111111111111111111111000000000000000000;
		7096: Delta = 69'sb000000000000000000000001000000000000000000000000001000000000000000000;
		8582: Delta = 69'sb111111111111111111111111000000000000000000000000001000000000000000000;
		42279: Delta = 69'sb000000000000000000000000111111111111111111111111111000000000000000000;
		43765: Delta = 69'sb111111111111111111111110111111111111111111111111111000000000000000000;
		6353: Delta = 69'sb000000000000000000000010000000000000000000000000001000000000000000000;
		9325: Delta = 69'sb111111111111111111111110000000000000000000000000001000000000000000000;
		41536: Delta = 69'sb000000000000000000000001111111111111111111111111111000000000000000000;
		44508: Delta = 69'sb111111111111111111111101111111111111111111111111111000000000000000000;
		4867: Delta = 69'sb000000000000000000000100000000000000000000000000001000000000000000000;
		10811: Delta = 69'sb111111111111111111111100000000000000000000000000001000000000000000000;
		40050: Delta = 69'sb000000000000000000000011111111111111111111111111111000000000000000000;
		45994: Delta = 69'sb111111111111111111111011111111111111111111111111111000000000000000000;
		1895: Delta = 69'sb000000000000000000001000000000000000000000000000001000000000000000000;
		13783: Delta = 69'sb111111111111111111111000000000000000000000000000001000000000000000000;
		37078: Delta = 69'sb000000000000000000000111111111111111111111111111111000000000000000000;
		48966: Delta = 69'sb111111111111111111110111111111111111111111111111111000000000000000000;
		46812: Delta = 69'sb000000000000000000010000000000000000000000000000001000000000000000000;
		19727: Delta = 69'sb111111111111111111110000000000000000000000000000001000000000000000000;
		31134: Delta = 69'sb000000000000000000001111111111111111111111111111111000000000000000000;
		4049: Delta = 69'sb111111111111111111101111111111111111111111111111111000000000000000000;
		34924: Delta = 69'sb000000000000000000100000000000000000000000000000001000000000000000000;
		31615: Delta = 69'sb111111111111111111100000000000000000000000000000001000000000000000000;
		19246: Delta = 69'sb000000000000000000011111111111111111111111111111111000000000000000000;
		15937: Delta = 69'sb111111111111111111011111111111111111111111111111111000000000000000000;
		11148: Delta = 69'sb000000000000000001000000000000000000000000000000001000000000000000000;
		4530: Delta = 69'sb111111111111111111000000000000000000000000000000001000000000000000000;
		46331: Delta = 69'sb000000000000000000111111111111111111111111111111111000000000000000000;
		39713: Delta = 69'sb111111111111111110111111111111111111111111111111111000000000000000000;
		14457: Delta = 69'sb000000000000000010000000000000000000000000000000001000000000000000000;
		1221: Delta = 69'sb111111111111111110000000000000000000000000000000001000000000000000000;
		49640: Delta = 69'sb000000000000000001111111111111111111111111111111111000000000000000000;
		36404: Delta = 69'sb111111111111111101111111111111111111111111111111111000000000000000000;
		21075: Delta = 69'sb000000000000000100000000000000000000000000000000001000000000000000000;
		45464: Delta = 69'sb111111111111111100000000000000000000000000000000001000000000000000000;
		5397: Delta = 69'sb000000000000000011111111111111111111111111111111111000000000000000000;
		29786: Delta = 69'sb111111111111111011111111111111111111111111111111111000000000000000000;
		34311: Delta = 69'sb000000000000001000000000000000000000000000000000001000000000000000000;
		32228: Delta = 69'sb111111111111111000000000000000000000000000000000001000000000000000000;
		18633: Delta = 69'sb000000000000000111111111111111111111111111111111111000000000000000000;
		16550: Delta = 69'sb111111111111110111111111111111111111111111111111111000000000000000000;
		9922: Delta = 69'sb000000000000010000000000000000000000000000000000001000000000000000000;
		5756: Delta = 69'sb111111111111110000000000000000000000000000000000001000000000000000000;
		45105: Delta = 69'sb000000000000001111111111111111111111111111111111111000000000000000000;
		40939: Delta = 69'sb111111111111101111111111111111111111111111111111111000000000000000000;
		12005: Delta = 69'sb000000000000100000000000000000000000000000000000001000000000000000000;
		3673: Delta = 69'sb111111111111100000000000000000000000000000000000001000000000000000000;
		47188: Delta = 69'sb000000000000011111111111111111111111111111111111111000000000000000000;
		38856: Delta = 69'sb111111111111011111111111111111111111111111111111111000000000000000000;
		16171: Delta = 69'sb000000000001000000000000000000000000000000000000001000000000000000000;
		50368: Delta = 69'sb111111111111000000000000000000000000000000000000001000000000000000000;
		493: Delta = 69'sb000000000000111111111111111111111111111111111111111000000000000000000;
		34690: Delta = 69'sb111111111110111111111111111111111111111111111111111000000000000000000;
		24503: Delta = 69'sb000000000010000000000000000000000000000000000000001000000000000000000;
		42036: Delta = 69'sb111111111110000000000000000000000000000000000000001000000000000000000;
		8825: Delta = 69'sb000000000001111111111111111111111111111111111111111000000000000000000;
		26358: Delta = 69'sb111111111101111111111111111111111111111111111111111000000000000000000;
		41167: Delta = 69'sb000000000100000000000000000000000000000000000000001000000000000000000;
		25372: Delta = 69'sb111111111100000000000000000000000000000000000000001000000000000000000;
		25489: Delta = 69'sb000000000011111111111111111111111111111111111111111000000000000000000;
		9694: Delta = 69'sb111111111011111111111111111111111111111111111111111000000000000000000;
		23634: Delta = 69'sb000000001000000000000000000000000000000000000000001000000000000000000;
		42905: Delta = 69'sb111111111000000000000000000000000000000000000000001000000000000000000;
		7956: Delta = 69'sb000000000111111111111111111111111111111111111111111000000000000000000;
		27227: Delta = 69'sb111111110111111111111111111111111111111111111111111000000000000000000;
		39429: Delta = 69'sb000000010000000000000000000000000000000000000000001000000000000000000;
		27110: Delta = 69'sb111111110000000000000000000000000000000000000000001000000000000000000;
		23751: Delta = 69'sb000000001111111111111111111111111111111111111111111000000000000000000;
		11432: Delta = 69'sb111111101111111111111111111111111111111111111111111000000000000000000;
		20158: Delta = 69'sb000000100000000000000000000000000000000000000000001000000000000000000;
		46381: Delta = 69'sb111111100000000000000000000000000000000000000000001000000000000000000;
		4480: Delta = 69'sb000000011111111111111111111111111111111111111111111000000000000000000;
		30703: Delta = 69'sb111111011111111111111111111111111111111111111111111000000000000000000;
		32477: Delta = 69'sb000001000000000000000000000000000000000000000000001000000000000000000;
		34062: Delta = 69'sb111111000000000000000000000000000000000000000000001000000000000000000;
		16799: Delta = 69'sb000000111111111111111111111111111111111111111111111000000000000000000;
		18384: Delta = 69'sb111110111111111111111111111111111111111111111111111000000000000000000;
		6254: Delta = 69'sb000010000000000000000000000000000000000000000000001000000000000000000;
		9424: Delta = 69'sb111110000000000000000000000000000000000000000000001000000000000000000;
		41437: Delta = 69'sb000001111111111111111111111111111111111111111111111000000000000000000;
		44607: Delta = 69'sb111101111111111111111111111111111111111111111111111000000000000000000;
		4669: Delta = 69'sb000100000000000000000000000000000000000000000000001000000000000000000;
		11009: Delta = 69'sb111100000000000000000000000000000000000000000000001000000000000000000;
		39852: Delta = 69'sb000011111111111111111111111111111111111111111111111000000000000000000;
		46192: Delta = 69'sb111011111111111111111111111111111111111111111111111000000000000000000;
		1499: Delta = 69'sb001000000000000000000000000000000000000000000000001000000000000000000;
		14179: Delta = 69'sb111000000000000000000000000000000000000000000000001000000000000000000;
		36682: Delta = 69'sb000111111111111111111111111111111111111111111111111000000000000000000;
		49362: Delta = 69'sb110111111111111111111111111111111111111111111111111000000000000000000;
		46020: Delta = 69'sb010000000000000000000000000000000000000000000000001000000000000000000;
		20519: Delta = 69'sb110000000000000000000000000000000000000000000000001000000000000000000;
		30342: Delta = 69'sb001111111111111111111111111111111111111111111111111000000000000000000;
		4841: Delta = 69'sb101111111111111111111111111111111111111111111111111000000000000000000;
		47034: Delta = 69'sb000000000000000000000000000000000000000000000000110000000000000000000;
		3827: Delta = 69'sb111111111111111111111111111111111111111111111111010000000000000000000;
		27529: Delta = 69'sb000000000000000000000000000000000000000000000001010000000000000000000;
		23332: Delta = 69'sb111111111111111111111111111111111111111111111110110000000000000000000;
		39380: Delta = 69'sb000000000000000000000000000000000000000000000010010000000000000000000;
		42837: Delta = 69'sb111111111111111111111111111111111111111111111110010000000000000000000;
		8024: Delta = 69'sb000000000000000000000000000000000000000000000001110000000000000000000;
		11481: Delta = 69'sb111111111111111111111111111111111111111111111101110000000000000000000;
		12221: Delta = 69'sb000000000000000000000000000000000000000000000100010000000000000000000;
		19135: Delta = 69'sb111111111111111111111111111111111111111111111100010000000000000000000;
		31726: Delta = 69'sb000000000000000000000000000000000000000000000011110000000000000000000;
		38640: Delta = 69'sb111111111111111111111111111111111111111111111011110000000000000000000;
		8764: Delta = 69'sb000000000000000000000000000000000000000000001000010000000000000000000;
		22592: Delta = 69'sb111111111111111111111111111111111111111111111000010000000000000000000;
		28269: Delta = 69'sb000000000000000000000000000000000000000000000111110000000000000000000;
		42097: Delta = 69'sb111111111111111111111111111111111111111111110111110000000000000000000;
		1850: Delta = 69'sb000000000000000000000000000000000000000000010000010000000000000000000;
		29506: Delta = 69'sb111111111111111111111111111111111111111111110000010000000000000000000;
		21355: Delta = 69'sb000000000000000000000000000000000000000000001111110000000000000000000;
		49011: Delta = 69'sb111111111111111111111111111111111111111111101111110000000000000000000;
		38883: Delta = 69'sb000000000000000000000000000000000000000000100000010000000000000000000;
		43334: Delta = 69'sb111111111111111111111111111111111111111111100000010000000000000000000;
		7527: Delta = 69'sb000000000000000000000000000000000000000000011111110000000000000000000;
		11978: Delta = 69'sb111111111111111111111111111111111111111111011111110000000000000000000;
		11227: Delta = 69'sb000000000000000000000000000000000000000001000000010000000000000000000;
		20129: Delta = 69'sb111111111111111111111111111111111111111111000000010000000000000000000;
		30732: Delta = 69'sb000000000000000000000000000000000000000000111111110000000000000000000;
		39634: Delta = 69'sb111111111111111111111111111111111111111110111111110000000000000000000;
		6776: Delta = 69'sb000000000000000000000000000000000000000010000000010000000000000000000;
		24580: Delta = 69'sb111111111111111111111111111111111111111110000000010000000000000000000;
		26281: Delta = 69'sb000000000000000000000000000000000000000001111111110000000000000000000;
		44085: Delta = 69'sb111111111111111111111111111111111111111101111111110000000000000000000;
		48735: Delta = 69'sb000000000000000000000000000000000000000100000000010000000000000000000;
		33482: Delta = 69'sb111111111111111111111111111111111111111100000000010000000000000000000;
		17379: Delta = 69'sb000000000000000000000000000000000000000011111111110000000000000000000;
		2126: Delta = 69'sb111111111111111111111111111111111111111011111111110000000000000000000;
		30931: Delta = 69'sb000000000000000000000000000000000000001000000000010000000000000000000;
		425: Delta = 69'sb111111111111111111111111111111111111111000000000010000000000000000000;
		50436: Delta = 69'sb000000000000000000000000000000000000000111111111110000000000000000000;
		19930: Delta = 69'sb111111111111111111111111111111111111110111111111110000000000000000000;
		46184: Delta = 69'sb000000000000000000000000000000000000010000000000010000000000000000000;
		36033: Delta = 69'sb111111111111111111111111111111111111110000000000010000000000000000000;
		14828: Delta = 69'sb000000000000000000000000000000000000001111111111110000000000000000000;
		4677: Delta = 69'sb111111111111111111111111111111111111101111111111110000000000000000000;
		25829: Delta = 69'sb000000000000000000000000000000000000100000000000010000000000000000000;
		5527: Delta = 69'sb111111111111111111111111111111111111100000000000010000000000000000000;
		45334: Delta = 69'sb000000000000000000000000000000000000011111111111110000000000000000000;
		25032: Delta = 69'sb111111111111111111111111111111111111011111111111110000000000000000000;
		35980: Delta = 69'sb000000000000000000000000000000000001000000000000010000000000000000000;
		46237: Delta = 69'sb111111111111111111111111111111111111000000000000010000000000000000000;
		4624: Delta = 69'sb000000000000000000000000000000000000111111111111110000000000000000000;
		14881: Delta = 69'sb111111111111111111111111111111111110111111111111110000000000000000000;
		5421: Delta = 69'sb000000000000000000000000000000000010000000000000010000000000000000000;
		25935: Delta = 69'sb111111111111111111111111111111111110000000000000010000000000000000000;
		24926: Delta = 69'sb000000000000000000000000000000000001111111111111110000000000000000000;
		45440: Delta = 69'sb111111111111111111111111111111111101111111111111110000000000000000000;
		46025: Delta = 69'sb000000000000000000000000000000000100000000000000010000000000000000000;
		36192: Delta = 69'sb111111111111111111111111111111111100000000000000010000000000000000000;
		14669: Delta = 69'sb000000000000000000000000000000000011111111111111110000000000000000000;
		4836: Delta = 69'sb111111111111111111111111111111111011111111111111110000000000000000000;
		25511: Delta = 69'sb000000000000000000000000000000001000000000000000010000000000000000000;
		5845: Delta = 69'sb111111111111111111111111111111111000000000000000010000000000000000000;
		45016: Delta = 69'sb000000000000000000000000000000000111111111111111110000000000000000000;
		25350: Delta = 69'sb111111111111111111111111111111110111111111111111110000000000000000000;
		35344: Delta = 69'sb000000000000000000000000000000010000000000000000010000000000000000000;
		46873: Delta = 69'sb111111111111111111111111111111110000000000000000010000000000000000000;
		3988: Delta = 69'sb000000000000000000000000000000001111111111111111110000000000000000000;
		15517: Delta = 69'sb111111111111111111111111111111101111111111111111110000000000000000000;
		4149: Delta = 69'sb000000000000000000000000000000100000000000000000010000000000000000000;
		27207: Delta = 69'sb111111111111111111111111111111100000000000000000010000000000000000000;
		23654: Delta = 69'sb000000000000000000000000000000011111111111111111110000000000000000000;
		46712: Delta = 69'sb111111111111111111111111111111011111111111111111110000000000000000000;
		43481: Delta = 69'sb000000000000000000000000000001000000000000000000010000000000000000000;
		38736: Delta = 69'sb111111111111111111111111111111000000000000000000010000000000000000000;
		12125: Delta = 69'sb000000000000000000000000000000111111111111111111110000000000000000000;
		7380: Delta = 69'sb111111111111111111111111111110111111111111111111110000000000000000000;
		20423: Delta = 69'sb000000000000000000000000000010000000000000000000010000000000000000000;
		10933: Delta = 69'sb111111111111111111111111111110000000000000000000010000000000000000000;
		39928: Delta = 69'sb000000000000000000000000000001111111111111111111110000000000000000000;
		30438: Delta = 69'sb111111111111111111111111111101111111111111111111110000000000000000000;
		25168: Delta = 69'sb000000000000000000000000000100000000000000000000010000000000000000000;
		6188: Delta = 69'sb111111111111111111111111111100000000000000000000010000000000000000000;
		44673: Delta = 69'sb000000000000000000000000000011111111111111111111110000000000000000000;
		25693: Delta = 69'sb111111111111111111111111111011111111111111111111110000000000000000000;
		34658: Delta = 69'sb000000000000000000000000001000000000000000000000010000000000000000000;
		47559: Delta = 69'sb111111111111111111111111111000000000000000000000010000000000000000000;
		3302: Delta = 69'sb000000000000000000000000000111111111111111111111110000000000000000000;
		16203: Delta = 69'sb111111111111111111111111110111111111111111111111110000000000000000000;
		2777: Delta = 69'sb000000000000000000000000010000000000000000000000010000000000000000000;
		28579: Delta = 69'sb111111111111111111111111110000000000000000000000010000000000000000000;
		22282: Delta = 69'sb000000000000000000000000001111111111111111111111110000000000000000000;
		48084: Delta = 69'sb111111111111111111111111101111111111111111111111110000000000000000000;
		40737: Delta = 69'sb000000000000000000000000100000000000000000000000010000000000000000000;
		41480: Delta = 69'sb111111111111111111111111100000000000000000000000010000000000000000000;
		9381: Delta = 69'sb000000000000000000000000011111111111111111111111110000000000000000000;
		10124: Delta = 69'sb111111111111111111111111011111111111111111111111110000000000000000000;
		14935: Delta = 69'sb000000000000000000000001000000000000000000000000010000000000000000000;
		16421: Delta = 69'sb111111111111111111111111000000000000000000000000010000000000000000000;
		34440: Delta = 69'sb000000000000000000000000111111111111111111111111110000000000000000000;
		35926: Delta = 69'sb111111111111111111111110111111111111111111111111110000000000000000000;
		14192: Delta = 69'sb000000000000000000000010000000000000000000000000010000000000000000000;
		17164: Delta = 69'sb111111111111111111111110000000000000000000000000010000000000000000000;
		33697: Delta = 69'sb000000000000000000000001111111111111111111111111110000000000000000000;
		36669: Delta = 69'sb111111111111111111111101111111111111111111111111110000000000000000000;
		12706: Delta = 69'sb000000000000000000000100000000000000000000000000010000000000000000000;
		18650: Delta = 69'sb111111111111111111111100000000000000000000000000010000000000000000000;
		32211: Delta = 69'sb000000000000000000000011111111111111111111111111110000000000000000000;
		38155: Delta = 69'sb111111111111111111111011111111111111111111111111110000000000000000000;
		9734: Delta = 69'sb000000000000000000001000000000000000000000000000010000000000000000000;
		21622: Delta = 69'sb111111111111111111111000000000000000000000000000010000000000000000000;
		29239: Delta = 69'sb000000000000000000000111111111111111111111111111110000000000000000000;
		41127: Delta = 69'sb111111111111111111110111111111111111111111111111110000000000000000000;
		3790: Delta = 69'sb000000000000000000010000000000000000000000000000010000000000000000000;
		27566: Delta = 69'sb111111111111111111110000000000000000000000000000010000000000000000000;
		23295: Delta = 69'sb000000000000000000001111111111111111111111111111110000000000000000000;
		47071: Delta = 69'sb111111111111111111101111111111111111111111111111110000000000000000000;
		42763: Delta = 69'sb000000000000000000100000000000000000000000000000010000000000000000000;
		39454: Delta = 69'sb111111111111111111100000000000000000000000000000010000000000000000000;
		11407: Delta = 69'sb000000000000000000011111111111111111111111111111110000000000000000000;
		8098: Delta = 69'sb111111111111111111011111111111111111111111111111110000000000000000000;
		18987: Delta = 69'sb000000000000000001000000000000000000000000000000010000000000000000000;
		12369: Delta = 69'sb111111111111111111000000000000000000000000000000010000000000000000000;
		38492: Delta = 69'sb000000000000000000111111111111111111111111111111110000000000000000000;
		31874: Delta = 69'sb111111111111111110111111111111111111111111111111110000000000000000000;
		22296: Delta = 69'sb000000000000000010000000000000000000000000000000010000000000000000000;
		9060: Delta = 69'sb111111111111111110000000000000000000000000000000010000000000000000000;
		41801: Delta = 69'sb000000000000000001111111111111111111111111111111110000000000000000000;
		28565: Delta = 69'sb111111111111111101111111111111111111111111111111110000000000000000000;
		28914: Delta = 69'sb000000000000000100000000000000000000000000000000010000000000000000000;
		2442: Delta = 69'sb111111111111111100000000000000000000000000000000010000000000000000000;
		48419: Delta = 69'sb000000000000000011111111111111111111111111111111110000000000000000000;
		21947: Delta = 69'sb111111111111111011111111111111111111111111111111110000000000000000000;
		42150: Delta = 69'sb000000000000001000000000000000000000000000000000010000000000000000000;
		40067: Delta = 69'sb111111111111111000000000000000000000000000000000010000000000000000000;
		10794: Delta = 69'sb000000000000000111111111111111111111111111111111110000000000000000000;
		8711: Delta = 69'sb111111111111110111111111111111111111111111111111110000000000000000000;
		17761: Delta = 69'sb000000000000010000000000000000000000000000000000010000000000000000000;
		13595: Delta = 69'sb111111111111110000000000000000000000000000000000010000000000000000000;
		37266: Delta = 69'sb000000000000001111111111111111111111111111111111110000000000000000000;
		33100: Delta = 69'sb111111111111101111111111111111111111111111111111110000000000000000000;
		19844: Delta = 69'sb000000000000100000000000000000000000000000000000010000000000000000000;
		11512: Delta = 69'sb111111111111100000000000000000000000000000000000010000000000000000000;
		39349: Delta = 69'sb000000000000011111111111111111111111111111111111110000000000000000000;
		31017: Delta = 69'sb111111111111011111111111111111111111111111111111110000000000000000000;
		24010: Delta = 69'sb000000000001000000000000000000000000000000000000010000000000000000000;
		7346: Delta = 69'sb111111111111000000000000000000000000000000000000010000000000000000000;
		43515: Delta = 69'sb000000000000111111111111111111111111111111111111110000000000000000000;
		26851: Delta = 69'sb111111111110111111111111111111111111111111111111110000000000000000000;
		32342: Delta = 69'sb000000000010000000000000000000000000000000000000010000000000000000000;
		49875: Delta = 69'sb111111111110000000000000000000000000000000000000010000000000000000000;
		986: Delta = 69'sb000000000001111111111111111111111111111111111111110000000000000000000;
		18519: Delta = 69'sb111111111101111111111111111111111111111111111111110000000000000000000;
		49006: Delta = 69'sb000000000100000000000000000000000000000000000000010000000000000000000;
		33211: Delta = 69'sb111111111100000000000000000000000000000000000000010000000000000000000;
		17650: Delta = 69'sb000000000011111111111111111111111111111111111111110000000000000000000;
		1855: Delta = 69'sb111111111011111111111111111111111111111111111111110000000000000000000;
		31473: Delta = 69'sb000000001000000000000000000000000000000000000000010000000000000000000;
		50744: Delta = 69'sb111111111000000000000000000000000000000000000000010000000000000000000;
		117: Delta = 69'sb000000000111111111111111111111111111111111111111110000000000000000000;
		19388: Delta = 69'sb111111110111111111111111111111111111111111111111110000000000000000000;
		47268: Delta = 69'sb000000010000000000000000000000000000000000000000010000000000000000000;
		34949: Delta = 69'sb111111110000000000000000000000000000000000000000010000000000000000000;
		15912: Delta = 69'sb000000001111111111111111111111111111111111111111110000000000000000000;
		3593: Delta = 69'sb111111101111111111111111111111111111111111111111110000000000000000000;
		27997: Delta = 69'sb000000100000000000000000000000000000000000000000010000000000000000000;
		3359: Delta = 69'sb111111100000000000000000000000000000000000000000010000000000000000000;
		47502: Delta = 69'sb000000011111111111111111111111111111111111111111110000000000000000000;
		22864: Delta = 69'sb111111011111111111111111111111111111111111111111110000000000000000000;
		40316: Delta = 69'sb000001000000000000000000000000000000000000000000010000000000000000000;
		41901: Delta = 69'sb111111000000000000000000000000000000000000000000010000000000000000000;
		8960: Delta = 69'sb000000111111111111111111111111111111111111111111110000000000000000000;
		10545: Delta = 69'sb111110111111111111111111111111111111111111111111110000000000000000000;
		14093: Delta = 69'sb000010000000000000000000000000000000000000000000010000000000000000000;
		17263: Delta = 69'sb111110000000000000000000000000000000000000000000010000000000000000000;
		33598: Delta = 69'sb000001111111111111111111111111111111111111111111110000000000000000000;
		36768: Delta = 69'sb111101111111111111111111111111111111111111111111110000000000000000000;
		12508: Delta = 69'sb000100000000000000000000000000000000000000000000010000000000000000000;
		18848: Delta = 69'sb111100000000000000000000000000000000000000000000010000000000000000000;
		32013: Delta = 69'sb000011111111111111111111111111111111111111111111110000000000000000000;
		38353: Delta = 69'sb111011111111111111111111111111111111111111111111110000000000000000000;
		9338: Delta = 69'sb001000000000000000000000000000000000000000000000010000000000000000000;
		22018: Delta = 69'sb111000000000000000000000000000000000000000000000010000000000000000000;
		28843: Delta = 69'sb000111111111111111111111111111111111111111111111110000000000000000000;
		41523: Delta = 69'sb110111111111111111111111111111111111111111111111110000000000000000000;
		2998: Delta = 69'sb010000000000000000000000000000000000000000000000010000000000000000000;
		28358: Delta = 69'sb110000000000000000000000000000000000000000000000010000000000000000000;
		22503: Delta = 69'sb001111111111111111111111111111111111111111111111110000000000000000000;
		47863: Delta = 69'sb101111111111111111111111111111111111111111111111110000000000000000000;
		43207: Delta = 69'sb000000000000000000000000000000000000000000000001100000000000000000000;
		7654: Delta = 69'sb111111111111111111111111111111111111111111111110100000000000000000000;
		4197: Delta = 69'sb000000000000000000000000000000000000000000000010100000000000000000000;
		46664: Delta = 69'sb111111111111111111111111111111111111111111111101100000000000000000000;
		27899: Delta = 69'sb000000000000000000000000000000000000000000000100100000000000000000000;
		34813: Delta = 69'sb111111111111111111111111111111111111111111111100100000000000000000000;
		16048: Delta = 69'sb000000000000000000000000000000000000000000000011100000000000000000000;
		22962: Delta = 69'sb111111111111111111111111111111111111111111111011100000000000000000000;
		24442: Delta = 69'sb000000000000000000000000000000000000000000001000100000000000000000000;
		38270: Delta = 69'sb111111111111111111111111111111111111111111111000100000000000000000000;
		12591: Delta = 69'sb000000000000000000000000000000000000000000000111100000000000000000000;
		26419: Delta = 69'sb111111111111111111111111111111111111111111110111100000000000000000000;
		17528: Delta = 69'sb000000000000000000000000000000000000000000010000100000000000000000000;
		45184: Delta = 69'sb111111111111111111111111111111111111111111110000100000000000000000000;
		5677: Delta = 69'sb000000000000000000000000000000000000000000001111100000000000000000000;
		33333: Delta = 69'sb111111111111111111111111111111111111111111101111100000000000000000000;
		3700: Delta = 69'sb000000000000000000000000000000000000000000100000100000000000000000000;
		8151: Delta = 69'sb111111111111111111111111111111111111111111100000100000000000000000000;
		42710: Delta = 69'sb000000000000000000000000000000000000000000011111100000000000000000000;
		47161: Delta = 69'sb111111111111111111111111111111111111111111011111100000000000000000000;
		26905: Delta = 69'sb000000000000000000000000000000000000000001000000100000000000000000000;
		35807: Delta = 69'sb111111111111111111111111111111111111111111000000100000000000000000000;
		15054: Delta = 69'sb000000000000000000000000000000000000000000111111100000000000000000000;
		23956: Delta = 69'sb111111111111111111111111111111111111111110111111100000000000000000000;
		22454: Delta = 69'sb000000000000000000000000000000000000000010000000100000000000000000000;
		40258: Delta = 69'sb111111111111111111111111111111111111111110000000100000000000000000000;
		10603: Delta = 69'sb000000000000000000000000000000000000000001111111100000000000000000000;
		28407: Delta = 69'sb111111111111111111111111111111111111111101111111100000000000000000000;
		13552: Delta = 69'sb000000000000000000000000000000000000000100000000100000000000000000000;
		49160: Delta = 69'sb111111111111111111111111111111111111111100000000100000000000000000000;
		1701: Delta = 69'sb000000000000000000000000000000000000000011111111100000000000000000000;
		37309: Delta = 69'sb111111111111111111111111111111111111111011111111100000000000000000000;
		46609: Delta = 69'sb000000000000000000000000000000000000001000000000100000000000000000000;
		16103: Delta = 69'sb111111111111111111111111111111111111111000000000100000000000000000000;
		34758: Delta = 69'sb000000000000000000000000000000000000000111111111100000000000000000000;
		4252: Delta = 69'sb111111111111111111111111111111111111110111111111100000000000000000000;
		11001: Delta = 69'sb000000000000000000000000000000000000010000000000100000000000000000000;
		850: Delta = 69'sb111111111111111111111111111111111111110000000000100000000000000000000;
		50011: Delta = 69'sb000000000000000000000000000000000000001111111111100000000000000000000;
		39860: Delta = 69'sb111111111111111111111111111111111111101111111111100000000000000000000;
		41507: Delta = 69'sb000000000000000000000000000000000000100000000000100000000000000000000;
		21205: Delta = 69'sb111111111111111111111111111111111111100000000000100000000000000000000;
		29656: Delta = 69'sb000000000000000000000000000000000000011111111111100000000000000000000;
		9354: Delta = 69'sb111111111111111111111111111111111111011111111111100000000000000000000;
		797: Delta = 69'sb000000000000000000000000000000000001000000000000100000000000000000000;
		11054: Delta = 69'sb111111111111111111111111111111111111000000000000100000000000000000000;
		39807: Delta = 69'sb000000000000000000000000000000000000111111111111100000000000000000000;
		50064: Delta = 69'sb111111111111111111111111111111111110111111111111100000000000000000000;
		21099: Delta = 69'sb000000000000000000000000000000000010000000000000100000000000000000000;
		41613: Delta = 69'sb111111111111111111111111111111111110000000000000100000000000000000000;
		9248: Delta = 69'sb000000000000000000000000000000000001111111111111100000000000000000000;
		29762: Delta = 69'sb111111111111111111111111111111111101111111111111100000000000000000000;
		10842: Delta = 69'sb000000000000000000000000000000000100000000000000100000000000000000000;
		1009: Delta = 69'sb111111111111111111111111111111111100000000000000100000000000000000000;
		49852: Delta = 69'sb000000000000000000000000000000000011111111111111100000000000000000000;
		40019: Delta = 69'sb111111111111111111111111111111111011111111111111100000000000000000000;
		41189: Delta = 69'sb000000000000000000000000000000001000000000000000100000000000000000000;
		21523: Delta = 69'sb111111111111111111111111111111111000000000000000100000000000000000000;
		29338: Delta = 69'sb000000000000000000000000000000000111111111111111100000000000000000000;
		9672: Delta = 69'sb111111111111111111111111111111110111111111111111100000000000000000000;
		161: Delta = 69'sb000000000000000000000000000000010000000000000000100000000000000000000;
		11690: Delta = 69'sb111111111111111111111111111111110000000000000000100000000000000000000;
		39171: Delta = 69'sb000000000000000000000000000000001111111111111111100000000000000000000;
		50700: Delta = 69'sb111111111111111111111111111111101111111111111111100000000000000000000;
		19827: Delta = 69'sb000000000000000000000000000000100000000000000000100000000000000000000;
		42885: Delta = 69'sb111111111111111111111111111111100000000000000000100000000000000000000;
		7976: Delta = 69'sb000000000000000000000000000000011111111111111111100000000000000000000;
		31034: Delta = 69'sb111111111111111111111111111111011111111111111111100000000000000000000;
		8298: Delta = 69'sb000000000000000000000000000001000000000000000000100000000000000000000;
		3553: Delta = 69'sb111111111111111111111111111111000000000000000000100000000000000000000;
		47308: Delta = 69'sb000000000000000000000000000000111111111111111111100000000000000000000;
		42563: Delta = 69'sb111111111111111111111111111110111111111111111111100000000000000000000;
		36101: Delta = 69'sb000000000000000000000000000010000000000000000000100000000000000000000;
		26611: Delta = 69'sb111111111111111111111111111110000000000000000000100000000000000000000;
		24250: Delta = 69'sb000000000000000000000000000001111111111111111111100000000000000000000;
		14760: Delta = 69'sb111111111111111111111111111101111111111111111111100000000000000000000;
		40846: Delta = 69'sb000000000000000000000000000100000000000000000000100000000000000000000;
		21866: Delta = 69'sb111111111111111111111111111100000000000000000000100000000000000000000;
		28995: Delta = 69'sb000000000000000000000000000011111111111111111111100000000000000000000;
		10015: Delta = 69'sb111111111111111111111111111011111111111111111111100000000000000000000;
		50336: Delta = 69'sb000000000000000000000000001000000000000000000000100000000000000000000;
		12376: Delta = 69'sb111111111111111111111111111000000000000000000000100000000000000000000;
		38485: Delta = 69'sb000000000000000000000000000111111111111111111111100000000000000000000;
		525: Delta = 69'sb111111111111111111111111110111111111111111111111100000000000000000000;
		18455: Delta = 69'sb000000000000000000000000010000000000000000000000100000000000000000000;
		44257: Delta = 69'sb111111111111111111111111110000000000000000000000100000000000000000000;
		6604: Delta = 69'sb000000000000000000000000001111111111111111111111100000000000000000000;
		32406: Delta = 69'sb111111111111111111111111101111111111111111111111100000000000000000000;
		5554: Delta = 69'sb000000000000000000000000100000000000000000000000100000000000000000000;
		6297: Delta = 69'sb111111111111111111111111100000000000000000000000100000000000000000000;
		44564: Delta = 69'sb000000000000000000000000011111111111111111111111100000000000000000000;
		45307: Delta = 69'sb111111111111111111111111011111111111111111111111100000000000000000000;
		30613: Delta = 69'sb000000000000000000000001000000000000000000000000100000000000000000000;
		32099: Delta = 69'sb111111111111111111111111000000000000000000000000100000000000000000000;
		18762: Delta = 69'sb000000000000000000000000111111111111111111111111100000000000000000000;
		20248: Delta = 69'sb111111111111111111111110111111111111111111111111100000000000000000000;
		29870: Delta = 69'sb000000000000000000000010000000000000000000000000100000000000000000000;
		32842: Delta = 69'sb111111111111111111111110000000000000000000000000100000000000000000000;
		18019: Delta = 69'sb000000000000000000000001111111111111111111111111100000000000000000000;
		20991: Delta = 69'sb111111111111111111111101111111111111111111111111100000000000000000000;
		28384: Delta = 69'sb000000000000000000000100000000000000000000000000100000000000000000000;
		34328: Delta = 69'sb111111111111111111111100000000000000000000000000100000000000000000000;
		16533: Delta = 69'sb000000000000000000000011111111111111111111111111100000000000000000000;
		22477: Delta = 69'sb111111111111111111111011111111111111111111111111100000000000000000000;
		25412: Delta = 69'sb000000000000000000001000000000000000000000000000100000000000000000000;
		37300: Delta = 69'sb111111111111111111111000000000000000000000000000100000000000000000000;
		13561: Delta = 69'sb000000000000000000000111111111111111111111111111100000000000000000000;
		25449: Delta = 69'sb111111111111111111110111111111111111111111111111100000000000000000000;
		19468: Delta = 69'sb000000000000000000010000000000000000000000000000100000000000000000000;
		43244: Delta = 69'sb111111111111111111110000000000000000000000000000100000000000000000000;
		7617: Delta = 69'sb000000000000000000001111111111111111111111111111100000000000000000000;
		31393: Delta = 69'sb111111111111111111101111111111111111111111111111100000000000000000000;
		7580: Delta = 69'sb000000000000000000100000000000000000000000000000100000000000000000000;
		4271: Delta = 69'sb111111111111111111100000000000000000000000000000100000000000000000000;
		46590: Delta = 69'sb000000000000000000011111111111111111111111111111100000000000000000000;
		43281: Delta = 69'sb111111111111111111011111111111111111111111111111100000000000000000000;
		34665: Delta = 69'sb000000000000000001000000000000000000000000000000100000000000000000000;
		28047: Delta = 69'sb111111111111111111000000000000000000000000000000100000000000000000000;
		22814: Delta = 69'sb000000000000000000111111111111111111111111111111100000000000000000000;
		16196: Delta = 69'sb111111111111111110111111111111111111111111111111100000000000000000000;
		37974: Delta = 69'sb000000000000000010000000000000000000000000000000100000000000000000000;
		24738: Delta = 69'sb111111111111111110000000000000000000000000000000100000000000000000000;
		26123: Delta = 69'sb000000000000000001111111111111111111111111111111100000000000000000000;
		12887: Delta = 69'sb111111111111111101111111111111111111111111111111100000000000000000000;
		44592: Delta = 69'sb000000000000000100000000000000000000000000000000100000000000000000000;
		18120: Delta = 69'sb111111111111111100000000000000000000000000000000100000000000000000000;
		32741: Delta = 69'sb000000000000000011111111111111111111111111111111100000000000000000000;
		6269: Delta = 69'sb111111111111111011111111111111111111111111111111100000000000000000000;
		6967: Delta = 69'sb000000000000001000000000000000000000000000000000100000000000000000000;
		4884: Delta = 69'sb111111111111111000000000000000000000000000000000100000000000000000000;
		45977: Delta = 69'sb000000000000000111111111111111111111111111111111100000000000000000000;
		43894: Delta = 69'sb111111111111110111111111111111111111111111111111100000000000000000000;
		33439: Delta = 69'sb000000000000010000000000000000000000000000000000100000000000000000000;
		29273: Delta = 69'sb111111111111110000000000000000000000000000000000100000000000000000000;
		21588: Delta = 69'sb000000000000001111111111111111111111111111111111100000000000000000000;
		17422: Delta = 69'sb111111111111101111111111111111111111111111111111100000000000000000000;
		35522: Delta = 69'sb000000000000100000000000000000000000000000000000100000000000000000000;
		27190: Delta = 69'sb111111111111100000000000000000000000000000000000100000000000000000000;
		23671: Delta = 69'sb000000000000011111111111111111111111111111111111100000000000000000000;
		15339: Delta = 69'sb111111111111011111111111111111111111111111111111100000000000000000000;
		39688: Delta = 69'sb000000000001000000000000000000000000000000000000100000000000000000000;
		23024: Delta = 69'sb111111111111000000000000000000000000000000000000100000000000000000000;
		27837: Delta = 69'sb000000000000111111111111111111111111111111111111100000000000000000000;
		11173: Delta = 69'sb111111111110111111111111111111111111111111111111100000000000000000000;
		48020: Delta = 69'sb000000000010000000000000000000000000000000000000100000000000000000000;
		14692: Delta = 69'sb111111111110000000000000000000000000000000000000100000000000000000000;
		36169: Delta = 69'sb000000000001111111111111111111111111111111111111100000000000000000000;
		2841: Delta = 69'sb111111111101111111111111111111111111111111111111100000000000000000000;
		13823: Delta = 69'sb000000000100000000000000000000000000000000000000100000000000000000000;
		48889: Delta = 69'sb111111111100000000000000000000000000000000000000100000000000000000000;
		1972: Delta = 69'sb000000000011111111111111111111111111111111111111100000000000000000000;
		37038: Delta = 69'sb111111111011111111111111111111111111111111111111100000000000000000000;
		47151: Delta = 69'sb000000001000000000000000000000000000000000000000100000000000000000000;
		15561: Delta = 69'sb111111111000000000000000000000000000000000000000100000000000000000000;
		35300: Delta = 69'sb000000000111111111111111111111111111111111111111100000000000000000000;
		3710: Delta = 69'sb111111110111111111111111111111111111111111111111100000000000000000000;
		12085: Delta = 69'sb000000010000000000000000000000000000000000000000100000000000000000000;
		50627: Delta = 69'sb111111110000000000000000000000000000000000000000100000000000000000000;
		234: Delta = 69'sb000000001111111111111111111111111111111111111111100000000000000000000;
		38776: Delta = 69'sb111111101111111111111111111111111111111111111111100000000000000000000;
		43675: Delta = 69'sb000000100000000000000000000000000000000000000000100000000000000000000;
		19037: Delta = 69'sb111111100000000000000000000000000000000000000000100000000000000000000;
		31824: Delta = 69'sb000000011111111111111111111111111111111111111111100000000000000000000;
		7186: Delta = 69'sb111111011111111111111111111111111111111111111111100000000000000000000;
		5133: Delta = 69'sb000001000000000000000000000000000000000000000000100000000000000000000;
		6718: Delta = 69'sb111111000000000000000000000000000000000000000000100000000000000000000;
		44143: Delta = 69'sb000000111111111111111111111111111111111111111111100000000000000000000;
		45728: Delta = 69'sb111110111111111111111111111111111111111111111111100000000000000000000;
		29771: Delta = 69'sb000010000000000000000000000000000000000000000000100000000000000000000;
		32941: Delta = 69'sb111110000000000000000000000000000000000000000000100000000000000000000;
		17920: Delta = 69'sb000001111111111111111111111111111111111111111111100000000000000000000;
		21090: Delta = 69'sb111101111111111111111111111111111111111111111111100000000000000000000;
		28186: Delta = 69'sb000100000000000000000000000000000000000000000000100000000000000000000;
		34526: Delta = 69'sb111100000000000000000000000000000000000000000000100000000000000000000;
		16335: Delta = 69'sb000011111111111111111111111111111111111111111111100000000000000000000;
		22675: Delta = 69'sb111011111111111111111111111111111111111111111111100000000000000000000;
		25016: Delta = 69'sb001000000000000000000000000000000000000000000000100000000000000000000;
		37696: Delta = 69'sb111000000000000000000000000000000000000000000000100000000000000000000;
		13165: Delta = 69'sb000111111111111111111111111111111111111111111111100000000000000000000;
		25845: Delta = 69'sb110111111111111111111111111111111111111111111111100000000000000000000;
		18676: Delta = 69'sb010000000000000000000000000000000000000000000000100000000000000000000;
		44036: Delta = 69'sb110000000000000000000000000000000000000000000000100000000000000000000;
		6825: Delta = 69'sb001111111111111111111111111111111111111111111111100000000000000000000;
		32185: Delta = 69'sb101111111111111111111111111111111111111111111111100000000000000000000;
		35553: Delta = 69'sb000000000000000000000000000000000000000000000011000000000000000000000;
		15308: Delta = 69'sb111111111111111111111111111111111111111111111101000000000000000000000;
		8394: Delta = 69'sb000000000000000000000000000000000000000000000101000000000000000000000;
		42467: Delta = 69'sb111111111111111111111111111111111111111111111011000000000000000000000;
		4937: Delta = 69'sb000000000000000000000000000000000000000000001001000000000000000000000;
		18765: Delta = 69'sb111111111111111111111111111111111111111111111001000000000000000000000;
		32096: Delta = 69'sb000000000000000000000000000000000000000000000111000000000000000000000;
		45924: Delta = 69'sb111111111111111111111111111111111111111111110111000000000000000000000;
		48884: Delta = 69'sb000000000000000000000000000000000000000000010001000000000000000000000;
		25679: Delta = 69'sb111111111111111111111111111111111111111111110001000000000000000000000;
		25182: Delta = 69'sb000000000000000000000000000000000000000000001111000000000000000000000;
		1977: Delta = 69'sb111111111111111111111111111111111111111111101111000000000000000000000;
		35056: Delta = 69'sb000000000000000000000000000000000000000000100001000000000000000000000;
		39507: Delta = 69'sb111111111111111111111111111111111111111111100001000000000000000000000;
		11354: Delta = 69'sb000000000000000000000000000000000000000000011111000000000000000000000;
		15805: Delta = 69'sb111111111111111111111111111111111111111111011111000000000000000000000;
		7400: Delta = 69'sb000000000000000000000000000000000000000001000001000000000000000000000;
		16302: Delta = 69'sb111111111111111111111111111111111111111111000001000000000000000000000;
		34559: Delta = 69'sb000000000000000000000000000000000000000000111111000000000000000000000;
		43461: Delta = 69'sb111111111111111111111111111111111111111110111111000000000000000000000;
		2949: Delta = 69'sb000000000000000000000000000000000000000010000001000000000000000000000;
		20753: Delta = 69'sb111111111111111111111111111111111111111110000001000000000000000000000;
		30108: Delta = 69'sb000000000000000000000000000000000000000001111111000000000000000000000;
		47912: Delta = 69'sb111111111111111111111111111111111111111101111111000000000000000000000;
		44908: Delta = 69'sb000000000000000000000000000000000000000100000001000000000000000000000;
		29655: Delta = 69'sb111111111111111111111111111111111111111100000001000000000000000000000;
		21206: Delta = 69'sb000000000000000000000000000000000000000011111111000000000000000000000;
		5953: Delta = 69'sb111111111111111111111111111111111111111011111111000000000000000000000;
		27104: Delta = 69'sb000000000000000000000000000000000000001000000001000000000000000000000;
		47459: Delta = 69'sb111111111111111111111111111111111111111000000001000000000000000000000;
		3402: Delta = 69'sb000000000000000000000000000000000000000111111111000000000000000000000;
		23757: Delta = 69'sb111111111111111111111111111111111111110111111111000000000000000000000;
		42357: Delta = 69'sb000000000000000000000000000000000000010000000001000000000000000000000;
		32206: Delta = 69'sb111111111111111111111111111111111111110000000001000000000000000000000;
		18655: Delta = 69'sb000000000000000000000000000000000000001111111111000000000000000000000;
		8504: Delta = 69'sb111111111111111111111111111111111111101111111111000000000000000000000;
		22002: Delta = 69'sb000000000000000000000000000000000000100000000001000000000000000000000;
		1700: Delta = 69'sb111111111111111111111111111111111111100000000001000000000000000000000;
		49161: Delta = 69'sb000000000000000000000000000000000000011111111111000000000000000000000;
		28859: Delta = 69'sb111111111111111111111111111111111111011111111111000000000000000000000;
		32153: Delta = 69'sb000000000000000000000000000000000001000000000001000000000000000000000;
		42410: Delta = 69'sb111111111111111111111111111111111111000000000001000000000000000000000;
		8451: Delta = 69'sb000000000000000000000000000000000000111111111111000000000000000000000;
		18708: Delta = 69'sb111111111111111111111111111111111110111111111111000000000000000000000;
		1594: Delta = 69'sb000000000000000000000000000000000010000000000001000000000000000000000;
		22108: Delta = 69'sb111111111111111111111111111111111110000000000001000000000000000000000;
		28753: Delta = 69'sb000000000000000000000000000000000001111111111111000000000000000000000;
		49267: Delta = 69'sb111111111111111111111111111111111101111111111111000000000000000000000;
		42198: Delta = 69'sb000000000000000000000000000000000100000000000001000000000000000000000;
		32365: Delta = 69'sb111111111111111111111111111111111100000000000001000000000000000000000;
		18496: Delta = 69'sb000000000000000000000000000000000011111111111111000000000000000000000;
		8663: Delta = 69'sb111111111111111111111111111111111011111111111111000000000000000000000;
		21684: Delta = 69'sb000000000000000000000000000000001000000000000001000000000000000000000;
		2018: Delta = 69'sb111111111111111111111111111111111000000000000001000000000000000000000;
		48843: Delta = 69'sb000000000000000000000000000000000111111111111111000000000000000000000;
		29177: Delta = 69'sb111111111111111111111111111111110111111111111111000000000000000000000;
		31517: Delta = 69'sb000000000000000000000000000000010000000000000001000000000000000000000;
		43046: Delta = 69'sb111111111111111111111111111111110000000000000001000000000000000000000;
		7815: Delta = 69'sb000000000000000000000000000000001111111111111111000000000000000000000;
		19344: Delta = 69'sb111111111111111111111111111111101111111111111111000000000000000000000;
		322: Delta = 69'sb000000000000000000000000000000100000000000000001000000000000000000000;
		23380: Delta = 69'sb111111111111111111111111111111100000000000000001000000000000000000000;
		27481: Delta = 69'sb000000000000000000000000000000011111111111111111000000000000000000000;
		50539: Delta = 69'sb111111111111111111111111111111011111111111111111000000000000000000000;
		39654: Delta = 69'sb000000000000000000000000000001000000000000000001000000000000000000000;
		34909: Delta = 69'sb111111111111111111111111111111000000000000000001000000000000000000000;
		15952: Delta = 69'sb000000000000000000000000000000111111111111111111000000000000000000000;
		11207: Delta = 69'sb111111111111111111111111111110111111111111111111000000000000000000000;
		16596: Delta = 69'sb000000000000000000000000000010000000000000000001000000000000000000000;
		7106: Delta = 69'sb111111111111111111111111111110000000000000000001000000000000000000000;
		43755: Delta = 69'sb000000000000000000000000000001111111111111111111000000000000000000000;
		34265: Delta = 69'sb111111111111111111111111111101111111111111111111000000000000000000000;
		21341: Delta = 69'sb000000000000000000000000000100000000000000000001000000000000000000000;
		2361: Delta = 69'sb111111111111111111111111111100000000000000000001000000000000000000000;
		48500: Delta = 69'sb000000000000000000000000000011111111111111111111000000000000000000000;
		29520: Delta = 69'sb111111111111111111111111111011111111111111111111000000000000000000000;
		30831: Delta = 69'sb000000000000000000000000001000000000000000000001000000000000000000000;
		43732: Delta = 69'sb111111111111111111111111111000000000000000000001000000000000000000000;
		7129: Delta = 69'sb000000000000000000000000000111111111111111111111000000000000000000000;
		20030: Delta = 69'sb111111111111111111111111110111111111111111111111000000000000000000000;
		49811: Delta = 69'sb000000000000000000000000010000000000000000000001000000000000000000000;
		24752: Delta = 69'sb111111111111111111111111110000000000000000000001000000000000000000000;
		26109: Delta = 69'sb000000000000000000000000001111111111111111111111000000000000000000000;
		1050: Delta = 69'sb111111111111111111111111101111111111111111111111000000000000000000000;
		36910: Delta = 69'sb000000000000000000000000100000000000000000000001000000000000000000000;
		37653: Delta = 69'sb111111111111111111111111100000000000000000000001000000000000000000000;
		13208: Delta = 69'sb000000000000000000000000011111111111111111111111000000000000000000000;
		13951: Delta = 69'sb111111111111111111111111011111111111111111111111000000000000000000000;
		11108: Delta = 69'sb000000000000000000000001000000000000000000000001000000000000000000000;
		12594: Delta = 69'sb111111111111111111111111000000000000000000000001000000000000000000000;
		38267: Delta = 69'sb000000000000000000000000111111111111111111111111000000000000000000000;
		39753: Delta = 69'sb111111111111111111111110111111111111111111111111000000000000000000000;
		10365: Delta = 69'sb000000000000000000000010000000000000000000000001000000000000000000000;
		13337: Delta = 69'sb111111111111111111111110000000000000000000000001000000000000000000000;
		37524: Delta = 69'sb000000000000000000000001111111111111111111111111000000000000000000000;
		40496: Delta = 69'sb111111111111111111111101111111111111111111111111000000000000000000000;
		8879: Delta = 69'sb000000000000000000000100000000000000000000000001000000000000000000000;
		14823: Delta = 69'sb111111111111111111111100000000000000000000000001000000000000000000000;
		36038: Delta = 69'sb000000000000000000000011111111111111111111111111000000000000000000000;
		41982: Delta = 69'sb111111111111111111111011111111111111111111111111000000000000000000000;
		5907: Delta = 69'sb000000000000000000001000000000000000000000000001000000000000000000000;
		17795: Delta = 69'sb111111111111111111111000000000000000000000000001000000000000000000000;
		33066: Delta = 69'sb000000000000000000000111111111111111111111111111000000000000000000000;
		44954: Delta = 69'sb111111111111111111110111111111111111111111111111000000000000000000000;
		50824: Delta = 69'sb000000000000000000010000000000000000000000000001000000000000000000000;
		23739: Delta = 69'sb111111111111111111110000000000000000000000000001000000000000000000000;
		27122: Delta = 69'sb000000000000000000001111111111111111111111111111000000000000000000000;
		37: Delta = 69'sb111111111111111111101111111111111111111111111111000000000000000000000;
		38936: Delta = 69'sb000000000000000000100000000000000000000000000001000000000000000000000;
		35627: Delta = 69'sb111111111111111111100000000000000000000000000001000000000000000000000;
		15234: Delta = 69'sb000000000000000000011111111111111111111111111111000000000000000000000;
		11925: Delta = 69'sb111111111111111111011111111111111111111111111111000000000000000000000;
		15160: Delta = 69'sb000000000000000001000000000000000000000000000001000000000000000000000;
		8542: Delta = 69'sb111111111111111111000000000000000000000000000001000000000000000000000;
		42319: Delta = 69'sb000000000000000000111111111111111111111111111111000000000000000000000;
		35701: Delta = 69'sb111111111111111110111111111111111111111111111111000000000000000000000;
		18469: Delta = 69'sb000000000000000010000000000000000000000000000001000000000000000000000;
		5233: Delta = 69'sb111111111111111110000000000000000000000000000001000000000000000000000;
		45628: Delta = 69'sb000000000000000001111111111111111111111111111111000000000000000000000;
		32392: Delta = 69'sb111111111111111101111111111111111111111111111111000000000000000000000;
		25087: Delta = 69'sb000000000000000100000000000000000000000000000001000000000000000000000;
		49476: Delta = 69'sb111111111111111100000000000000000000000000000001000000000000000000000;
		1385: Delta = 69'sb000000000000000011111111111111111111111111111111000000000000000000000;
		25774: Delta = 69'sb111111111111111011111111111111111111111111111111000000000000000000000;
		38323: Delta = 69'sb000000000000001000000000000000000000000000000001000000000000000000000;
		36240: Delta = 69'sb111111111111111000000000000000000000000000000001000000000000000000000;
		14621: Delta = 69'sb000000000000000111111111111111111111111111111111000000000000000000000;
		12538: Delta = 69'sb111111111111110111111111111111111111111111111111000000000000000000000;
		13934: Delta = 69'sb000000000000010000000000000000000000000000000001000000000000000000000;
		9768: Delta = 69'sb111111111111110000000000000000000000000000000001000000000000000000000;
		41093: Delta = 69'sb000000000000001111111111111111111111111111111111000000000000000000000;
		36927: Delta = 69'sb111111111111101111111111111111111111111111111111000000000000000000000;
		16017: Delta = 69'sb000000000000100000000000000000000000000000000001000000000000000000000;
		7685: Delta = 69'sb111111111111100000000000000000000000000000000001000000000000000000000;
		43176: Delta = 69'sb000000000000011111111111111111111111111111111111000000000000000000000;
		34844: Delta = 69'sb111111111111011111111111111111111111111111111111000000000000000000000;
		20183: Delta = 69'sb000000000001000000000000000000000000000000000001000000000000000000000;
		3519: Delta = 69'sb111111111111000000000000000000000000000000000001000000000000000000000;
		47342: Delta = 69'sb000000000000111111111111111111111111111111111111000000000000000000000;
		30678: Delta = 69'sb111111111110111111111111111111111111111111111111000000000000000000000;
		28515: Delta = 69'sb000000000010000000000000000000000000000000000001000000000000000000000;
		46048: Delta = 69'sb111111111110000000000000000000000000000000000001000000000000000000000;
		4813: Delta = 69'sb000000000001111111111111111111111111111111111111000000000000000000000;
		22346: Delta = 69'sb111111111101111111111111111111111111111111111111000000000000000000000;
		45179: Delta = 69'sb000000000100000000000000000000000000000000000001000000000000000000000;
		29384: Delta = 69'sb111111111100000000000000000000000000000000000001000000000000000000000;
		21477: Delta = 69'sb000000000011111111111111111111111111111111111111000000000000000000000;
		5682: Delta = 69'sb111111111011111111111111111111111111111111111111000000000000000000000;
		27646: Delta = 69'sb000000001000000000000000000000000000000000000001000000000000000000000;
		46917: Delta = 69'sb111111111000000000000000000000000000000000000001000000000000000000000;
		3944: Delta = 69'sb000000000111111111111111111111111111111111111111000000000000000000000;
		23215: Delta = 69'sb111111110111111111111111111111111111111111111111000000000000000000000;
		43441: Delta = 69'sb000000010000000000000000000000000000000000000001000000000000000000000;
		31122: Delta = 69'sb111111110000000000000000000000000000000000000001000000000000000000000;
		19739: Delta = 69'sb000000001111111111111111111111111111111111111111000000000000000000000;
		7420: Delta = 69'sb111111101111111111111111111111111111111111111111000000000000000000000;
		24170: Delta = 69'sb000000100000000000000000000000000000000000000001000000000000000000000;
		50393: Delta = 69'sb111111100000000000000000000000000000000000000001000000000000000000000;
		468: Delta = 69'sb000000011111111111111111111111111111111111111111000000000000000000000;
		26691: Delta = 69'sb111111011111111111111111111111111111111111111111000000000000000000000;
		36489: Delta = 69'sb000001000000000000000000000000000000000000000001000000000000000000000;
		38074: Delta = 69'sb111111000000000000000000000000000000000000000001000000000000000000000;
		12787: Delta = 69'sb000000111111111111111111111111111111111111111111000000000000000000000;
		14372: Delta = 69'sb111110111111111111111111111111111111111111111111000000000000000000000;
		10266: Delta = 69'sb000010000000000000000000000000000000000000000001000000000000000000000;
		13436: Delta = 69'sb111110000000000000000000000000000000000000000001000000000000000000000;
		37425: Delta = 69'sb000001111111111111111111111111111111111111111111000000000000000000000;
		40595: Delta = 69'sb111101111111111111111111111111111111111111111111000000000000000000000;
		8681: Delta = 69'sb000100000000000000000000000000000000000000000001000000000000000000000;
		15021: Delta = 69'sb111100000000000000000000000000000000000000000001000000000000000000000;
		35840: Delta = 69'sb000011111111111111111111111111111111111111111111000000000000000000000;
		42180: Delta = 69'sb111011111111111111111111111111111111111111111111000000000000000000000;
		5511: Delta = 69'sb001000000000000000000000000000000000000000000001000000000000000000000;
		18191: Delta = 69'sb111000000000000000000000000000000000000000000001000000000000000000000;
		32670: Delta = 69'sb000111111111111111111111111111111111111111111111000000000000000000000;
		45350: Delta = 69'sb110111111111111111111111111111111111111111111111000000000000000000000;
		50032: Delta = 69'sb010000000000000000000000000000000000000000000001000000000000000000000;
		24531: Delta = 69'sb110000000000000000000000000000000000000000000001000000000000000000000;
		26330: Delta = 69'sb001111111111111111111111111111111111111111111111000000000000000000000;
		829: Delta = 69'sb101111111111111111111111111111111111111111111111000000000000000000000;
		20245: Delta = 69'sb000000000000000000000000000000000000000000000110000000000000000000000;
		30616: Delta = 69'sb111111111111111111111111111111111111111111111010000000000000000000000;
		16788: Delta = 69'sb000000000000000000000000000000000000000000001010000000000000000000000;
		34073: Delta = 69'sb111111111111111111111111111111111111111111110110000000000000000000000;
		9874: Delta = 69'sb000000000000000000000000000000000000000000010010000000000000000000000;
		37530: Delta = 69'sb111111111111111111111111111111111111111111110010000000000000000000000;
		13331: Delta = 69'sb000000000000000000000000000000000000000000001110000000000000000000000;
		40987: Delta = 69'sb111111111111111111111111111111111111111111101110000000000000000000000;
		46907: Delta = 69'sb000000000000000000000000000000000000000000100010000000000000000000000;
		497: Delta = 69'sb111111111111111111111111111111111111111111100010000000000000000000000;
		50364: Delta = 69'sb000000000000000000000000000000000000000000011110000000000000000000000;
		3954: Delta = 69'sb111111111111111111111111111111111111111111011110000000000000000000000;
		19251: Delta = 69'sb000000000000000000000000000000000000000001000010000000000000000000000;
		28153: Delta = 69'sb111111111111111111111111111111111111111111000010000000000000000000000;
		22708: Delta = 69'sb000000000000000000000000000000000000000000111110000000000000000000000;
		31610: Delta = 69'sb111111111111111111111111111111111111111110111110000000000000000000000;
		14800: Delta = 69'sb000000000000000000000000000000000000000010000010000000000000000000000;
		32604: Delta = 69'sb111111111111111111111111111111111111111110000010000000000000000000000;
		18257: Delta = 69'sb000000000000000000000000000000000000000001111110000000000000000000000;
		36061: Delta = 69'sb111111111111111111111111111111111111111101111110000000000000000000000;
		5898: Delta = 69'sb000000000000000000000000000000000000000100000010000000000000000000000;
		41506: Delta = 69'sb111111111111111111111111111111111111111100000010000000000000000000000;
		9355: Delta = 69'sb000000000000000000000000000000000000000011111110000000000000000000000;
		44963: Delta = 69'sb111111111111111111111111111111111111111011111110000000000000000000000;
		38955: Delta = 69'sb000000000000000000000000000000000000001000000010000000000000000000000;
		8449: Delta = 69'sb111111111111111111111111111111111111111000000010000000000000000000000;
		42412: Delta = 69'sb000000000000000000000000000000000000000111111110000000000000000000000;
		11906: Delta = 69'sb111111111111111111111111111111111111110111111110000000000000000000000;
		3347: Delta = 69'sb000000000000000000000000000000000000010000000010000000000000000000000;
		44057: Delta = 69'sb111111111111111111111111111111111111110000000010000000000000000000000;
		6804: Delta = 69'sb000000000000000000000000000000000000001111111110000000000000000000000;
		47514: Delta = 69'sb111111111111111111111111111111111111101111111110000000000000000000000;
		33853: Delta = 69'sb000000000000000000000000000000000000100000000010000000000000000000000;
		13551: Delta = 69'sb111111111111111111111111111111111111100000000010000000000000000000000;
		37310: Delta = 69'sb000000000000000000000000000000000000011111111110000000000000000000000;
		17008: Delta = 69'sb111111111111111111111111111111111111011111111110000000000000000000000;
		44004: Delta = 69'sb000000000000000000000000000000000001000000000010000000000000000000000;
		3400: Delta = 69'sb111111111111111111111111111111111111000000000010000000000000000000000;
		47461: Delta = 69'sb000000000000000000000000000000000000111111111110000000000000000000000;
		6857: Delta = 69'sb111111111111111111111111111111111110111111111110000000000000000000000;
		13445: Delta = 69'sb000000000000000000000000000000000010000000000010000000000000000000000;
		33959: Delta = 69'sb111111111111111111111111111111111110000000000010000000000000000000000;
		16902: Delta = 69'sb000000000000000000000000000000000001111111111110000000000000000000000;
		37416: Delta = 69'sb111111111111111111111111111111111101111111111110000000000000000000000;
		3188: Delta = 69'sb000000000000000000000000000000000100000000000010000000000000000000000;
		44216: Delta = 69'sb111111111111111111111111111111111100000000000010000000000000000000000;
		6645: Delta = 69'sb000000000000000000000000000000000011111111111110000000000000000000000;
		47673: Delta = 69'sb111111111111111111111111111111111011111111111110000000000000000000000;
		33535: Delta = 69'sb000000000000000000000000000000001000000000000010000000000000000000000;
		13869: Delta = 69'sb111111111111111111111111111111111000000000000010000000000000000000000;
		36992: Delta = 69'sb000000000000000000000000000000000111111111111110000000000000000000000;
		17326: Delta = 69'sb111111111111111111111111111111110111111111111110000000000000000000000;
		43368: Delta = 69'sb000000000000000000000000000000010000000000000010000000000000000000000;
		4036: Delta = 69'sb111111111111111111111111111111110000000000000010000000000000000000000;
		46825: Delta = 69'sb000000000000000000000000000000001111111111111110000000000000000000000;
		7493: Delta = 69'sb111111111111111111111111111111101111111111111110000000000000000000000;
		12173: Delta = 69'sb000000000000000000000000000000100000000000000010000000000000000000000;
		35231: Delta = 69'sb111111111111111111111111111111100000000000000010000000000000000000000;
		15630: Delta = 69'sb000000000000000000000000000000011111111111111110000000000000000000000;
		38688: Delta = 69'sb111111111111111111111111111111011111111111111110000000000000000000000;
		644: Delta = 69'sb000000000000000000000000000001000000000000000010000000000000000000000;
		46760: Delta = 69'sb111111111111111111111111111111000000000000000010000000000000000000000;
		4101: Delta = 69'sb000000000000000000000000000000111111111111111110000000000000000000000;
		50217: Delta = 69'sb111111111111111111111111111110111111111111111110000000000000000000000;
		28447: Delta = 69'sb000000000000000000000000000010000000000000000010000000000000000000000;
		18957: Delta = 69'sb111111111111111111111111111110000000000000000010000000000000000000000;
		31904: Delta = 69'sb000000000000000000000000000001111111111111111110000000000000000000000;
		22414: Delta = 69'sb111111111111111111111111111101111111111111111110000000000000000000000;
		33192: Delta = 69'sb000000000000000000000000000100000000000000000010000000000000000000000;
		14212: Delta = 69'sb111111111111111111111111111100000000000000000010000000000000000000000;
		36649: Delta = 69'sb000000000000000000000000000011111111111111111110000000000000000000000;
		17669: Delta = 69'sb111111111111111111111111111011111111111111111110000000000000000000000;
		42682: Delta = 69'sb000000000000000000000000001000000000000000000010000000000000000000000;
		4722: Delta = 69'sb111111111111111111111111111000000000000000000010000000000000000000000;
		46139: Delta = 69'sb000000000000000000000000000111111111111111111110000000000000000000000;
		8179: Delta = 69'sb111111111111111111111111110111111111111111111110000000000000000000000;
		10801: Delta = 69'sb000000000000000000000000010000000000000000000010000000000000000000000;
		36603: Delta = 69'sb111111111111111111111111110000000000000000000010000000000000000000000;
		14258: Delta = 69'sb000000000000000000000000001111111111111111111110000000000000000000000;
		40060: Delta = 69'sb111111111111111111111111101111111111111111111110000000000000000000000;
		48761: Delta = 69'sb000000000000000000000000100000000000000000000010000000000000000000000;
		49504: Delta = 69'sb111111111111111111111111100000000000000000000010000000000000000000000;
		1357: Delta = 69'sb000000000000000000000000011111111111111111111110000000000000000000000;
		2100: Delta = 69'sb111111111111111111111111011111111111111111111110000000000000000000000;
		22959: Delta = 69'sb000000000000000000000001000000000000000000000010000000000000000000000;
		24445: Delta = 69'sb111111111111111111111111000000000000000000000010000000000000000000000;
		26416: Delta = 69'sb000000000000000000000000111111111111111111111110000000000000000000000;
		27902: Delta = 69'sb111111111111111111111110111111111111111111111110000000000000000000000;
		22216: Delta = 69'sb000000000000000000000010000000000000000000000010000000000000000000000;
		25188: Delta = 69'sb111111111111111111111110000000000000000000000010000000000000000000000;
		25673: Delta = 69'sb000000000000000000000001111111111111111111111110000000000000000000000;
		28645: Delta = 69'sb111111111111111111111101111111111111111111111110000000000000000000000;
		20730: Delta = 69'sb000000000000000000000100000000000000000000000010000000000000000000000;
		26674: Delta = 69'sb111111111111111111111100000000000000000000000010000000000000000000000;
		24187: Delta = 69'sb000000000000000000000011111111111111111111111110000000000000000000000;
		30131: Delta = 69'sb111111111111111111111011111111111111111111111110000000000000000000000;
		17758: Delta = 69'sb000000000000000000001000000000000000000000000010000000000000000000000;
		29646: Delta = 69'sb111111111111111111111000000000000000000000000010000000000000000000000;
		21215: Delta = 69'sb000000000000000000000111111111111111111111111110000000000000000000000;
		33103: Delta = 69'sb111111111111111111110111111111111111111111111110000000000000000000000;
		11814: Delta = 69'sb000000000000000000010000000000000000000000000010000000000000000000000;
		35590: Delta = 69'sb111111111111111111110000000000000000000000000010000000000000000000000;
		15271: Delta = 69'sb000000000000000000001111111111111111111111111110000000000000000000000;
		39047: Delta = 69'sb111111111111111111101111111111111111111111111110000000000000000000000;
		50787: Delta = 69'sb000000000000000000100000000000000000000000000010000000000000000000000;
		47478: Delta = 69'sb111111111111111111100000000000000000000000000010000000000000000000000;
		3383: Delta = 69'sb000000000000000000011111111111111111111111111110000000000000000000000;
		74: Delta = 69'sb111111111111111111011111111111111111111111111110000000000000000000000;
		27011: Delta = 69'sb000000000000000001000000000000000000000000000010000000000000000000000;
		20393: Delta = 69'sb111111111111111111000000000000000000000000000010000000000000000000000;
		30468: Delta = 69'sb000000000000000000111111111111111111111111111110000000000000000000000;
		23850: Delta = 69'sb111111111111111110111111111111111111111111111110000000000000000000000;
		30320: Delta = 69'sb000000000000000010000000000000000000000000000010000000000000000000000;
		17084: Delta = 69'sb111111111111111110000000000000000000000000000010000000000000000000000;
		33777: Delta = 69'sb000000000000000001111111111111111111111111111110000000000000000000000;
		20541: Delta = 69'sb111111111111111101111111111111111111111111111110000000000000000000000;
		36938: Delta = 69'sb000000000000000100000000000000000000000000000010000000000000000000000;
		10466: Delta = 69'sb111111111111111100000000000000000000000000000010000000000000000000000;
		40395: Delta = 69'sb000000000000000011111111111111111111111111111110000000000000000000000;
		13923: Delta = 69'sb111111111111111011111111111111111111111111111110000000000000000000000;
		50174: Delta = 69'sb000000000000001000000000000000000000000000000010000000000000000000000;
		48091: Delta = 69'sb111111111111111000000000000000000000000000000010000000000000000000000;
		2770: Delta = 69'sb000000000000000111111111111111111111111111111110000000000000000000000;
		687: Delta = 69'sb111111111111110111111111111111111111111111111110000000000000000000000;
		25785: Delta = 69'sb000000000000010000000000000000000000000000000010000000000000000000000;
		21619: Delta = 69'sb111111111111110000000000000000000000000000000010000000000000000000000;
		29242: Delta = 69'sb000000000000001111111111111111111111111111111110000000000000000000000;
		25076: Delta = 69'sb111111111111101111111111111111111111111111111110000000000000000000000;
		27868: Delta = 69'sb000000000000100000000000000000000000000000000010000000000000000000000;
		19536: Delta = 69'sb111111111111100000000000000000000000000000000010000000000000000000000;
		31325: Delta = 69'sb000000000000011111111111111111111111111111111110000000000000000000000;
		22993: Delta = 69'sb111111111111011111111111111111111111111111111110000000000000000000000;
		32034: Delta = 69'sb000000000001000000000000000000000000000000000010000000000000000000000;
		15370: Delta = 69'sb111111111111000000000000000000000000000000000010000000000000000000000;
		35491: Delta = 69'sb000000000000111111111111111111111111111111111110000000000000000000000;
		18827: Delta = 69'sb111111111110111111111111111111111111111111111110000000000000000000000;
		40366: Delta = 69'sb000000000010000000000000000000000000000000000010000000000000000000000;
		7038: Delta = 69'sb111111111110000000000000000000000000000000000010000000000000000000000;
		43823: Delta = 69'sb000000000001111111111111111111111111111111111110000000000000000000000;
		10495: Delta = 69'sb111111111101111111111111111111111111111111111110000000000000000000000;
		6169: Delta = 69'sb000000000100000000000000000000000000000000000010000000000000000000000;
		41235: Delta = 69'sb111111111100000000000000000000000000000000000010000000000000000000000;
		9626: Delta = 69'sb000000000011111111111111111111111111111111111110000000000000000000000;
		44692: Delta = 69'sb111111111011111111111111111111111111111111111110000000000000000000000;
		39497: Delta = 69'sb000000001000000000000000000000000000000000000010000000000000000000000;
		7907: Delta = 69'sb111111111000000000000000000000000000000000000010000000000000000000000;
		42954: Delta = 69'sb000000000111111111111111111111111111111111111110000000000000000000000;
		11364: Delta = 69'sb111111110111111111111111111111111111111111111110000000000000000000000;
		4431: Delta = 69'sb000000010000000000000000000000000000000000000010000000000000000000000;
		42973: Delta = 69'sb111111110000000000000000000000000000000000000010000000000000000000000;
		7888: Delta = 69'sb000000001111111111111111111111111111111111111110000000000000000000000;
		46430: Delta = 69'sb111111101111111111111111111111111111111111111110000000000000000000000;
		36021: Delta = 69'sb000000100000000000000000000000000000000000000010000000000000000000000;
		11383: Delta = 69'sb111111100000000000000000000000000000000000000010000000000000000000000;
		39478: Delta = 69'sb000000011111111111111111111111111111111111111110000000000000000000000;
		14840: Delta = 69'sb111111011111111111111111111111111111111111111110000000000000000000000;
		48340: Delta = 69'sb000001000000000000000000000000000000000000000010000000000000000000000;
		49925: Delta = 69'sb111111000000000000000000000000000000000000000010000000000000000000000;
		936: Delta = 69'sb000000111111111111111111111111111111111111111110000000000000000000000;
		2521: Delta = 69'sb111110111111111111111111111111111111111111111110000000000000000000000;
		22117: Delta = 69'sb000010000000000000000000000000000000000000000010000000000000000000000;
		25287: Delta = 69'sb111110000000000000000000000000000000000000000010000000000000000000000;
		25574: Delta = 69'sb000001111111111111111111111111111111111111111110000000000000000000000;
		28744: Delta = 69'sb111101111111111111111111111111111111111111111110000000000000000000000;
		20532: Delta = 69'sb000100000000000000000000000000000000000000000010000000000000000000000;
		26872: Delta = 69'sb111100000000000000000000000000000000000000000010000000000000000000000;
		23989: Delta = 69'sb000011111111111111111111111111111111111111111110000000000000000000000;
		30329: Delta = 69'sb111011111111111111111111111111111111111111111110000000000000000000000;
		17362: Delta = 69'sb001000000000000000000000000000000000000000000010000000000000000000000;
		30042: Delta = 69'sb111000000000000000000000000000000000000000000010000000000000000000000;
		20819: Delta = 69'sb000111111111111111111111111111111111111111111110000000000000000000000;
		33499: Delta = 69'sb110111111111111111111111111111111111111111111110000000000000000000000;
		11022: Delta = 69'sb010000000000000000000000000000000000000000000010000000000000000000000;
		36382: Delta = 69'sb110000000000000000000000000000000000000000000010000000000000000000000;
		14479: Delta = 69'sb001111111111111111111111111111111111111111111110000000000000000000000;
		39839: Delta = 69'sb101111111111111111111111111111111111111111111110000000000000000000000;
		40490: Delta = 69'sb000000000000000000000000000000000000000000001100000000000000000000000;
		10371: Delta = 69'sb111111111111111111111111111111111111111111110100000000000000000000000;
		33576: Delta = 69'sb000000000000000000000000000000000000000000010100000000000000000000000;
		17285: Delta = 69'sb111111111111111111111111111111111111111111101100000000000000000000000;
		19748: Delta = 69'sb000000000000000000000000000000000000000000100100000000000000000000000;
		24199: Delta = 69'sb111111111111111111111111111111111111111111100100000000000000000000000;
		26662: Delta = 69'sb000000000000000000000000000000000000000000011100000000000000000000000;
		31113: Delta = 69'sb111111111111111111111111111111111111111111011100000000000000000000000;
		42953: Delta = 69'sb000000000000000000000000000000000000000001000100000000000000000000000;
		994: Delta = 69'sb111111111111111111111111111111111111111111000100000000000000000000000;
		49867: Delta = 69'sb000000000000000000000000000000000000000000111100000000000000000000000;
		7908: Delta = 69'sb111111111111111111111111111111111111111110111100000000000000000000000;
		38502: Delta = 69'sb000000000000000000000000000000000000000010000100000000000000000000000;
		5445: Delta = 69'sb111111111111111111111111111111111111111110000100000000000000000000000;
		45416: Delta = 69'sb000000000000000000000000000000000000000001111100000000000000000000000;
		12359: Delta = 69'sb111111111111111111111111111111111111111101111100000000000000000000000;
		29600: Delta = 69'sb000000000000000000000000000000000000000100000100000000000000000000000;
		14347: Delta = 69'sb111111111111111111111111111111111111111100000100000000000000000000000;
		36514: Delta = 69'sb000000000000000000000000000000000000000011111100000000000000000000000;
		21261: Delta = 69'sb111111111111111111111111111111111111111011111100000000000000000000000;
		11796: Delta = 69'sb000000000000000000000000000000000000001000000100000000000000000000000;
		32151: Delta = 69'sb111111111111111111111111111111111111111000000100000000000000000000000;
		18710: Delta = 69'sb000000000000000000000000000000000000000111111100000000000000000000000;
		39065: Delta = 69'sb111111111111111111111111111111111111110111111100000000000000000000000;
		27049: Delta = 69'sb000000000000000000000000000000000000010000000100000000000000000000000;
		16898: Delta = 69'sb111111111111111111111111111111111111110000000100000000000000000000000;
		33963: Delta = 69'sb000000000000000000000000000000000000001111111100000000000000000000000;
		23812: Delta = 69'sb111111111111111111111111111111111111101111111100000000000000000000000;
		6694: Delta = 69'sb000000000000000000000000000000000000100000000100000000000000000000000;
		37253: Delta = 69'sb111111111111111111111111111111111111100000000100000000000000000000000;
		13608: Delta = 69'sb000000000000000000000000000000000000011111111100000000000000000000000;
		44167: Delta = 69'sb111111111111111111111111111111111111011111111100000000000000000000000;
		16845: Delta = 69'sb000000000000000000000000000000000001000000000100000000000000000000000;
		27102: Delta = 69'sb111111111111111111111111111111111111000000000100000000000000000000000;
		23759: Delta = 69'sb000000000000000000000000000000000000111111111100000000000000000000000;
		34016: Delta = 69'sb111111111111111111111111111111111110111111111100000000000000000000000;
		37147: Delta = 69'sb000000000000000000000000000000000010000000000100000000000000000000000;
		6800: Delta = 69'sb111111111111111111111111111111111110000000000100000000000000000000000;
		44061: Delta = 69'sb000000000000000000000000000000000001111111111100000000000000000000000;
		13714: Delta = 69'sb111111111111111111111111111111111101111111111100000000000000000000000;
		26890: Delta = 69'sb000000000000000000000000000000000100000000000100000000000000000000000;
		17057: Delta = 69'sb111111111111111111111111111111111100000000000100000000000000000000000;
		33804: Delta = 69'sb000000000000000000000000000000000011111111111100000000000000000000000;
		23971: Delta = 69'sb111111111111111111111111111111111011111111111100000000000000000000000;
		6376: Delta = 69'sb000000000000000000000000000000001000000000000100000000000000000000000;
		37571: Delta = 69'sb111111111111111111111111111111111000000000000100000000000000000000000;
		13290: Delta = 69'sb000000000000000000000000000000000111111111111100000000000000000000000;
		44485: Delta = 69'sb111111111111111111111111111111110111111111111100000000000000000000000;
		16209: Delta = 69'sb000000000000000000000000000000010000000000000100000000000000000000000;
		27738: Delta = 69'sb111111111111111111111111111111110000000000000100000000000000000000000;
		23123: Delta = 69'sb000000000000000000000000000000001111111111111100000000000000000000000;
		34652: Delta = 69'sb111111111111111111111111111111101111111111111100000000000000000000000;
		35875: Delta = 69'sb000000000000000000000000000000100000000000000100000000000000000000000;
		8072: Delta = 69'sb111111111111111111111111111111100000000000000100000000000000000000000;
		42789: Delta = 69'sb000000000000000000000000000000011111111111111100000000000000000000000;
		14986: Delta = 69'sb111111111111111111111111111111011111111111111100000000000000000000000;
		24346: Delta = 69'sb000000000000000000000000000001000000000000000100000000000000000000000;
		19601: Delta = 69'sb111111111111111111111111111111000000000000000100000000000000000000000;
		31260: Delta = 69'sb000000000000000000000000000000111111111111111100000000000000000000000;
		26515: Delta = 69'sb111111111111111111111111111110111111111111111100000000000000000000000;
		1288: Delta = 69'sb000000000000000000000000000010000000000000000100000000000000000000000;
		42659: Delta = 69'sb111111111111111111111111111110000000000000000100000000000000000000000;
		8202: Delta = 69'sb000000000000000000000000000001111111111111111100000000000000000000000;
		49573: Delta = 69'sb111111111111111111111111111101111111111111111100000000000000000000000;
		6033: Delta = 69'sb000000000000000000000000000100000000000000000100000000000000000000000;
		37914: Delta = 69'sb111111111111111111111111111100000000000000000100000000000000000000000;
		12947: Delta = 69'sb000000000000000000000000000011111111111111111100000000000000000000000;
		44828: Delta = 69'sb111111111111111111111111111011111111111111111100000000000000000000000;
		15523: Delta = 69'sb000000000000000000000000001000000000000000000100000000000000000000000;
		28424: Delta = 69'sb111111111111111111111111111000000000000000000100000000000000000000000;
		22437: Delta = 69'sb000000000000000000000000000111111111111111111100000000000000000000000;
		35338: Delta = 69'sb111111111111111111111111110111111111111111111100000000000000000000000;
		34503: Delta = 69'sb000000000000000000000000010000000000000000000100000000000000000000000;
		9444: Delta = 69'sb111111111111111111111111110000000000000000000100000000000000000000000;
		41417: Delta = 69'sb000000000000000000000000001111111111111111111100000000000000000000000;
		16358: Delta = 69'sb111111111111111111111111101111111111111111111100000000000000000000000;
		21602: Delta = 69'sb000000000000000000000000100000000000000000000100000000000000000000000;
		22345: Delta = 69'sb111111111111111111111111100000000000000000000100000000000000000000000;
		28516: Delta = 69'sb000000000000000000000000011111111111111111111100000000000000000000000;
		29259: Delta = 69'sb111111111111111111111111011111111111111111111100000000000000000000000;
		46661: Delta = 69'sb000000000000000000000001000000000000000000000100000000000000000000000;
		48147: Delta = 69'sb111111111111111111111111000000000000000000000100000000000000000000000;
		2714: Delta = 69'sb000000000000000000000000111111111111111111111100000000000000000000000;
		4200: Delta = 69'sb111111111111111111111110111111111111111111111100000000000000000000000;
		45918: Delta = 69'sb000000000000000000000010000000000000000000000100000000000000000000000;
		48890: Delta = 69'sb111111111111111111111110000000000000000000000100000000000000000000000;
		1971: Delta = 69'sb000000000000000000000001111111111111111111111100000000000000000000000;
		4943: Delta = 69'sb111111111111111111111101111111111111111111111100000000000000000000000;
		44432: Delta = 69'sb000000000000000000000100000000000000000000000100000000000000000000000;
		50376: Delta = 69'sb111111111111111111111100000000000000000000000100000000000000000000000;
		485: Delta = 69'sb000000000000000000000011111111111111111111111100000000000000000000000;
		6429: Delta = 69'sb111111111111111111111011111111111111111111111100000000000000000000000;
		41460: Delta = 69'sb000000000000000000001000000000000000000000000100000000000000000000000;
		2487: Delta = 69'sb111111111111111111111000000000000000000000000100000000000000000000000;
		48374: Delta = 69'sb000000000000000000000111111111111111111111111100000000000000000000000;
		9401: Delta = 69'sb111111111111111111110111111111111111111111111100000000000000000000000;
		35516: Delta = 69'sb000000000000000000010000000000000000000000000100000000000000000000000;
		8431: Delta = 69'sb111111111111111111110000000000000000000000000100000000000000000000000;
		42430: Delta = 69'sb000000000000000000001111111111111111111111111100000000000000000000000;
		15345: Delta = 69'sb111111111111111111101111111111111111111111111100000000000000000000000;
		23628: Delta = 69'sb000000000000000000100000000000000000000000000100000000000000000000000;
		20319: Delta = 69'sb111111111111111111100000000000000000000000000100000000000000000000000;
		30542: Delta = 69'sb000000000000000000011111111111111111111111111100000000000000000000000;
		27233: Delta = 69'sb111111111111111111011111111111111111111111111100000000000000000000000;
		50713: Delta = 69'sb000000000000000001000000000000000000000000000100000000000000000000000;
		44095: Delta = 69'sb111111111111111111000000000000000000000000000100000000000000000000000;
		6766: Delta = 69'sb000000000000000000111111111111111111111111111100000000000000000000000;
		148: Delta = 69'sb111111111111111110111111111111111111111111111100000000000000000000000;
		3161: Delta = 69'sb000000000000000010000000000000000000000000000100000000000000000000000;
		40786: Delta = 69'sb111111111111111110000000000000000000000000000100000000000000000000000;
		10075: Delta = 69'sb000000000000000001111111111111111111111111111100000000000000000000000;
		47700: Delta = 69'sb111111111111111101111111111111111111111111111100000000000000000000000;
		9779: Delta = 69'sb000000000000000100000000000000000000000000000100000000000000000000000;
		34168: Delta = 69'sb111111111111111100000000000000000000000000000100000000000000000000000;
		16693: Delta = 69'sb000000000000000011111111111111111111111111111100000000000000000000000;
		41082: Delta = 69'sb111111111111111011111111111111111111111111111100000000000000000000000;
		23015: Delta = 69'sb000000000000001000000000000000000000000000000100000000000000000000000;
		20932: Delta = 69'sb111111111111111000000000000000000000000000000100000000000000000000000;
		29929: Delta = 69'sb000000000000000111111111111111111111111111111100000000000000000000000;
		27846: Delta = 69'sb111111111111110111111111111111111111111111111100000000000000000000000;
		49487: Delta = 69'sb000000000000010000000000000000000000000000000100000000000000000000000;
		45321: Delta = 69'sb111111111111110000000000000000000000000000000100000000000000000000000;
		5540: Delta = 69'sb000000000000001111111111111111111111111111111100000000000000000000000;
		1374: Delta = 69'sb111111111111101111111111111111111111111111111100000000000000000000000;
		709: Delta = 69'sb000000000000100000000000000000000000000000000100000000000000000000000;
		43238: Delta = 69'sb111111111111100000000000000000000000000000000100000000000000000000000;
		7623: Delta = 69'sb000000000000011111111111111111111111111111111100000000000000000000000;
		50152: Delta = 69'sb111111111111011111111111111111111111111111111100000000000000000000000;
		4875: Delta = 69'sb000000000001000000000000000000000000000000000100000000000000000000000;
		39072: Delta = 69'sb111111111111000000000000000000000000000000000100000000000000000000000;
		11789: Delta = 69'sb000000000000111111111111111111111111111111111100000000000000000000000;
		45986: Delta = 69'sb111111111110111111111111111111111111111111111100000000000000000000000;
		13207: Delta = 69'sb000000000010000000000000000000000000000000000100000000000000000000000;
		30740: Delta = 69'sb111111111110000000000000000000000000000000000100000000000000000000000;
		20121: Delta = 69'sb000000000001111111111111111111111111111111111100000000000000000000000;
		37654: Delta = 69'sb111111111101111111111111111111111111111111111100000000000000000000000;
		29871: Delta = 69'sb000000000100000000000000000000000000000000000100000000000000000000000;
		14076: Delta = 69'sb111111111100000000000000000000000000000000000100000000000000000000000;
		36785: Delta = 69'sb000000000011111111111111111111111111111111111100000000000000000000000;
		20990: Delta = 69'sb111111111011111111111111111111111111111111111100000000000000000000000;
		12338: Delta = 69'sb000000001000000000000000000000000000000000000100000000000000000000000;
		31609: Delta = 69'sb111111111000000000000000000000000000000000000100000000000000000000000;
		19252: Delta = 69'sb000000000111111111111111111111111111111111111100000000000000000000000;
		38523: Delta = 69'sb111111110111111111111111111111111111111111111100000000000000000000000;
		28133: Delta = 69'sb000000010000000000000000000000000000000000000100000000000000000000000;
		15814: Delta = 69'sb111111110000000000000000000000000000000000000100000000000000000000000;
		35047: Delta = 69'sb000000001111111111111111111111111111111111111100000000000000000000000;
		22728: Delta = 69'sb111111101111111111111111111111111111111111111100000000000000000000000;
		8862: Delta = 69'sb000000100000000000000000000000000000000000000100000000000000000000000;
		35085: Delta = 69'sb111111100000000000000000000000000000000000000100000000000000000000000;
		15776: Delta = 69'sb000000011111111111111111111111111111111111111100000000000000000000000;
		41999: Delta = 69'sb111111011111111111111111111111111111111111111100000000000000000000000;
		21181: Delta = 69'sb000001000000000000000000000000000000000000000100000000000000000000000;
		22766: Delta = 69'sb111111000000000000000000000000000000000000000100000000000000000000000;
		28095: Delta = 69'sb000000111111111111111111111111111111111111111100000000000000000000000;
		29680: Delta = 69'sb111110111111111111111111111111111111111111111100000000000000000000000;
		45819: Delta = 69'sb000010000000000000000000000000000000000000000100000000000000000000000;
		48989: Delta = 69'sb111110000000000000000000000000000000000000000100000000000000000000000;
		1872: Delta = 69'sb000001111111111111111111111111111111111111111100000000000000000000000;
		5042: Delta = 69'sb111101111111111111111111111111111111111111111100000000000000000000000;
		44234: Delta = 69'sb000100000000000000000000000000000000000000000100000000000000000000000;
		50574: Delta = 69'sb111100000000000000000000000000000000000000000100000000000000000000000;
		287: Delta = 69'sb000011111111111111111111111111111111111111111100000000000000000000000;
		6627: Delta = 69'sb111011111111111111111111111111111111111111111100000000000000000000000;
		41064: Delta = 69'sb001000000000000000000000000000000000000000000100000000000000000000000;
		2883: Delta = 69'sb111000000000000000000000000000000000000000000100000000000000000000000;
		47978: Delta = 69'sb000111111111111111111111111111111111111111111100000000000000000000000;
		9797: Delta = 69'sb110111111111111111111111111111111111111111111100000000000000000000000;
		34724: Delta = 69'sb010000000000000000000000000000000000000000000100000000000000000000000;
		9223: Delta = 69'sb110000000000000000000000000000000000000000000100000000000000000000000;
		41638: Delta = 69'sb001111111111111111111111111111111111111111111100000000000000000000000;
		16137: Delta = 69'sb101111111111111111111111111111111111111111111100000000000000000000000;
		30119: Delta = 69'sb000000000000000000000000000000000000000000011000000000000000000000000;
		20742: Delta = 69'sb111111111111111111111111111111111111111111101000000000000000000000000;
		16291: Delta = 69'sb000000000000000000000000000000000000000000101000000000000000000000000;
		34570: Delta = 69'sb111111111111111111111111111111111111111111011000000000000000000000000;
		39496: Delta = 69'sb000000000000000000000000000000000000000001001000000000000000000000000;
		48398: Delta = 69'sb111111111111111111111111111111111111111111001000000000000000000000000;
		2463: Delta = 69'sb000000000000000000000000000000000000000000111000000000000000000000000;
		11365: Delta = 69'sb111111111111111111111111111111111111111110111000000000000000000000000;
		35045: Delta = 69'sb000000000000000000000000000000000000000010001000000000000000000000000;
		1988: Delta = 69'sb111111111111111111111111111111111111111110001000000000000000000000000;
		48873: Delta = 69'sb000000000000000000000000000000000000000001111000000000000000000000000;
		15816: Delta = 69'sb111111111111111111111111111111111111111101111000000000000000000000000;
		26143: Delta = 69'sb000000000000000000000000000000000000000100001000000000000000000000000;
		10890: Delta = 69'sb111111111111111111111111111111111111111100001000000000000000000000000;
		39971: Delta = 69'sb000000000000000000000000000000000000000011111000000000000000000000000;
		24718: Delta = 69'sb111111111111111111111111111111111111111011111000000000000000000000000;
		8339: Delta = 69'sb000000000000000000000000000000000000001000001000000000000000000000000;
		28694: Delta = 69'sb111111111111111111111111111111111111111000001000000000000000000000000;
		22167: Delta = 69'sb000000000000000000000000000000000000000111111000000000000000000000000;
		42522: Delta = 69'sb111111111111111111111111111111111111110111111000000000000000000000000;
		23592: Delta = 69'sb000000000000000000000000000000000000010000001000000000000000000000000;
		13441: Delta = 69'sb111111111111111111111111111111111111110000001000000000000000000000000;
		37420: Delta = 69'sb000000000000000000000000000000000000001111111000000000000000000000000;
		27269: Delta = 69'sb111111111111111111111111111111111111101111111000000000000000000000000;
		3237: Delta = 69'sb000000000000000000000000000000000000100000001000000000000000000000000;
		33796: Delta = 69'sb111111111111111111111111111111111111100000001000000000000000000000000;
		17065: Delta = 69'sb000000000000000000000000000000000000011111111000000000000000000000000;
		47624: Delta = 69'sb111111111111111111111111111111111111011111111000000000000000000000000;
		13388: Delta = 69'sb000000000000000000000000000000000001000000001000000000000000000000000;
		23645: Delta = 69'sb111111111111111111111111111111111111000000001000000000000000000000000;
		27216: Delta = 69'sb000000000000000000000000000000000000111111111000000000000000000000000;
		37473: Delta = 69'sb111111111111111111111111111111111110111111111000000000000000000000000;
		33690: Delta = 69'sb000000000000000000000000000000000010000000001000000000000000000000000;
		3343: Delta = 69'sb111111111111111111111111111111111110000000001000000000000000000000000;
		47518: Delta = 69'sb000000000000000000000000000000000001111111111000000000000000000000000;
		17171: Delta = 69'sb111111111111111111111111111111111101111111111000000000000000000000000;
		23433: Delta = 69'sb000000000000000000000000000000000100000000001000000000000000000000000;
		13600: Delta = 69'sb111111111111111111111111111111111100000000001000000000000000000000000;
		37261: Delta = 69'sb000000000000000000000000000000000011111111111000000000000000000000000;
		27428: Delta = 69'sb111111111111111111111111111111111011111111111000000000000000000000000;
		2919: Delta = 69'sb000000000000000000000000000000001000000000001000000000000000000000000;
		34114: Delta = 69'sb111111111111111111111111111111111000000000001000000000000000000000000;
		16747: Delta = 69'sb000000000000000000000000000000000111111111111000000000000000000000000;
		47942: Delta = 69'sb111111111111111111111111111111110111111111111000000000000000000000000;
		12752: Delta = 69'sb000000000000000000000000000000010000000000001000000000000000000000000;
		24281: Delta = 69'sb111111111111111111111111111111110000000000001000000000000000000000000;
		26580: Delta = 69'sb000000000000000000000000000000001111111111111000000000000000000000000;
		38109: Delta = 69'sb111111111111111111111111111111101111111111111000000000000000000000000;
		32418: Delta = 69'sb000000000000000000000000000000100000000000001000000000000000000000000;
		4615: Delta = 69'sb111111111111111111111111111111100000000000001000000000000000000000000;
		46246: Delta = 69'sb000000000000000000000000000000011111111111111000000000000000000000000;
		18443: Delta = 69'sb111111111111111111111111111111011111111111111000000000000000000000000;
		20889: Delta = 69'sb000000000000000000000000000001000000000000001000000000000000000000000;
		16144: Delta = 69'sb111111111111111111111111111111000000000000001000000000000000000000000;
		34717: Delta = 69'sb000000000000000000000000000000111111111111111000000000000000000000000;
		29972: Delta = 69'sb111111111111111111111111111110111111111111111000000000000000000000000;
		48692: Delta = 69'sb000000000000000000000000000010000000000000001000000000000000000000000;
		39202: Delta = 69'sb111111111111111111111111111110000000000000001000000000000000000000000;
		11659: Delta = 69'sb000000000000000000000000000001111111111111111000000000000000000000000;
		2169: Delta = 69'sb111111111111111111111111111101111111111111111000000000000000000000000;
		2576: Delta = 69'sb000000000000000000000000000100000000000000001000000000000000000000000;
		34457: Delta = 69'sb111111111111111111111111111100000000000000001000000000000000000000000;
		16404: Delta = 69'sb000000000000000000000000000011111111111111111000000000000000000000000;
		48285: Delta = 69'sb111111111111111111111111111011111111111111111000000000000000000000000;
		12066: Delta = 69'sb000000000000000000000000001000000000000000001000000000000000000000000;
		24967: Delta = 69'sb111111111111111111111111111000000000000000001000000000000000000000000;
		25894: Delta = 69'sb000000000000000000000000000111111111111111111000000000000000000000000;
		38795: Delta = 69'sb111111111111111111111111110111111111111111111000000000000000000000000;
		31046: Delta = 69'sb000000000000000000000000010000000000000000001000000000000000000000000;
		5987: Delta = 69'sb111111111111111111111111110000000000000000001000000000000000000000000;
		44874: Delta = 69'sb000000000000000000000000001111111111111111111000000000000000000000000;
		19815: Delta = 69'sb111111111111111111111111101111111111111111111000000000000000000000000;
		18145: Delta = 69'sb000000000000000000000000100000000000000000001000000000000000000000000;
		18888: Delta = 69'sb111111111111111111111111100000000000000000001000000000000000000000000;
		31973: Delta = 69'sb000000000000000000000000011111111111111111111000000000000000000000000;
		32716: Delta = 69'sb111111111111111111111111011111111111111111111000000000000000000000000;
		43204: Delta = 69'sb000000000000000000000001000000000000000000001000000000000000000000000;
		44690: Delta = 69'sb111111111111111111111111000000000000000000001000000000000000000000000;
		6171: Delta = 69'sb000000000000000000000000111111111111111111111000000000000000000000000;
		7657: Delta = 69'sb111111111111111111111110111111111111111111111000000000000000000000000;
		42461: Delta = 69'sb000000000000000000000010000000000000000000001000000000000000000000000;
		45433: Delta = 69'sb111111111111111111111110000000000000000000001000000000000000000000000;
		5428: Delta = 69'sb000000000000000000000001111111111111111111111000000000000000000000000;
		8400: Delta = 69'sb111111111111111111111101111111111111111111111000000000000000000000000;
		40975: Delta = 69'sb000000000000000000000100000000000000000000001000000000000000000000000;
		46919: Delta = 69'sb111111111111111111111100000000000000000000001000000000000000000000000;
		3942: Delta = 69'sb000000000000000000000011111111111111111111111000000000000000000000000;
		9886: Delta = 69'sb111111111111111111111011111111111111111111111000000000000000000000000;
		38003: Delta = 69'sb000000000000000000001000000000000000000000001000000000000000000000000;
		49891: Delta = 69'sb111111111111111111111000000000000000000000001000000000000000000000000;
		970: Delta = 69'sb000000000000000000000111111111111111111111111000000000000000000000000;
		12858: Delta = 69'sb111111111111111111110111111111111111111111111000000000000000000000000;
		32059: Delta = 69'sb000000000000000000010000000000000000000000001000000000000000000000000;
		4974: Delta = 69'sb111111111111111111110000000000000000000000001000000000000000000000000;
		45887: Delta = 69'sb000000000000000000001111111111111111111111111000000000000000000000000;
		18802: Delta = 69'sb111111111111111111101111111111111111111111111000000000000000000000000;
		20171: Delta = 69'sb000000000000000000100000000000000000000000001000000000000000000000000;
		16862: Delta = 69'sb111111111111111111100000000000000000000000001000000000000000000000000;
		33999: Delta = 69'sb000000000000000000011111111111111111111111111000000000000000000000000;
		30690: Delta = 69'sb111111111111111111011111111111111111111111111000000000000000000000000;
		47256: Delta = 69'sb000000000000000001000000000000000000000000001000000000000000000000000;
		40638: Delta = 69'sb111111111111111111000000000000000000000000001000000000000000000000000;
		10223: Delta = 69'sb000000000000000000111111111111111111111111111000000000000000000000000;
		3605: Delta = 69'sb111111111111111110111111111111111111111111111000000000000000000000000;
		50565: Delta = 69'sb000000000000000010000000000000000000000000001000000000000000000000000;
		37329: Delta = 69'sb111111111111111110000000000000000000000000001000000000000000000000000;
		13532: Delta = 69'sb000000000000000001111111111111111111111111111000000000000000000000000;
		296: Delta = 69'sb111111111111111101111111111111111111111111111000000000000000000000000;
		6322: Delta = 69'sb000000000000000100000000000000000000000000001000000000000000000000000;
		30711: Delta = 69'sb111111111111111100000000000000000000000000001000000000000000000000000;
		20150: Delta = 69'sb000000000000000011111111111111111111111111111000000000000000000000000;
		44539: Delta = 69'sb111111111111111011111111111111111111111111111000000000000000000000000;
		19558: Delta = 69'sb000000000000001000000000000000000000000000001000000000000000000000000;
		17475: Delta = 69'sb111111111111111000000000000000000000000000001000000000000000000000000;
		33386: Delta = 69'sb000000000000000111111111111111111111111111111000000000000000000000000;
		31303: Delta = 69'sb111111111111110111111111111111111111111111111000000000000000000000000;
		46030: Delta = 69'sb000000000000010000000000000000000000000000001000000000000000000000000;
		41864: Delta = 69'sb111111111111110000000000000000000000000000001000000000000000000000000;
		8997: Delta = 69'sb000000000000001111111111111111111111111111111000000000000000000000000;
		4831: Delta = 69'sb111111111111101111111111111111111111111111111000000000000000000000000;
		48113: Delta = 69'sb000000000000100000000000000000000000000000001000000000000000000000000;
		39781: Delta = 69'sb111111111111100000000000000000000000000000001000000000000000000000000;
		11080: Delta = 69'sb000000000000011111111111111111111111111111111000000000000000000000000;
		2748: Delta = 69'sb111111111111011111111111111111111111111111111000000000000000000000000;
		1418: Delta = 69'sb000000000001000000000000000000000000000000001000000000000000000000000;
		35615: Delta = 69'sb111111111111000000000000000000000000000000001000000000000000000000000;
		15246: Delta = 69'sb000000000000111111111111111111111111111111111000000000000000000000000;
		49443: Delta = 69'sb111111111110111111111111111111111111111111111000000000000000000000000;
		9750: Delta = 69'sb000000000010000000000000000000000000000000001000000000000000000000000;
		27283: Delta = 69'sb111111111110000000000000000000000000000000001000000000000000000000000;
		23578: Delta = 69'sb000000000001111111111111111111111111111111111000000000000000000000000;
		41111: Delta = 69'sb111111111101111111111111111111111111111111111000000000000000000000000;
		26414: Delta = 69'sb000000000100000000000000000000000000000000001000000000000000000000000;
		10619: Delta = 69'sb111111111100000000000000000000000000000000001000000000000000000000000;
		40242: Delta = 69'sb000000000011111111111111111111111111111111111000000000000000000000000;
		24447: Delta = 69'sb111111111011111111111111111111111111111111111000000000000000000000000;
		8881: Delta = 69'sb000000001000000000000000000000000000000000001000000000000000000000000;
		28152: Delta = 69'sb111111111000000000000000000000000000000000001000000000000000000000000;
		22709: Delta = 69'sb000000000111111111111111111111111111111111111000000000000000000000000;
		41980: Delta = 69'sb111111110111111111111111111111111111111111111000000000000000000000000;
		24676: Delta = 69'sb000000010000000000000000000000000000000000001000000000000000000000000;
		12357: Delta = 69'sb111111110000000000000000000000000000000000001000000000000000000000000;
		38504: Delta = 69'sb000000001111111111111111111111111111111111111000000000000000000000000;
		26185: Delta = 69'sb111111101111111111111111111111111111111111111000000000000000000000000;
		5405: Delta = 69'sb000000100000000000000000000000000000000000001000000000000000000000000;
		31628: Delta = 69'sb111111100000000000000000000000000000000000001000000000000000000000000;
		19233: Delta = 69'sb000000011111111111111111111111111111111111111000000000000000000000000;
		45456: Delta = 69'sb111111011111111111111111111111111111111111111000000000000000000000000;
		17724: Delta = 69'sb000001000000000000000000000000000000000000001000000000000000000000000;
		19309: Delta = 69'sb111111000000000000000000000000000000000000001000000000000000000000000;
		31552: Delta = 69'sb000000111111111111111111111111111111111111111000000000000000000000000;
		33137: Delta = 69'sb111110111111111111111111111111111111111111111000000000000000000000000;
		42362: Delta = 69'sb000010000000000000000000000000000000000000001000000000000000000000000;
		45532: Delta = 69'sb111110000000000000000000000000000000000000001000000000000000000000000;
		5329: Delta = 69'sb000001111111111111111111111111111111111111111000000000000000000000000;
		8499: Delta = 69'sb111101111111111111111111111111111111111111111000000000000000000000000;
		40777: Delta = 69'sb000100000000000000000000000000000000000000001000000000000000000000000;
		47117: Delta = 69'sb111100000000000000000000000000000000000000001000000000000000000000000;
		3744: Delta = 69'sb000011111111111111111111111111111111111111111000000000000000000000000;
		10084: Delta = 69'sb111011111111111111111111111111111111111111111000000000000000000000000;
		37607: Delta = 69'sb001000000000000000000000000000000000000000001000000000000000000000000;
		50287: Delta = 69'sb111000000000000000000000000000000000000000001000000000000000000000000;
		574: Delta = 69'sb000111111111111111111111111111111111111111111000000000000000000000000;
		13254: Delta = 69'sb110111111111111111111111111111111111111111111000000000000000000000000;
		31267: Delta = 69'sb010000000000000000000000000000000000000000001000000000000000000000000;
		5766: Delta = 69'sb110000000000000000000000000000000000000000001000000000000000000000000;
		45095: Delta = 69'sb001111111111111111111111111111111111111111111000000000000000000000000;
		19594: Delta = 69'sb101111111111111111111111111111111111111111111000000000000000000000000;
		9377: Delta = 69'sb000000000000000000000000000000000000000000110000000000000000000000000;
		41484: Delta = 69'sb111111111111111111111111111111111111111111010000000000000000000000000;
		32582: Delta = 69'sb000000000000000000000000000000000000000001010000000000000000000000000;
		18279: Delta = 69'sb111111111111111111111111111111111111111110110000000000000000000000000;
		28131: Delta = 69'sb000000000000000000000000000000000000000010010000000000000000000000000;
		45935: Delta = 69'sb111111111111111111111111111111111111111110010000000000000000000000000;
		4926: Delta = 69'sb000000000000000000000000000000000000000001110000000000000000000000000;
		22730: Delta = 69'sb111111111111111111111111111111111111111101110000000000000000000000000;
		19229: Delta = 69'sb000000000000000000000000000000000000000100010000000000000000000000000;
		3976: Delta = 69'sb111111111111111111111111111111111111111100010000000000000000000000000;
		46885: Delta = 69'sb000000000000000000000000000000000000000011110000000000000000000000000;
		31632: Delta = 69'sb111111111111111111111111111111111111111011110000000000000000000000000;
		1425: Delta = 69'sb000000000000000000000000000000000000001000010000000000000000000000000;
		21780: Delta = 69'sb111111111111111111111111111111111111111000010000000000000000000000000;
		29081: Delta = 69'sb000000000000000000000000000000000000000111110000000000000000000000000;
		49436: Delta = 69'sb111111111111111111111111111111111111110111110000000000000000000000000;
		16678: Delta = 69'sb000000000000000000000000000000000000010000010000000000000000000000000;
		6527: Delta = 69'sb111111111111111111111111111111111111110000010000000000000000000000000;
		44334: Delta = 69'sb000000000000000000000000000000000000001111110000000000000000000000000;
		34183: Delta = 69'sb111111111111111111111111111111111111101111110000000000000000000000000;
		47184: Delta = 69'sb000000000000000000000000000000000000100000010000000000000000000000000;
		26882: Delta = 69'sb111111111111111111111111111111111111100000010000000000000000000000000;
		23979: Delta = 69'sb000000000000000000000000000000000000011111110000000000000000000000000;
		3677: Delta = 69'sb111111111111111111111111111111111111011111110000000000000000000000000;
		6474: Delta = 69'sb000000000000000000000000000000000001000000010000000000000000000000000;
		16731: Delta = 69'sb111111111111111111111111111111111111000000010000000000000000000000000;
		34130: Delta = 69'sb000000000000000000000000000000000000111111110000000000000000000000000;
		44387: Delta = 69'sb111111111111111111111111111111111110111111110000000000000000000000000;
		26776: Delta = 69'sb000000000000000000000000000000000010000000010000000000000000000000000;
		47290: Delta = 69'sb111111111111111111111111111111111110000000010000000000000000000000000;
		3571: Delta = 69'sb000000000000000000000000000000000001111111110000000000000000000000000;
		24085: Delta = 69'sb111111111111111111111111111111111101111111110000000000000000000000000;
		16519: Delta = 69'sb000000000000000000000000000000000100000000010000000000000000000000000;
		6686: Delta = 69'sb111111111111111111111111111111111100000000010000000000000000000000000;
		44175: Delta = 69'sb000000000000000000000000000000000011111111110000000000000000000000000;
		34342: Delta = 69'sb111111111111111111111111111111111011111111110000000000000000000000000;
		46866: Delta = 69'sb000000000000000000000000000000001000000000010000000000000000000000000;
		27200: Delta = 69'sb111111111111111111111111111111111000000000010000000000000000000000000;
		23661: Delta = 69'sb000000000000000000000000000000000111111111110000000000000000000000000;
		3995: Delta = 69'sb111111111111111111111111111111110111111111110000000000000000000000000;
		5838: Delta = 69'sb000000000000000000000000000000010000000000010000000000000000000000000;
		17367: Delta = 69'sb111111111111111111111111111111110000000000010000000000000000000000000;
		33494: Delta = 69'sb000000000000000000000000000000001111111111110000000000000000000000000;
		45023: Delta = 69'sb111111111111111111111111111111101111111111110000000000000000000000000;
		25504: Delta = 69'sb000000000000000000000000000000100000000000010000000000000000000000000;
		48562: Delta = 69'sb111111111111111111111111111111100000000000010000000000000000000000000;
		2299: Delta = 69'sb000000000000000000000000000000011111111111110000000000000000000000000;
		25357: Delta = 69'sb111111111111111111111111111111011111111111110000000000000000000000000;
		13975: Delta = 69'sb000000000000000000000000000001000000000000010000000000000000000000000;
		9230: Delta = 69'sb111111111111111111111111111111000000000000010000000000000000000000000;
		41631: Delta = 69'sb000000000000000000000000000000111111111111110000000000000000000000000;
		36886: Delta = 69'sb111111111111111111111111111110111111111111110000000000000000000000000;
		41778: Delta = 69'sb000000000000000000000000000010000000000000010000000000000000000000000;
		32288: Delta = 69'sb111111111111111111111111111110000000000000010000000000000000000000000;
		18573: Delta = 69'sb000000000000000000000000000001111111111111110000000000000000000000000;
		9083: Delta = 69'sb111111111111111111111111111101111111111111110000000000000000000000000;
		46523: Delta = 69'sb000000000000000000000000000100000000000000010000000000000000000000000;
		27543: Delta = 69'sb111111111111111111111111111100000000000000010000000000000000000000000;
		23318: Delta = 69'sb000000000000000000000000000011111111111111110000000000000000000000000;
		4338: Delta = 69'sb111111111111111111111111111011111111111111110000000000000000000000000;
		5152: Delta = 69'sb000000000000000000000000001000000000000000010000000000000000000000000;
		18053: Delta = 69'sb111111111111111111111111111000000000000000010000000000000000000000000;
		32808: Delta = 69'sb000000000000000000000000000111111111111111110000000000000000000000000;
		45709: Delta = 69'sb111111111111111111111111110111111111111111110000000000000000000000000;
		24132: Delta = 69'sb000000000000000000000000010000000000000000010000000000000000000000000;
		49934: Delta = 69'sb111111111111111111111111110000000000000000010000000000000000000000000;
		927: Delta = 69'sb000000000000000000000000001111111111111111110000000000000000000000000;
		26729: Delta = 69'sb111111111111111111111111101111111111111111110000000000000000000000000;
		11231: Delta = 69'sb000000000000000000000000100000000000000000010000000000000000000000000;
		11974: Delta = 69'sb111111111111111111111111100000000000000000010000000000000000000000000;
		38887: Delta = 69'sb000000000000000000000000011111111111111111110000000000000000000000000;
		39630: Delta = 69'sb111111111111111111111111011111111111111111110000000000000000000000000;
		36290: Delta = 69'sb000000000000000000000001000000000000000000010000000000000000000000000;
		37776: Delta = 69'sb111111111111111111111111000000000000000000010000000000000000000000000;
		13085: Delta = 69'sb000000000000000000000000111111111111111111110000000000000000000000000;
		14571: Delta = 69'sb111111111111111111111110111111111111111111110000000000000000000000000;
		35547: Delta = 69'sb000000000000000000000010000000000000000000010000000000000000000000000;
		38519: Delta = 69'sb111111111111111111111110000000000000000000010000000000000000000000000;
		12342: Delta = 69'sb000000000000000000000001111111111111111111110000000000000000000000000;
		15314: Delta = 69'sb111111111111111111111101111111111111111111110000000000000000000000000;
		34061: Delta = 69'sb000000000000000000000100000000000000000000010000000000000000000000000;
		40005: Delta = 69'sb111111111111111111111100000000000000000000010000000000000000000000000;
		10856: Delta = 69'sb000000000000000000000011111111111111111111110000000000000000000000000;
		16800: Delta = 69'sb111111111111111111111011111111111111111111110000000000000000000000000;
		31089: Delta = 69'sb000000000000000000001000000000000000000000010000000000000000000000000;
		42977: Delta = 69'sb111111111111111111111000000000000000000000010000000000000000000000000;
		7884: Delta = 69'sb000000000000000000000111111111111111111111110000000000000000000000000;
		19772: Delta = 69'sb111111111111111111110111111111111111111111110000000000000000000000000;
		25145: Delta = 69'sb000000000000000000010000000000000000000000010000000000000000000000000;
		48921: Delta = 69'sb111111111111111111110000000000000000000000010000000000000000000000000;
		1940: Delta = 69'sb000000000000000000001111111111111111111111110000000000000000000000000;
		25716: Delta = 69'sb111111111111111111101111111111111111111111110000000000000000000000000;
		13257: Delta = 69'sb000000000000000000100000000000000000000000010000000000000000000000000;
		9948: Delta = 69'sb111111111111111111100000000000000000000000010000000000000000000000000;
		40913: Delta = 69'sb000000000000000000011111111111111111111111110000000000000000000000000;
		37604: Delta = 69'sb111111111111111111011111111111111111111111110000000000000000000000000;
		40342: Delta = 69'sb000000000000000001000000000000000000000000010000000000000000000000000;
		33724: Delta = 69'sb111111111111111111000000000000000000000000010000000000000000000000000;
		17137: Delta = 69'sb000000000000000000111111111111111111111111110000000000000000000000000;
		10519: Delta = 69'sb111111111111111110111111111111111111111111110000000000000000000000000;
		43651: Delta = 69'sb000000000000000010000000000000000000000000010000000000000000000000000;
		30415: Delta = 69'sb111111111111111110000000000000000000000000010000000000000000000000000;
		20446: Delta = 69'sb000000000000000001111111111111111111111111110000000000000000000000000;
		7210: Delta = 69'sb111111111111111101111111111111111111111111110000000000000000000000000;
		50269: Delta = 69'sb000000000000000100000000000000000000000000010000000000000000000000000;
		23797: Delta = 69'sb111111111111111100000000000000000000000000010000000000000000000000000;
		27064: Delta = 69'sb000000000000000011111111111111111111111111110000000000000000000000000;
		592: Delta = 69'sb111111111111111011111111111111111111111111110000000000000000000000000;
		12644: Delta = 69'sb000000000000001000000000000000000000000000010000000000000000000000000;
		10561: Delta = 69'sb111111111111111000000000000000000000000000010000000000000000000000000;
		40300: Delta = 69'sb000000000000000111111111111111111111111111110000000000000000000000000;
		38217: Delta = 69'sb111111111111110111111111111111111111111111110000000000000000000000000;
		39116: Delta = 69'sb000000000000010000000000000000000000000000010000000000000000000000000;
		34950: Delta = 69'sb111111111111110000000000000000000000000000010000000000000000000000000;
		15911: Delta = 69'sb000000000000001111111111111111111111111111110000000000000000000000000;
		11745: Delta = 69'sb111111111111101111111111111111111111111111110000000000000000000000000;
		41199: Delta = 69'sb000000000000100000000000000000000000000000010000000000000000000000000;
		32867: Delta = 69'sb111111111111100000000000000000000000000000010000000000000000000000000;
		17994: Delta = 69'sb000000000000011111111111111111111111111111110000000000000000000000000;
		9662: Delta = 69'sb111111111111011111111111111111111111111111110000000000000000000000000;
		45365: Delta = 69'sb000000000001000000000000000000000000000000010000000000000000000000000;
		28701: Delta = 69'sb111111111111000000000000000000000000000000010000000000000000000000000;
		22160: Delta = 69'sb000000000000111111111111111111111111111111110000000000000000000000000;
		5496: Delta = 69'sb111111111110111111111111111111111111111111110000000000000000000000000;
		2836: Delta = 69'sb000000000010000000000000000000000000000000010000000000000000000000000;
		20369: Delta = 69'sb111111111110000000000000000000000000000000010000000000000000000000000;
		30492: Delta = 69'sb000000000001111111111111111111111111111111110000000000000000000000000;
		48025: Delta = 69'sb111111111101111111111111111111111111111111110000000000000000000000000;
		19500: Delta = 69'sb000000000100000000000000000000000000000000010000000000000000000000000;
		3705: Delta = 69'sb111111111100000000000000000000000000000000010000000000000000000000000;
		47156: Delta = 69'sb000000000011111111111111111111111111111111110000000000000000000000000;
		31361: Delta = 69'sb111111111011111111111111111111111111111111110000000000000000000000000;
		1967: Delta = 69'sb000000001000000000000000000000000000000000010000000000000000000000000;
		21238: Delta = 69'sb111111111000000000000000000000000000000000010000000000000000000000000;
		29623: Delta = 69'sb000000000111111111111111111111111111111111110000000000000000000000000;
		48894: Delta = 69'sb111111110111111111111111111111111111111111110000000000000000000000000;
		17762: Delta = 69'sb000000010000000000000000000000000000000000010000000000000000000000000;
		5443: Delta = 69'sb111111110000000000000000000000000000000000010000000000000000000000000;
		45418: Delta = 69'sb000000001111111111111111111111111111111111110000000000000000000000000;
		33099: Delta = 69'sb111111101111111111111111111111111111111111110000000000000000000000000;
		49352: Delta = 69'sb000000100000000000000000000000000000000000010000000000000000000000000;
		24714: Delta = 69'sb111111100000000000000000000000000000000000010000000000000000000000000;
		26147: Delta = 69'sb000000011111111111111111111111111111111111110000000000000000000000000;
		1509: Delta = 69'sb111111011111111111111111111111111111111111110000000000000000000000000;
		10810: Delta = 69'sb000001000000000000000000000000000000000000010000000000000000000000000;
		12395: Delta = 69'sb111111000000000000000000000000000000000000010000000000000000000000000;
		38466: Delta = 69'sb000000111111111111111111111111111111111111110000000000000000000000000;
		40051: Delta = 69'sb111110111111111111111111111111111111111111110000000000000000000000000;
		35448: Delta = 69'sb000010000000000000000000000000000000000000010000000000000000000000000;
		38618: Delta = 69'sb111110000000000000000000000000000000000000010000000000000000000000000;
		12243: Delta = 69'sb000001111111111111111111111111111111111111110000000000000000000000000;
		15413: Delta = 69'sb111101111111111111111111111111111111111111110000000000000000000000000;
		33863: Delta = 69'sb000100000000000000000000000000000000000000010000000000000000000000000;
		40203: Delta = 69'sb111100000000000000000000000000000000000000010000000000000000000000000;
		10658: Delta = 69'sb000011111111111111111111111111111111111111110000000000000000000000000;
		16998: Delta = 69'sb111011111111111111111111111111111111111111110000000000000000000000000;
		30693: Delta = 69'sb001000000000000000000000000000000000000000010000000000000000000000000;
		43373: Delta = 69'sb111000000000000000000000000000000000000000010000000000000000000000000;
		7488: Delta = 69'sb000111111111111111111111111111111111111111110000000000000000000000000;
		20168: Delta = 69'sb110111111111111111111111111111111111111111110000000000000000000000000;
		24353: Delta = 69'sb010000000000000000000000000000000000000000010000000000000000000000000;
		49713: Delta = 69'sb110000000000000000000000000000000000000000010000000000000000000000000;
		1148: Delta = 69'sb001111111111111111111111111111111111111111110000000000000000000000000;
		26508: Delta = 69'sb101111111111111111111111111111111111111111110000000000000000000000000;
		18754: Delta = 69'sb000000000000000000000000000000000000000001100000000000000000000000000;
		32107: Delta = 69'sb111111111111111111111111111111111111111110100000000000000000000000000;
		14303: Delta = 69'sb000000000000000000000000000000000000000010100000000000000000000000000;
		36558: Delta = 69'sb111111111111111111111111111111111111111101100000000000000000000000000;
		5401: Delta = 69'sb000000000000000000000000000000000000000100100000000000000000000000000;
		41009: Delta = 69'sb111111111111111111111111111111111111111100100000000000000000000000000;
		9852: Delta = 69'sb000000000000000000000000000000000000000011100000000000000000000000000;
		45460: Delta = 69'sb111111111111111111111111111111111111111011100000000000000000000000000;
		38458: Delta = 69'sb000000000000000000000000000000000000001000100000000000000000000000000;
		7952: Delta = 69'sb111111111111111111111111111111111111111000100000000000000000000000000;
		42909: Delta = 69'sb000000000000000000000000000000000000000111100000000000000000000000000;
		12403: Delta = 69'sb111111111111111111111111111111111111110111100000000000000000000000000;
		2850: Delta = 69'sb000000000000000000000000000000000000010000100000000000000000000000000;
		43560: Delta = 69'sb111111111111111111111111111111111111110000100000000000000000000000000;
		7301: Delta = 69'sb000000000000000000000000000000000000001111100000000000000000000000000;
		48011: Delta = 69'sb111111111111111111111111111111111111101111100000000000000000000000000;
		33356: Delta = 69'sb000000000000000000000000000000000000100000100000000000000000000000000;
		13054: Delta = 69'sb111111111111111111111111111111111111100000100000000000000000000000000;
		37807: Delta = 69'sb000000000000000000000000000000000000011111100000000000000000000000000;
		17505: Delta = 69'sb111111111111111111111111111111111111011111100000000000000000000000000;
		43507: Delta = 69'sb000000000000000000000000000000000001000000100000000000000000000000000;
		2903: Delta = 69'sb111111111111111111111111111111111111000000100000000000000000000000000;
		47958: Delta = 69'sb000000000000000000000000000000000000111111100000000000000000000000000;
		7354: Delta = 69'sb111111111111111111111111111111111110111111100000000000000000000000000;
		12948: Delta = 69'sb000000000000000000000000000000000010000000100000000000000000000000000;
		33462: Delta = 69'sb111111111111111111111111111111111110000000100000000000000000000000000;
		17399: Delta = 69'sb000000000000000000000000000000000001111111100000000000000000000000000;
		37913: Delta = 69'sb111111111111111111111111111111111101111111100000000000000000000000000;
		2691: Delta = 69'sb000000000000000000000000000000000100000000100000000000000000000000000;
		43719: Delta = 69'sb111111111111111111111111111111111100000000100000000000000000000000000;
		7142: Delta = 69'sb000000000000000000000000000000000011111111100000000000000000000000000;
		48170: Delta = 69'sb111111111111111111111111111111111011111111100000000000000000000000000;
		33038: Delta = 69'sb000000000000000000000000000000001000000000100000000000000000000000000;
		13372: Delta = 69'sb111111111111111111111111111111111000000000100000000000000000000000000;
		37489: Delta = 69'sb000000000000000000000000000000000111111111100000000000000000000000000;
		17823: Delta = 69'sb111111111111111111111111111111110111111111100000000000000000000000000;
		42871: Delta = 69'sb000000000000000000000000000000010000000000100000000000000000000000000;
		3539: Delta = 69'sb111111111111111111111111111111110000000000100000000000000000000000000;
		47322: Delta = 69'sb000000000000000000000000000000001111111111100000000000000000000000000;
		7990: Delta = 69'sb111111111111111111111111111111101111111111100000000000000000000000000;
		11676: Delta = 69'sb000000000000000000000000000000100000000000100000000000000000000000000;
		34734: Delta = 69'sb111111111111111111111111111111100000000000100000000000000000000000000;
		16127: Delta = 69'sb000000000000000000000000000000011111111111100000000000000000000000000;
		39185: Delta = 69'sb111111111111111111111111111111011111111111100000000000000000000000000;
		147: Delta = 69'sb000000000000000000000000000001000000000000100000000000000000000000000;
		46263: Delta = 69'sb111111111111111111111111111111000000000000100000000000000000000000000;
		4598: Delta = 69'sb000000000000000000000000000000111111111111100000000000000000000000000;
		50714: Delta = 69'sb111111111111111111111111111110111111111111100000000000000000000000000;
		27950: Delta = 69'sb000000000000000000000000000010000000000000100000000000000000000000000;
		18460: Delta = 69'sb111111111111111111111111111110000000000000100000000000000000000000000;
		32401: Delta = 69'sb000000000000000000000000000001111111111111100000000000000000000000000;
		22911: Delta = 69'sb111111111111111111111111111101111111111111100000000000000000000000000;
		32695: Delta = 69'sb000000000000000000000000000100000000000000100000000000000000000000000;
		13715: Delta = 69'sb111111111111111111111111111100000000000000100000000000000000000000000;
		37146: Delta = 69'sb000000000000000000000000000011111111111111100000000000000000000000000;
		18166: Delta = 69'sb111111111111111111111111111011111111111111100000000000000000000000000;
		42185: Delta = 69'sb000000000000000000000000001000000000000000100000000000000000000000000;
		4225: Delta = 69'sb111111111111111111111111111000000000000000100000000000000000000000000;
		46636: Delta = 69'sb000000000000000000000000000111111111111111100000000000000000000000000;
		8676: Delta = 69'sb111111111111111111111111110111111111111111100000000000000000000000000;
		10304: Delta = 69'sb000000000000000000000000010000000000000000100000000000000000000000000;
		36106: Delta = 69'sb111111111111111111111111110000000000000000100000000000000000000000000;
		14755: Delta = 69'sb000000000000000000000000001111111111111111100000000000000000000000000;
		40557: Delta = 69'sb111111111111111111111111101111111111111111100000000000000000000000000;
		48264: Delta = 69'sb000000000000000000000000100000000000000000100000000000000000000000000;
		49007: Delta = 69'sb111111111111111111111111100000000000000000100000000000000000000000000;
		1854: Delta = 69'sb000000000000000000000000011111111111111111100000000000000000000000000;
		2597: Delta = 69'sb111111111111111111111111011111111111111111100000000000000000000000000;
		22462: Delta = 69'sb000000000000000000000001000000000000000000100000000000000000000000000;
		23948: Delta = 69'sb111111111111111111111111000000000000000000100000000000000000000000000;
		26913: Delta = 69'sb000000000000000000000000111111111111111111100000000000000000000000000;
		28399: Delta = 69'sb111111111111111111111110111111111111111111100000000000000000000000000;
		21719: Delta = 69'sb000000000000000000000010000000000000000000100000000000000000000000000;
		24691: Delta = 69'sb111111111111111111111110000000000000000000100000000000000000000000000;
		26170: Delta = 69'sb000000000000000000000001111111111111111111100000000000000000000000000;
		29142: Delta = 69'sb111111111111111111111101111111111111111111100000000000000000000000000;
		20233: Delta = 69'sb000000000000000000000100000000000000000000100000000000000000000000000;
		26177: Delta = 69'sb111111111111111111111100000000000000000000100000000000000000000000000;
		24684: Delta = 69'sb000000000000000000000011111111111111111111100000000000000000000000000;
		30628: Delta = 69'sb111111111111111111111011111111111111111111100000000000000000000000000;
		17261: Delta = 69'sb000000000000000000001000000000000000000000100000000000000000000000000;
		29149: Delta = 69'sb111111111111111111111000000000000000000000100000000000000000000000000;
		21712: Delta = 69'sb000000000000000000000111111111111111111111100000000000000000000000000;
		33600: Delta = 69'sb111111111111111111110111111111111111111111100000000000000000000000000;
		11317: Delta = 69'sb000000000000000000010000000000000000000000100000000000000000000000000;
		35093: Delta = 69'sb111111111111111111110000000000000000000000100000000000000000000000000;
		15768: Delta = 69'sb000000000000000000001111111111111111111111100000000000000000000000000;
		39544: Delta = 69'sb111111111111111111101111111111111111111111100000000000000000000000000;
		50290: Delta = 69'sb000000000000000000100000000000000000000000100000000000000000000000000;
		46981: Delta = 69'sb111111111111111111100000000000000000000000100000000000000000000000000;
		3880: Delta = 69'sb000000000000000000011111111111111111111111100000000000000000000000000;
		571: Delta = 69'sb111111111111111111011111111111111111111111100000000000000000000000000;
		26514: Delta = 69'sb000000000000000001000000000000000000000000100000000000000000000000000;
		19896: Delta = 69'sb111111111111111111000000000000000000000000100000000000000000000000000;
		30965: Delta = 69'sb000000000000000000111111111111111111111111100000000000000000000000000;
		24347: Delta = 69'sb111111111111111110111111111111111111111111100000000000000000000000000;
		29823: Delta = 69'sb000000000000000010000000000000000000000000100000000000000000000000000;
		16587: Delta = 69'sb111111111111111110000000000000000000000000100000000000000000000000000;
		34274: Delta = 69'sb000000000000000001111111111111111111111111100000000000000000000000000;
		21038: Delta = 69'sb111111111111111101111111111111111111111111100000000000000000000000000;
		36441: Delta = 69'sb000000000000000100000000000000000000000000100000000000000000000000000;
		9969: Delta = 69'sb111111111111111100000000000000000000000000100000000000000000000000000;
		40892: Delta = 69'sb000000000000000011111111111111111111111111100000000000000000000000000;
		14420: Delta = 69'sb111111111111111011111111111111111111111111100000000000000000000000000;
		49677: Delta = 69'sb000000000000001000000000000000000000000000100000000000000000000000000;
		47594: Delta = 69'sb111111111111111000000000000000000000000000100000000000000000000000000;
		3267: Delta = 69'sb000000000000000111111111111111111111111111100000000000000000000000000;
		1184: Delta = 69'sb111111111111110111111111111111111111111111100000000000000000000000000;
		25288: Delta = 69'sb000000000000010000000000000000000000000000100000000000000000000000000;
		21122: Delta = 69'sb111111111111110000000000000000000000000000100000000000000000000000000;
		29739: Delta = 69'sb000000000000001111111111111111111111111111100000000000000000000000000;
		25573: Delta = 69'sb111111111111101111111111111111111111111111100000000000000000000000000;
		27371: Delta = 69'sb000000000000100000000000000000000000000000100000000000000000000000000;
		19039: Delta = 69'sb111111111111100000000000000000000000000000100000000000000000000000000;
		31822: Delta = 69'sb000000000000011111111111111111111111111111100000000000000000000000000;
		23490: Delta = 69'sb111111111111011111111111111111111111111111100000000000000000000000000;
		31537: Delta = 69'sb000000000001000000000000000000000000000000100000000000000000000000000;
		14873: Delta = 69'sb111111111111000000000000000000000000000000100000000000000000000000000;
		35988: Delta = 69'sb000000000000111111111111111111111111111111100000000000000000000000000;
		19324: Delta = 69'sb111111111110111111111111111111111111111111100000000000000000000000000;
		39869: Delta = 69'sb000000000010000000000000000000000000000000100000000000000000000000000;
		6541: Delta = 69'sb111111111110000000000000000000000000000000100000000000000000000000000;
		44320: Delta = 69'sb000000000001111111111111111111111111111111100000000000000000000000000;
		10992: Delta = 69'sb111111111101111111111111111111111111111111100000000000000000000000000;
		5672: Delta = 69'sb000000000100000000000000000000000000000000100000000000000000000000000;
		40738: Delta = 69'sb111111111100000000000000000000000000000000100000000000000000000000000;
		10123: Delta = 69'sb000000000011111111111111111111111111111111100000000000000000000000000;
		45189: Delta = 69'sb111111111011111111111111111111111111111111100000000000000000000000000;
		39000: Delta = 69'sb000000001000000000000000000000000000000000100000000000000000000000000;
		7410: Delta = 69'sb111111111000000000000000000000000000000000100000000000000000000000000;
		43451: Delta = 69'sb000000000111111111111111111111111111111111100000000000000000000000000;
		11861: Delta = 69'sb111111110111111111111111111111111111111111100000000000000000000000000;
		3934: Delta = 69'sb000000010000000000000000000000000000000000100000000000000000000000000;
		42476: Delta = 69'sb111111110000000000000000000000000000000000100000000000000000000000000;
		8385: Delta = 69'sb000000001111111111111111111111111111111111100000000000000000000000000;
		46927: Delta = 69'sb111111101111111111111111111111111111111111100000000000000000000000000;
		35524: Delta = 69'sb000000100000000000000000000000000000000000100000000000000000000000000;
		10886: Delta = 69'sb111111100000000000000000000000000000000000100000000000000000000000000;
		39975: Delta = 69'sb000000011111111111111111111111111111111111100000000000000000000000000;
		15337: Delta = 69'sb111111011111111111111111111111111111111111100000000000000000000000000;
		47843: Delta = 69'sb000001000000000000000000000000000000000000100000000000000000000000000;
		49428: Delta = 69'sb111111000000000000000000000000000000000000100000000000000000000000000;
		1433: Delta = 69'sb000000111111111111111111111111111111111111100000000000000000000000000;
		3018: Delta = 69'sb111110111111111111111111111111111111111111100000000000000000000000000;
		21620: Delta = 69'sb000010000000000000000000000000000000000000100000000000000000000000000;
		24790: Delta = 69'sb111110000000000000000000000000000000000000100000000000000000000000000;
		26071: Delta = 69'sb000001111111111111111111111111111111111111100000000000000000000000000;
		29241: Delta = 69'sb111101111111111111111111111111111111111111100000000000000000000000000;
		20035: Delta = 69'sb000100000000000000000000000000000000000000100000000000000000000000000;
		26375: Delta = 69'sb111100000000000000000000000000000000000000100000000000000000000000000;
		24486: Delta = 69'sb000011111111111111111111111111111111111111100000000000000000000000000;
		30826: Delta = 69'sb111011111111111111111111111111111111111111100000000000000000000000000;
		16865: Delta = 69'sb001000000000000000000000000000000000000000100000000000000000000000000;
		29545: Delta = 69'sb111000000000000000000000000000000000000000100000000000000000000000000;
		21316: Delta = 69'sb000111111111111111111111111111111111111111100000000000000000000000000;
		33996: Delta = 69'sb110111111111111111111111111111111111111111100000000000000000000000000;
		10525: Delta = 69'sb010000000000000000000000000000000000000000100000000000000000000000000;
		35885: Delta = 69'sb110000000000000000000000000000000000000000100000000000000000000000000;
		14976: Delta = 69'sb001111111111111111111111111111111111111111100000000000000000000000000;
		40336: Delta = 69'sb101111111111111111111111111111111111111111100000000000000000000000000;
		37508: Delta = 69'sb000000000000000000000000000000000000000011000000000000000000000000000;
		13353: Delta = 69'sb111111111111111111111111111111111111111101000000000000000000000000000;
		28606: Delta = 69'sb000000000000000000000000000000000000000101000000000000000000000000000;
		22255: Delta = 69'sb111111111111111111111111111111111111111011000000000000000000000000000;
		10802: Delta = 69'sb000000000000000000000000000000000000001001000000000000000000000000000;
		31157: Delta = 69'sb111111111111111111111111111111111111111001000000000000000000000000000;
		19704: Delta = 69'sb000000000000000000000000000000000000000111000000000000000000000000000;
		40059: Delta = 69'sb111111111111111111111111111111111111110111000000000000000000000000000;
		26055: Delta = 69'sb000000000000000000000000000000000000010001000000000000000000000000000;
		15904: Delta = 69'sb111111111111111111111111111111111111110001000000000000000000000000000;
		34957: Delta = 69'sb000000000000000000000000000000000000001111000000000000000000000000000;
		24806: Delta = 69'sb111111111111111111111111111111111111101111000000000000000000000000000;
		5700: Delta = 69'sb000000000000000000000000000000000000100001000000000000000000000000000;
		36259: Delta = 69'sb111111111111111111111111111111111111100001000000000000000000000000000;
		14602: Delta = 69'sb000000000000000000000000000000000000011111000000000000000000000000000;
		45161: Delta = 69'sb111111111111111111111111111111111111011111000000000000000000000000000;
		15851: Delta = 69'sb000000000000000000000000000000000001000001000000000000000000000000000;
		26108: Delta = 69'sb111111111111111111111111111111111111000001000000000000000000000000000;
		24753: Delta = 69'sb000000000000000000000000000000000000111111000000000000000000000000000;
		35010: Delta = 69'sb111111111111111111111111111111111110111111000000000000000000000000000;
		36153: Delta = 69'sb000000000000000000000000000000000010000001000000000000000000000000000;
		5806: Delta = 69'sb111111111111111111111111111111111110000001000000000000000000000000000;
		45055: Delta = 69'sb000000000000000000000000000000000001111111000000000000000000000000000;
		14708: Delta = 69'sb111111111111111111111111111111111101111111000000000000000000000000000;
		25896: Delta = 69'sb000000000000000000000000000000000100000001000000000000000000000000000;
		16063: Delta = 69'sb111111111111111111111111111111111100000001000000000000000000000000000;
		34798: Delta = 69'sb000000000000000000000000000000000011111111000000000000000000000000000;
		24965: Delta = 69'sb111111111111111111111111111111111011111111000000000000000000000000000;
		5382: Delta = 69'sb000000000000000000000000000000001000000001000000000000000000000000000;
		36577: Delta = 69'sb111111111111111111111111111111111000000001000000000000000000000000000;
		14284: Delta = 69'sb000000000000000000000000000000000111111111000000000000000000000000000;
		45479: Delta = 69'sb111111111111111111111111111111110111111111000000000000000000000000000;
		15215: Delta = 69'sb000000000000000000000000000000010000000001000000000000000000000000000;
		26744: Delta = 69'sb111111111111111111111111111111110000000001000000000000000000000000000;
		24117: Delta = 69'sb000000000000000000000000000000001111111111000000000000000000000000000;
		35646: Delta = 69'sb111111111111111111111111111111101111111111000000000000000000000000000;
		34881: Delta = 69'sb000000000000000000000000000000100000000001000000000000000000000000000;
		7078: Delta = 69'sb111111111111111111111111111111100000000001000000000000000000000000000;
		43783: Delta = 69'sb000000000000000000000000000000011111111111000000000000000000000000000;
		15980: Delta = 69'sb111111111111111111111111111111011111111111000000000000000000000000000;
		23352: Delta = 69'sb000000000000000000000000000001000000000001000000000000000000000000000;
		18607: Delta = 69'sb111111111111111111111111111111000000000001000000000000000000000000000;
		32254: Delta = 69'sb000000000000000000000000000000111111111111000000000000000000000000000;
		27509: Delta = 69'sb111111111111111111111111111110111111111111000000000000000000000000000;
		294: Delta = 69'sb000000000000000000000000000010000000000001000000000000000000000000000;
		41665: Delta = 69'sb111111111111111111111111111110000000000001000000000000000000000000000;
		9196: Delta = 69'sb000000000000000000000000000001111111111111000000000000000000000000000;
		50567: Delta = 69'sb111111111111111111111111111101111111111111000000000000000000000000000;
		5039: Delta = 69'sb000000000000000000000000000100000000000001000000000000000000000000000;
		36920: Delta = 69'sb111111111111111111111111111100000000000001000000000000000000000000000;
		13941: Delta = 69'sb000000000000000000000000000011111111111111000000000000000000000000000;
		45822: Delta = 69'sb111111111111111111111111111011111111111111000000000000000000000000000;
		14529: Delta = 69'sb000000000000000000000000001000000000000001000000000000000000000000000;
		27430: Delta = 69'sb111111111111111111111111111000000000000001000000000000000000000000000;
		23431: Delta = 69'sb000000000000000000000000000111111111111111000000000000000000000000000;
		36332: Delta = 69'sb111111111111111111111111110111111111111111000000000000000000000000000;
		33509: Delta = 69'sb000000000000000000000000010000000000000001000000000000000000000000000;
		8450: Delta = 69'sb111111111111111111111111110000000000000001000000000000000000000000000;
		42411: Delta = 69'sb000000000000000000000000001111111111111111000000000000000000000000000;
		17352: Delta = 69'sb111111111111111111111111101111111111111111000000000000000000000000000;
		20608: Delta = 69'sb000000000000000000000000100000000000000001000000000000000000000000000;
		21351: Delta = 69'sb111111111111111111111111100000000000000001000000000000000000000000000;
		29510: Delta = 69'sb000000000000000000000000011111111111111111000000000000000000000000000;
		30253: Delta = 69'sb111111111111111111111111011111111111111111000000000000000000000000000;
		45667: Delta = 69'sb000000000000000000000001000000000000000001000000000000000000000000000;
		47153: Delta = 69'sb111111111111111111111111000000000000000001000000000000000000000000000;
		3708: Delta = 69'sb000000000000000000000000111111111111111111000000000000000000000000000;
		5194: Delta = 69'sb111111111111111111111110111111111111111111000000000000000000000000000;
		44924: Delta = 69'sb000000000000000000000010000000000000000001000000000000000000000000000;
		47896: Delta = 69'sb111111111111111111111110000000000000000001000000000000000000000000000;
		2965: Delta = 69'sb000000000000000000000001111111111111111111000000000000000000000000000;
		5937: Delta = 69'sb111111111111111111111101111111111111111111000000000000000000000000000;
		43438: Delta = 69'sb000000000000000000000100000000000000000001000000000000000000000000000;
		49382: Delta = 69'sb111111111111111111111100000000000000000001000000000000000000000000000;
		1479: Delta = 69'sb000000000000000000000011111111111111111111000000000000000000000000000;
		7423: Delta = 69'sb111111111111111111111011111111111111111111000000000000000000000000000;
		40466: Delta = 69'sb000000000000000000001000000000000000000001000000000000000000000000000;
		1493: Delta = 69'sb111111111111111111111000000000000000000001000000000000000000000000000;
		49368: Delta = 69'sb000000000000000000000111111111111111111111000000000000000000000000000;
		10395: Delta = 69'sb111111111111111111110111111111111111111111000000000000000000000000000;
		34522: Delta = 69'sb000000000000000000010000000000000000000001000000000000000000000000000;
		7437: Delta = 69'sb111111111111111111110000000000000000000001000000000000000000000000000;
		43424: Delta = 69'sb000000000000000000001111111111111111111111000000000000000000000000000;
		16339: Delta = 69'sb111111111111111111101111111111111111111111000000000000000000000000000;
		22634: Delta = 69'sb000000000000000000100000000000000000000001000000000000000000000000000;
		19325: Delta = 69'sb111111111111111111100000000000000000000001000000000000000000000000000;
		31536: Delta = 69'sb000000000000000000011111111111111111111111000000000000000000000000000;
		28227: Delta = 69'sb111111111111111111011111111111111111111111000000000000000000000000000;
		49719: Delta = 69'sb000000000000000001000000000000000000000001000000000000000000000000000;
		43101: Delta = 69'sb111111111111111111000000000000000000000001000000000000000000000000000;
		7760: Delta = 69'sb000000000000000000111111111111111111111111000000000000000000000000000;
		1142: Delta = 69'sb111111111111111110111111111111111111111111000000000000000000000000000;
		2167: Delta = 69'sb000000000000000010000000000000000000000001000000000000000000000000000;
		39792: Delta = 69'sb111111111111111110000000000000000000000001000000000000000000000000000;
		11069: Delta = 69'sb000000000000000001111111111111111111111111000000000000000000000000000;
		48694: Delta = 69'sb111111111111111101111111111111111111111111000000000000000000000000000;
		8785: Delta = 69'sb000000000000000100000000000000000000000001000000000000000000000000000;
		33174: Delta = 69'sb111111111111111100000000000000000000000001000000000000000000000000000;
		17687: Delta = 69'sb000000000000000011111111111111111111111111000000000000000000000000000;
		42076: Delta = 69'sb111111111111111011111111111111111111111111000000000000000000000000000;
		22021: Delta = 69'sb000000000000001000000000000000000000000001000000000000000000000000000;
		19938: Delta = 69'sb111111111111111000000000000000000000000001000000000000000000000000000;
		30923: Delta = 69'sb000000000000000111111111111111111111111111000000000000000000000000000;
		28840: Delta = 69'sb111111111111110111111111111111111111111111000000000000000000000000000;
		48493: Delta = 69'sb000000000000010000000000000000000000000001000000000000000000000000000;
		44327: Delta = 69'sb111111111111110000000000000000000000000001000000000000000000000000000;
		6534: Delta = 69'sb000000000000001111111111111111111111111111000000000000000000000000000;
		2368: Delta = 69'sb111111111111101111111111111111111111111111000000000000000000000000000;
		50576: Delta = 69'sb000000000000100000000000000000000000000001000000000000000000000000000;
		42244: Delta = 69'sb111111111111100000000000000000000000000001000000000000000000000000000;
		8617: Delta = 69'sb000000000000011111111111111111111111111111000000000000000000000000000;
		285: Delta = 69'sb111111111111011111111111111111111111111111000000000000000000000000000;
		3881: Delta = 69'sb000000000001000000000000000000000000000001000000000000000000000000000;
		38078: Delta = 69'sb111111111111000000000000000000000000000001000000000000000000000000000;
		12783: Delta = 69'sb000000000000111111111111111111111111111111000000000000000000000000000;
		46980: Delta = 69'sb111111111110111111111111111111111111111111000000000000000000000000000;
		12213: Delta = 69'sb000000000010000000000000000000000000000001000000000000000000000000000;
		29746: Delta = 69'sb111111111110000000000000000000000000000001000000000000000000000000000;
		21115: Delta = 69'sb000000000001111111111111111111111111111111000000000000000000000000000;
		38648: Delta = 69'sb111111111101111111111111111111111111111111000000000000000000000000000;
		28877: Delta = 69'sb000000000100000000000000000000000000000001000000000000000000000000000;
		13082: Delta = 69'sb111111111100000000000000000000000000000001000000000000000000000000000;
		37779: Delta = 69'sb000000000011111111111111111111111111111111000000000000000000000000000;
		21984: Delta = 69'sb111111111011111111111111111111111111111111000000000000000000000000000;
		11344: Delta = 69'sb000000001000000000000000000000000000000001000000000000000000000000000;
		30615: Delta = 69'sb111111111000000000000000000000000000000001000000000000000000000000000;
		20246: Delta = 69'sb000000000111111111111111111111111111111111000000000000000000000000000;
		39517: Delta = 69'sb111111110111111111111111111111111111111111000000000000000000000000000;
		27139: Delta = 69'sb000000010000000000000000000000000000000001000000000000000000000000000;
		14820: Delta = 69'sb111111110000000000000000000000000000000001000000000000000000000000000;
		36041: Delta = 69'sb000000001111111111111111111111111111111111000000000000000000000000000;
		23722: Delta = 69'sb111111101111111111111111111111111111111111000000000000000000000000000;
		7868: Delta = 69'sb000000100000000000000000000000000000000001000000000000000000000000000;
		34091: Delta = 69'sb111111100000000000000000000000000000000001000000000000000000000000000;
		16770: Delta = 69'sb000000011111111111111111111111111111111111000000000000000000000000000;
		42993: Delta = 69'sb111111011111111111111111111111111111111111000000000000000000000000000;
		20187: Delta = 69'sb000001000000000000000000000000000000000001000000000000000000000000000;
		21772: Delta = 69'sb111111000000000000000000000000000000000001000000000000000000000000000;
		29089: Delta = 69'sb000000111111111111111111111111111111111111000000000000000000000000000;
		30674: Delta = 69'sb111110111111111111111111111111111111111111000000000000000000000000000;
		44825: Delta = 69'sb000010000000000000000000000000000000000001000000000000000000000000000;
		47995: Delta = 69'sb111110000000000000000000000000000000000001000000000000000000000000000;
		2866: Delta = 69'sb000001111111111111111111111111111111111111000000000000000000000000000;
		6036: Delta = 69'sb111101111111111111111111111111111111111111000000000000000000000000000;
		43240: Delta = 69'sb000100000000000000000000000000000000000001000000000000000000000000000;
		49580: Delta = 69'sb111100000000000000000000000000000000000001000000000000000000000000000;
		1281: Delta = 69'sb000011111111111111111111111111111111111111000000000000000000000000000;
		7621: Delta = 69'sb111011111111111111111111111111111111111111000000000000000000000000000;
		40070: Delta = 69'sb001000000000000000000000000000000000000001000000000000000000000000000;
		1889: Delta = 69'sb111000000000000000000000000000000000000001000000000000000000000000000;
		48972: Delta = 69'sb000111111111111111111111111111111111111111000000000000000000000000000;
		10791: Delta = 69'sb110111111111111111111111111111111111111111000000000000000000000000000;
		33730: Delta = 69'sb010000000000000000000000000000000000000001000000000000000000000000000;
		8229: Delta = 69'sb110000000000000000000000000000000000000001000000000000000000000000000;
		42632: Delta = 69'sb001111111111111111111111111111111111111111000000000000000000000000000;
		17131: Delta = 69'sb101111111111111111111111111111111111111111000000000000000000000000000;
		24155: Delta = 69'sb000000000000000000000000000000000000000110000000000000000000000000000;
		26706: Delta = 69'sb111111111111111111111111111111111111111010000000000000000000000000000;
		6351: Delta = 69'sb000000000000000000000000000000000000001010000000000000000000000000000;
		44510: Delta = 69'sb111111111111111111111111111111111111110110000000000000000000000000000;
		21604: Delta = 69'sb000000000000000000000000000000000000010010000000000000000000000000000;
		11453: Delta = 69'sb111111111111111111111111111111111111110010000000000000000000000000000;
		39408: Delta = 69'sb000000000000000000000000000000000000001110000000000000000000000000000;
		29257: Delta = 69'sb111111111111111111111111111111111111101110000000000000000000000000000;
		1249: Delta = 69'sb000000000000000000000000000000000000100010000000000000000000000000000;
		31808: Delta = 69'sb111111111111111111111111111111111111100010000000000000000000000000000;
		19053: Delta = 69'sb000000000000000000000000000000000000011110000000000000000000000000000;
		49612: Delta = 69'sb111111111111111111111111111111111111011110000000000000000000000000000;
		11400: Delta = 69'sb000000000000000000000000000000000001000010000000000000000000000000000;
		21657: Delta = 69'sb111111111111111111111111111111111111000010000000000000000000000000000;
		29204: Delta = 69'sb000000000000000000000000000000000000111110000000000000000000000000000;
		39461: Delta = 69'sb111111111111111111111111111111111110111110000000000000000000000000000;
		31702: Delta = 69'sb000000000000000000000000000000000010000010000000000000000000000000000;
		1355: Delta = 69'sb111111111111111111111111111111111110000010000000000000000000000000000;
		49506: Delta = 69'sb000000000000000000000000000000000001111110000000000000000000000000000;
		19159: Delta = 69'sb111111111111111111111111111111111101111110000000000000000000000000000;
		21445: Delta = 69'sb000000000000000000000000000000000100000010000000000000000000000000000;
		11612: Delta = 69'sb111111111111111111111111111111111100000010000000000000000000000000000;
		39249: Delta = 69'sb000000000000000000000000000000000011111110000000000000000000000000000;
		29416: Delta = 69'sb111111111111111111111111111111111011111110000000000000000000000000000;
		931: Delta = 69'sb000000000000000000000000000000001000000010000000000000000000000000000;
		32126: Delta = 69'sb111111111111111111111111111111111000000010000000000000000000000000000;
		18735: Delta = 69'sb000000000000000000000000000000000111111110000000000000000000000000000;
		49930: Delta = 69'sb111111111111111111111111111111110111111110000000000000000000000000000;
		10764: Delta = 69'sb000000000000000000000000000000010000000010000000000000000000000000000;
		22293: Delta = 69'sb111111111111111111111111111111110000000010000000000000000000000000000;
		28568: Delta = 69'sb000000000000000000000000000000001111111110000000000000000000000000000;
		40097: Delta = 69'sb111111111111111111111111111111101111111110000000000000000000000000000;
		30430: Delta = 69'sb000000000000000000000000000000100000000010000000000000000000000000000;
		2627: Delta = 69'sb111111111111111111111111111111100000000010000000000000000000000000000;
		48234: Delta = 69'sb000000000000000000000000000000011111111110000000000000000000000000000;
		20431: Delta = 69'sb111111111111111111111111111111011111111110000000000000000000000000000;
		18901: Delta = 69'sb000000000000000000000000000001000000000010000000000000000000000000000;
		14156: Delta = 69'sb111111111111111111111111111111000000000010000000000000000000000000000;
		36705: Delta = 69'sb000000000000000000000000000000111111111110000000000000000000000000000;
		31960: Delta = 69'sb111111111111111111111111111110111111111110000000000000000000000000000;
		46704: Delta = 69'sb000000000000000000000000000010000000000010000000000000000000000000000;
		37214: Delta = 69'sb111111111111111111111111111110000000000010000000000000000000000000000;
		13647: Delta = 69'sb000000000000000000000000000001111111111110000000000000000000000000000;
		4157: Delta = 69'sb111111111111111111111111111101111111111110000000000000000000000000000;
		588: Delta = 69'sb000000000000000000000000000100000000000010000000000000000000000000000;
		32469: Delta = 69'sb111111111111111111111111111100000000000010000000000000000000000000000;
		18392: Delta = 69'sb000000000000000000000000000011111111111110000000000000000000000000000;
		50273: Delta = 69'sb111111111111111111111111111011111111111110000000000000000000000000000;
		10078: Delta = 69'sb000000000000000000000000001000000000000010000000000000000000000000000;
		22979: Delta = 69'sb111111111111111111111111111000000000000010000000000000000000000000000;
		27882: Delta = 69'sb000000000000000000000000000111111111111110000000000000000000000000000;
		40783: Delta = 69'sb111111111111111111111111110111111111111110000000000000000000000000000;
		29058: Delta = 69'sb000000000000000000000000010000000000000010000000000000000000000000000;
		3999: Delta = 69'sb111111111111111111111111110000000000000010000000000000000000000000000;
		46862: Delta = 69'sb000000000000000000000000001111111111111110000000000000000000000000000;
		21803: Delta = 69'sb111111111111111111111111101111111111111110000000000000000000000000000;
		16157: Delta = 69'sb000000000000000000000000100000000000000010000000000000000000000000000;
		16900: Delta = 69'sb111111111111111111111111100000000000000010000000000000000000000000000;
		33961: Delta = 69'sb000000000000000000000000011111111111111110000000000000000000000000000;
		34704: Delta = 69'sb111111111111111111111111011111111111111110000000000000000000000000000;
		41216: Delta = 69'sb000000000000000000000001000000000000000010000000000000000000000000000;
		42702: Delta = 69'sb111111111111111111111111000000000000000010000000000000000000000000000;
		8159: Delta = 69'sb000000000000000000000000111111111111111110000000000000000000000000000;
		9645: Delta = 69'sb111111111111111111111110111111111111111110000000000000000000000000000;
		40473: Delta = 69'sb000000000000000000000010000000000000000010000000000000000000000000000;
		43445: Delta = 69'sb111111111111111111111110000000000000000010000000000000000000000000000;
		7416: Delta = 69'sb000000000000000000000001111111111111111110000000000000000000000000000;
		10388: Delta = 69'sb111111111111111111111101111111111111111110000000000000000000000000000;
		38987: Delta = 69'sb000000000000000000000100000000000000000010000000000000000000000000000;
		44931: Delta = 69'sb111111111111111111111100000000000000000010000000000000000000000000000;
		5930: Delta = 69'sb000000000000000000000011111111111111111110000000000000000000000000000;
		11874: Delta = 69'sb111111111111111111111011111111111111111110000000000000000000000000000;
		36015: Delta = 69'sb000000000000000000001000000000000000000010000000000000000000000000000;
		47903: Delta = 69'sb111111111111111111111000000000000000000010000000000000000000000000000;
		2958: Delta = 69'sb000000000000000000000111111111111111111110000000000000000000000000000;
		14846: Delta = 69'sb111111111111111111110111111111111111111110000000000000000000000000000;
		30071: Delta = 69'sb000000000000000000010000000000000000000010000000000000000000000000000;
		2986: Delta = 69'sb111111111111111111110000000000000000000010000000000000000000000000000;
		47875: Delta = 69'sb000000000000000000001111111111111111111110000000000000000000000000000;
		20790: Delta = 69'sb111111111111111111101111111111111111111110000000000000000000000000000;
		18183: Delta = 69'sb000000000000000000100000000000000000000010000000000000000000000000000;
		14874: Delta = 69'sb111111111111111111100000000000000000000010000000000000000000000000000;
		35987: Delta = 69'sb000000000000000000011111111111111111111110000000000000000000000000000;
		32678: Delta = 69'sb111111111111111111011111111111111111111110000000000000000000000000000;
		45268: Delta = 69'sb000000000000000001000000000000000000000010000000000000000000000000000;
		38650: Delta = 69'sb111111111111111111000000000000000000000010000000000000000000000000000;
		12211: Delta = 69'sb000000000000000000111111111111111111111110000000000000000000000000000;
		5593: Delta = 69'sb111111111111111110111111111111111111111110000000000000000000000000000;
		48577: Delta = 69'sb000000000000000010000000000000000000000010000000000000000000000000000;
		35341: Delta = 69'sb111111111111111110000000000000000000000010000000000000000000000000000;
		15520: Delta = 69'sb000000000000000001111111111111111111111110000000000000000000000000000;
		2284: Delta = 69'sb111111111111111101111111111111111111111110000000000000000000000000000;
		4334: Delta = 69'sb000000000000000100000000000000000000000010000000000000000000000000000;
		28723: Delta = 69'sb111111111111111100000000000000000000000010000000000000000000000000000;
		22138: Delta = 69'sb000000000000000011111111111111111111111110000000000000000000000000000;
		46527: Delta = 69'sb111111111111111011111111111111111111111110000000000000000000000000000;
		17570: Delta = 69'sb000000000000001000000000000000000000000010000000000000000000000000000;
		15487: Delta = 69'sb111111111111111000000000000000000000000010000000000000000000000000000;
		35374: Delta = 69'sb000000000000000111111111111111111111111110000000000000000000000000000;
		33291: Delta = 69'sb111111111111110111111111111111111111111110000000000000000000000000000;
		44042: Delta = 69'sb000000000000010000000000000000000000000010000000000000000000000000000;
		39876: Delta = 69'sb111111111111110000000000000000000000000010000000000000000000000000000;
		10985: Delta = 69'sb000000000000001111111111111111111111111110000000000000000000000000000;
		6819: Delta = 69'sb111111111111101111111111111111111111111110000000000000000000000000000;
		46125: Delta = 69'sb000000000000100000000000000000000000000010000000000000000000000000000;
		37793: Delta = 69'sb111111111111100000000000000000000000000010000000000000000000000000000;
		13068: Delta = 69'sb000000000000011111111111111111111111111110000000000000000000000000000;
		4736: Delta = 69'sb111111111111011111111111111111111111111110000000000000000000000000000;
		50291: Delta = 69'sb000000000001000000000000000000000000000010000000000000000000000000000;
		33627: Delta = 69'sb111111111111000000000000000000000000000010000000000000000000000000000;
		17234: Delta = 69'sb000000000000111111111111111111111111111110000000000000000000000000000;
		570: Delta = 69'sb111111111110111111111111111111111111111110000000000000000000000000000;
		7762: Delta = 69'sb000000000010000000000000000000000000000010000000000000000000000000000;
		25295: Delta = 69'sb111111111110000000000000000000000000000010000000000000000000000000000;
		25566: Delta = 69'sb000000000001111111111111111111111111111110000000000000000000000000000;
		43099: Delta = 69'sb111111111101111111111111111111111111111110000000000000000000000000000;
		24426: Delta = 69'sb000000000100000000000000000000000000000010000000000000000000000000000;
		8631: Delta = 69'sb111111111100000000000000000000000000000010000000000000000000000000000;
		42230: Delta = 69'sb000000000011111111111111111111111111111110000000000000000000000000000;
		26435: Delta = 69'sb111111111011111111111111111111111111111110000000000000000000000000000;
		6893: Delta = 69'sb000000001000000000000000000000000000000010000000000000000000000000000;
		26164: Delta = 69'sb111111111000000000000000000000000000000010000000000000000000000000000;
		24697: Delta = 69'sb000000000111111111111111111111111111111110000000000000000000000000000;
		43968: Delta = 69'sb111111110111111111111111111111111111111110000000000000000000000000000;
		22688: Delta = 69'sb000000010000000000000000000000000000000010000000000000000000000000000;
		10369: Delta = 69'sb111111110000000000000000000000000000000010000000000000000000000000000;
		40492: Delta = 69'sb000000001111111111111111111111111111111110000000000000000000000000000;
		28173: Delta = 69'sb111111101111111111111111111111111111111110000000000000000000000000000;
		3417: Delta = 69'sb000000100000000000000000000000000000000010000000000000000000000000000;
		29640: Delta = 69'sb111111100000000000000000000000000000000010000000000000000000000000000;
		21221: Delta = 69'sb000000011111111111111111111111111111111110000000000000000000000000000;
		47444: Delta = 69'sb111111011111111111111111111111111111111110000000000000000000000000000;
		15736: Delta = 69'sb000001000000000000000000000000000000000010000000000000000000000000000;
		17321: Delta = 69'sb111111000000000000000000000000000000000010000000000000000000000000000;
		33540: Delta = 69'sb000000111111111111111111111111111111111110000000000000000000000000000;
		35125: Delta = 69'sb111110111111111111111111111111111111111110000000000000000000000000000;
		40374: Delta = 69'sb000010000000000000000000000000000000000010000000000000000000000000000;
		43544: Delta = 69'sb111110000000000000000000000000000000000010000000000000000000000000000;
		7317: Delta = 69'sb000001111111111111111111111111111111111110000000000000000000000000000;
		10487: Delta = 69'sb111101111111111111111111111111111111111110000000000000000000000000000;
		38789: Delta = 69'sb000100000000000000000000000000000000000010000000000000000000000000000;
		45129: Delta = 69'sb111100000000000000000000000000000000000010000000000000000000000000000;
		5732: Delta = 69'sb000011111111111111111111111111111111111110000000000000000000000000000;
		12072: Delta = 69'sb111011111111111111111111111111111111111110000000000000000000000000000;
		35619: Delta = 69'sb001000000000000000000000000000000000000010000000000000000000000000000;
		48299: Delta = 69'sb111000000000000000000000000000000000000010000000000000000000000000000;
		2562: Delta = 69'sb000111111111111111111111111111111111111110000000000000000000000000000;
		15242: Delta = 69'sb110111111111111111111111111111111111111110000000000000000000000000000;
		29279: Delta = 69'sb010000000000000000000000000000000000000010000000000000000000000000000;
		3778: Delta = 69'sb110000000000000000000000000000000000000010000000000000000000000000000;
		47083: Delta = 69'sb001111111111111111111111111111111111111110000000000000000000000000000;
		21582: Delta = 69'sb101111111111111111111111111111111111111110000000000000000000000000000;
		48310: Delta = 69'sb000000000000000000000000000000000000001100000000000000000000000000000;
		2551: Delta = 69'sb111111111111111111111111111111111111110100000000000000000000000000000;
		12702: Delta = 69'sb000000000000000000000000000000000000010100000000000000000000000000000;
		38159: Delta = 69'sb111111111111111111111111111111111111101100000000000000000000000000000;
		43208: Delta = 69'sb000000000000000000000000000000000000100100000000000000000000000000000;
		22906: Delta = 69'sb111111111111111111111111111111111111100100000000000000000000000000000;
		27955: Delta = 69'sb000000000000000000000000000000000000011100000000000000000000000000000;
		7653: Delta = 69'sb111111111111111111111111111111111111011100000000000000000000000000000;
		2498: Delta = 69'sb000000000000000000000000000000000001000100000000000000000000000000000;
		12755: Delta = 69'sb111111111111111111111111111111111111000100000000000000000000000000000;
		38106: Delta = 69'sb000000000000000000000000000000000000111100000000000000000000000000000;
		48363: Delta = 69'sb111111111111111111111111111111111110111100000000000000000000000000000;
		22800: Delta = 69'sb000000000000000000000000000000000010000100000000000000000000000000000;
		43314: Delta = 69'sb111111111111111111111111111111111110000100000000000000000000000000000;
		7547: Delta = 69'sb000000000000000000000000000000000001111100000000000000000000000000000;
		28061: Delta = 69'sb111111111111111111111111111111111101111100000000000000000000000000000;
		12543: Delta = 69'sb000000000000000000000000000000000100000100000000000000000000000000000;
		2710: Delta = 69'sb111111111111111111111111111111111100000100000000000000000000000000000;
		48151: Delta = 69'sb000000000000000000000000000000000011111100000000000000000000000000000;
		38318: Delta = 69'sb111111111111111111111111111111111011111100000000000000000000000000000;
		42890: Delta = 69'sb000000000000000000000000000000001000000100000000000000000000000000000;
		23224: Delta = 69'sb111111111111111111111111111111111000000100000000000000000000000000000;
		27637: Delta = 69'sb000000000000000000000000000000000111111100000000000000000000000000000;
		7971: Delta = 69'sb111111111111111111111111111111110111111100000000000000000000000000000;
		1862: Delta = 69'sb000000000000000000000000000000010000000100000000000000000000000000000;
		13391: Delta = 69'sb111111111111111111111111111111110000000100000000000000000000000000000;
		37470: Delta = 69'sb000000000000000000000000000000001111111100000000000000000000000000000;
		48999: Delta = 69'sb111111111111111111111111111111101111111100000000000000000000000000000;
		21528: Delta = 69'sb000000000000000000000000000000100000000100000000000000000000000000000;
		44586: Delta = 69'sb111111111111111111111111111111100000000100000000000000000000000000000;
		6275: Delta = 69'sb000000000000000000000000000000011111111100000000000000000000000000000;
		29333: Delta = 69'sb111111111111111111111111111111011111111100000000000000000000000000000;
		9999: Delta = 69'sb000000000000000000000000000001000000000100000000000000000000000000000;
		5254: Delta = 69'sb111111111111111111111111111111000000000100000000000000000000000000000;
		45607: Delta = 69'sb000000000000000000000000000000111111111100000000000000000000000000000;
		40862: Delta = 69'sb111111111111111111111111111110111111111100000000000000000000000000000;
		37802: Delta = 69'sb000000000000000000000000000010000000000100000000000000000000000000000;
		28312: Delta = 69'sb111111111111111111111111111110000000000100000000000000000000000000000;
		22549: Delta = 69'sb000000000000000000000000000001111111111100000000000000000000000000000;
		13059: Delta = 69'sb111111111111111111111111111101111111111100000000000000000000000000000;
		42547: Delta = 69'sb000000000000000000000000000100000000000100000000000000000000000000000;
		23567: Delta = 69'sb111111111111111111111111111100000000000100000000000000000000000000000;
		27294: Delta = 69'sb000000000000000000000000000011111111111100000000000000000000000000000;
		8314: Delta = 69'sb111111111111111111111111111011111111111100000000000000000000000000000;
		1176: Delta = 69'sb000000000000000000000000001000000000000100000000000000000000000000000;
		14077: Delta = 69'sb111111111111111111111111111000000000000100000000000000000000000000000;
		36784: Delta = 69'sb000000000000000000000000000111111111111100000000000000000000000000000;
		49685: Delta = 69'sb111111111111111111111111110111111111111100000000000000000000000000000;
		20156: Delta = 69'sb000000000000000000000000010000000000000100000000000000000000000000000;
		45958: Delta = 69'sb111111111111111111111111110000000000000100000000000000000000000000000;
		4903: Delta = 69'sb000000000000000000000000001111111111111100000000000000000000000000000;
		30705: Delta = 69'sb111111111111111111111111101111111111111100000000000000000000000000000;
		7255: Delta = 69'sb000000000000000000000000100000000000000100000000000000000000000000000;
		7998: Delta = 69'sb111111111111111111111111100000000000000100000000000000000000000000000;
		42863: Delta = 69'sb000000000000000000000000011111111111111100000000000000000000000000000;
		43606: Delta = 69'sb111111111111111111111111011111111111111100000000000000000000000000000;
		32314: Delta = 69'sb000000000000000000000001000000000000000100000000000000000000000000000;
		33800: Delta = 69'sb111111111111111111111111000000000000000100000000000000000000000000000;
		17061: Delta = 69'sb000000000000000000000000111111111111111100000000000000000000000000000;
		18547: Delta = 69'sb111111111111111111111110111111111111111100000000000000000000000000000;
		31571: Delta = 69'sb000000000000000000000010000000000000000100000000000000000000000000000;
		34543: Delta = 69'sb111111111111111111111110000000000000000100000000000000000000000000000;
		16318: Delta = 69'sb000000000000000000000001111111111111111100000000000000000000000000000;
		19290: Delta = 69'sb111111111111111111111101111111111111111100000000000000000000000000000;
		30085: Delta = 69'sb000000000000000000000100000000000000000100000000000000000000000000000;
		36029: Delta = 69'sb111111111111111111111100000000000000000100000000000000000000000000000;
		14832: Delta = 69'sb000000000000000000000011111111111111111100000000000000000000000000000;
		20776: Delta = 69'sb111111111111111111111011111111111111111100000000000000000000000000000;
		27113: Delta = 69'sb000000000000000000001000000000000000000100000000000000000000000000000;
		39001: Delta = 69'sb111111111111111111111000000000000000000100000000000000000000000000000;
		11860: Delta = 69'sb000000000000000000000111111111111111111100000000000000000000000000000;
		23748: Delta = 69'sb111111111111111111110111111111111111111100000000000000000000000000000;
		21169: Delta = 69'sb000000000000000000010000000000000000000100000000000000000000000000000;
		44945: Delta = 69'sb111111111111111111110000000000000000000100000000000000000000000000000;
		5916: Delta = 69'sb000000000000000000001111111111111111111100000000000000000000000000000;
		29692: Delta = 69'sb111111111111111111101111111111111111111100000000000000000000000000000;
		9281: Delta = 69'sb000000000000000000100000000000000000000100000000000000000000000000000;
		5972: Delta = 69'sb111111111111111111100000000000000000000100000000000000000000000000000;
		44889: Delta = 69'sb000000000000000000011111111111111111111100000000000000000000000000000;
		41580: Delta = 69'sb111111111111111111011111111111111111111100000000000000000000000000000;
		36366: Delta = 69'sb000000000000000001000000000000000000000100000000000000000000000000000;
		29748: Delta = 69'sb111111111111111111000000000000000000000100000000000000000000000000000;
		21113: Delta = 69'sb000000000000000000111111111111111111111100000000000000000000000000000;
		14495: Delta = 69'sb111111111111111110111111111111111111111100000000000000000000000000000;
		39675: Delta = 69'sb000000000000000010000000000000000000000100000000000000000000000000000;
		26439: Delta = 69'sb111111111111111110000000000000000000000100000000000000000000000000000;
		24422: Delta = 69'sb000000000000000001111111111111111111111100000000000000000000000000000;
		11186: Delta = 69'sb111111111111111101111111111111111111111100000000000000000000000000000;
		46293: Delta = 69'sb000000000000000100000000000000000000000100000000000000000000000000000;
		19821: Delta = 69'sb111111111111111100000000000000000000000100000000000000000000000000000;
		31040: Delta = 69'sb000000000000000011111111111111111111111100000000000000000000000000000;
		4568: Delta = 69'sb111111111111111011111111111111111111111100000000000000000000000000000;
		8668: Delta = 69'sb000000000000001000000000000000000000000100000000000000000000000000000;
		6585: Delta = 69'sb111111111111111000000000000000000000000100000000000000000000000000000;
		44276: Delta = 69'sb000000000000000111111111111111111111111100000000000000000000000000000;
		42193: Delta = 69'sb111111111111110111111111111111111111111100000000000000000000000000000;
		35140: Delta = 69'sb000000000000010000000000000000000000000100000000000000000000000000000;
		30974: Delta = 69'sb111111111111110000000000000000000000000100000000000000000000000000000;
		19887: Delta = 69'sb000000000000001111111111111111111111111100000000000000000000000000000;
		15721: Delta = 69'sb111111111111101111111111111111111111111100000000000000000000000000000;
		37223: Delta = 69'sb000000000000100000000000000000000000000100000000000000000000000000000;
		28891: Delta = 69'sb111111111111100000000000000000000000000100000000000000000000000000000;
		21970: Delta = 69'sb000000000000011111111111111111111111111100000000000000000000000000000;
		13638: Delta = 69'sb111111111111011111111111111111111111111100000000000000000000000000000;
		41389: Delta = 69'sb000000000001000000000000000000000000000100000000000000000000000000000;
		24725: Delta = 69'sb111111111111000000000000000000000000000100000000000000000000000000000;
		26136: Delta = 69'sb000000000000111111111111111111111111111100000000000000000000000000000;
		9472: Delta = 69'sb111111111110111111111111111111111111111100000000000000000000000000000;
		49721: Delta = 69'sb000000000010000000000000000000000000000100000000000000000000000000000;
		16393: Delta = 69'sb111111111110000000000000000000000000000100000000000000000000000000000;
		34468: Delta = 69'sb000000000001111111111111111111111111111100000000000000000000000000000;
		1140: Delta = 69'sb111111111101111111111111111111111111111100000000000000000000000000000;
		15524: Delta = 69'sb000000000100000000000000000000000000000100000000000000000000000000000;
		50590: Delta = 69'sb111111111100000000000000000000000000000100000000000000000000000000000;
		271: Delta = 69'sb000000000011111111111111111111111111111100000000000000000000000000000;
		35337: Delta = 69'sb111111111011111111111111111111111111111100000000000000000000000000000;
		48852: Delta = 69'sb000000001000000000000000000000000000000100000000000000000000000000000;
		17262: Delta = 69'sb111111111000000000000000000000000000000100000000000000000000000000000;
		33599: Delta = 69'sb000000000111111111111111111111111111111100000000000000000000000000000;
		2009: Delta = 69'sb111111110111111111111111111111111111111100000000000000000000000000000;
		13786: Delta = 69'sb000000010000000000000000000000000000000100000000000000000000000000000;
		1467: Delta = 69'sb111111110000000000000000000000000000000100000000000000000000000000000;
		49394: Delta = 69'sb000000001111111111111111111111111111111100000000000000000000000000000;
		37075: Delta = 69'sb111111101111111111111111111111111111111100000000000000000000000000000;
		45376: Delta = 69'sb000000100000000000000000000000000000000100000000000000000000000000000;
		20738: Delta = 69'sb111111100000000000000000000000000000000100000000000000000000000000000;
		30123: Delta = 69'sb000000011111111111111111111111111111111100000000000000000000000000000;
		5485: Delta = 69'sb111111011111111111111111111111111111111100000000000000000000000000000;
		6834: Delta = 69'sb000001000000000000000000000000000000000100000000000000000000000000000;
		8419: Delta = 69'sb111111000000000000000000000000000000000100000000000000000000000000000;
		42442: Delta = 69'sb000000111111111111111111111111111111111100000000000000000000000000000;
		44027: Delta = 69'sb111110111111111111111111111111111111111100000000000000000000000000000;
		31472: Delta = 69'sb000010000000000000000000000000000000000100000000000000000000000000000;
		34642: Delta = 69'sb111110000000000000000000000000000000000100000000000000000000000000000;
		16219: Delta = 69'sb000001111111111111111111111111111111111100000000000000000000000000000;
		19389: Delta = 69'sb111101111111111111111111111111111111111100000000000000000000000000000;
		29887: Delta = 69'sb000100000000000000000000000000000000000100000000000000000000000000000;
		36227: Delta = 69'sb111100000000000000000000000000000000000100000000000000000000000000000;
		14634: Delta = 69'sb000011111111111111111111111111111111111100000000000000000000000000000;
		20974: Delta = 69'sb111011111111111111111111111111111111111100000000000000000000000000000;
		26717: Delta = 69'sb001000000000000000000000000000000000000100000000000000000000000000000;
		39397: Delta = 69'sb111000000000000000000000000000000000000100000000000000000000000000000;
		11464: Delta = 69'sb000111111111111111111111111111111111111100000000000000000000000000000;
		24144: Delta = 69'sb110111111111111111111111111111111111111100000000000000000000000000000;
		20377: Delta = 69'sb010000000000000000000000000000000000000100000000000000000000000000000;
		45737: Delta = 69'sb110000000000000000000000000000000000000100000000000000000000000000000;
		5124: Delta = 69'sb001111111111111111111111111111111111111100000000000000000000000000000;
		30484: Delta = 69'sb101111111111111111111111111111111111111100000000000000000000000000000;
		45759: Delta = 69'sb000000000000000000000000000000000000011000000000000000000000000000000;
		5102: Delta = 69'sb111111111111111111111111111111111111101000000000000000000000000000000;
		25404: Delta = 69'sb000000000000000000000000000000000000101000000000000000000000000000000;
		25457: Delta = 69'sb111111111111111111111111111111111111011000000000000000000000000000000;
		35555: Delta = 69'sb000000000000000000000000000000000001001000000000000000000000000000000;
		45812: Delta = 69'sb111111111111111111111111111111111111001000000000000000000000000000000;
		5049: Delta = 69'sb000000000000000000000000000000000000111000000000000000000000000000000;
		15306: Delta = 69'sb111111111111111111111111111111111110111000000000000000000000000000000;
		4996: Delta = 69'sb000000000000000000000000000000000010001000000000000000000000000000000;
		25510: Delta = 69'sb111111111111111111111111111111111110001000000000000000000000000000000;
		25351: Delta = 69'sb000000000000000000000000000000000001111000000000000000000000000000000;
		45865: Delta = 69'sb111111111111111111111111111111111101111000000000000000000000000000000;
		45600: Delta = 69'sb000000000000000000000000000000000100001000000000000000000000000000000;
		35767: Delta = 69'sb111111111111111111111111111111111100001000000000000000000000000000000;
		15094: Delta = 69'sb000000000000000000000000000000000011111000000000000000000000000000000;
		5261: Delta = 69'sb111111111111111111111111111111111011111000000000000000000000000000000;
		25086: Delta = 69'sb000000000000000000000000000000001000001000000000000000000000000000000;
		5420: Delta = 69'sb111111111111111111111111111111111000001000000000000000000000000000000;
		45441: Delta = 69'sb000000000000000000000000000000000111111000000000000000000000000000000;
		25775: Delta = 69'sb111111111111111111111111111111110111111000000000000000000000000000000;
		34919: Delta = 69'sb000000000000000000000000000000010000001000000000000000000000000000000;
		46448: Delta = 69'sb111111111111111111111111111111110000001000000000000000000000000000000;
		4413: Delta = 69'sb000000000000000000000000000000001111111000000000000000000000000000000;
		15942: Delta = 69'sb111111111111111111111111111111101111111000000000000000000000000000000;
		3724: Delta = 69'sb000000000000000000000000000000100000001000000000000000000000000000000;
		26782: Delta = 69'sb111111111111111111111111111111100000001000000000000000000000000000000;
		24079: Delta = 69'sb000000000000000000000000000000011111111000000000000000000000000000000;
		47137: Delta = 69'sb111111111111111111111111111111011111111000000000000000000000000000000;
		43056: Delta = 69'sb000000000000000000000000000001000000001000000000000000000000000000000;
		38311: Delta = 69'sb111111111111111111111111111111000000001000000000000000000000000000000;
		12550: Delta = 69'sb000000000000000000000000000000111111111000000000000000000000000000000;
		7805: Delta = 69'sb111111111111111111111111111110111111111000000000000000000000000000000;
		19998: Delta = 69'sb000000000000000000000000000010000000001000000000000000000000000000000;
		10508: Delta = 69'sb111111111111111111111111111110000000001000000000000000000000000000000;
		40353: Delta = 69'sb000000000000000000000000000001111111111000000000000000000000000000000;
		30863: Delta = 69'sb111111111111111111111111111101111111111000000000000000000000000000000;
		24743: Delta = 69'sb000000000000000000000000000100000000001000000000000000000000000000000;
		5763: Delta = 69'sb111111111111111111111111111100000000001000000000000000000000000000000;
		45098: Delta = 69'sb000000000000000000000000000011111111111000000000000000000000000000000;
		26118: Delta = 69'sb111111111111111111111111111011111111111000000000000000000000000000000;
		34233: Delta = 69'sb000000000000000000000000001000000000001000000000000000000000000000000;
		47134: Delta = 69'sb111111111111111111111111111000000000001000000000000000000000000000000;
		3727: Delta = 69'sb000000000000000000000000000111111111111000000000000000000000000000000;
		16628: Delta = 69'sb111111111111111111111111110111111111111000000000000000000000000000000;
		2352: Delta = 69'sb000000000000000000000000010000000000001000000000000000000000000000000;
		28154: Delta = 69'sb111111111111111111111111110000000000001000000000000000000000000000000;
		22707: Delta = 69'sb000000000000000000000000001111111111111000000000000000000000000000000;
		48509: Delta = 69'sb111111111111111111111111101111111111111000000000000000000000000000000;
		40312: Delta = 69'sb000000000000000000000000100000000000001000000000000000000000000000000;
		41055: Delta = 69'sb111111111111111111111111100000000000001000000000000000000000000000000;
		9806: Delta = 69'sb000000000000000000000000011111111111111000000000000000000000000000000;
		10549: Delta = 69'sb111111111111111111111111011111111111111000000000000000000000000000000;
		14510: Delta = 69'sb000000000000000000000001000000000000001000000000000000000000000000000;
		15996: Delta = 69'sb111111111111111111111111000000000000001000000000000000000000000000000;
		34865: Delta = 69'sb000000000000000000000000111111111111111000000000000000000000000000000;
		36351: Delta = 69'sb111111111111111111111110111111111111111000000000000000000000000000000;
		13767: Delta = 69'sb000000000000000000000010000000000000001000000000000000000000000000000;
		16739: Delta = 69'sb111111111111111111111110000000000000001000000000000000000000000000000;
		34122: Delta = 69'sb000000000000000000000001111111111111111000000000000000000000000000000;
		37094: Delta = 69'sb111111111111111111111101111111111111111000000000000000000000000000000;
		12281: Delta = 69'sb000000000000000000000100000000000000001000000000000000000000000000000;
		18225: Delta = 69'sb111111111111111111111100000000000000001000000000000000000000000000000;
		32636: Delta = 69'sb000000000000000000000011111111111111111000000000000000000000000000000;
		38580: Delta = 69'sb111111111111111111111011111111111111111000000000000000000000000000000;
		9309: Delta = 69'sb000000000000000000001000000000000000001000000000000000000000000000000;
		21197: Delta = 69'sb111111111111111111111000000000000000001000000000000000000000000000000;
		29664: Delta = 69'sb000000000000000000000111111111111111111000000000000000000000000000000;
		41552: Delta = 69'sb111111111111111111110111111111111111111000000000000000000000000000000;
		3365: Delta = 69'sb000000000000000000010000000000000000001000000000000000000000000000000;
		27141: Delta = 69'sb111111111111111111110000000000000000001000000000000000000000000000000;
		23720: Delta = 69'sb000000000000000000001111111111111111111000000000000000000000000000000;
		47496: Delta = 69'sb111111111111111111101111111111111111111000000000000000000000000000000;
		42338: Delta = 69'sb000000000000000000100000000000000000001000000000000000000000000000000;
		39029: Delta = 69'sb111111111111111111100000000000000000001000000000000000000000000000000;
		11832: Delta = 69'sb000000000000000000011111111111111111111000000000000000000000000000000;
		8523: Delta = 69'sb111111111111111111011111111111111111111000000000000000000000000000000;
		18562: Delta = 69'sb000000000000000001000000000000000000001000000000000000000000000000000;
		11944: Delta = 69'sb111111111111111111000000000000000000001000000000000000000000000000000;
		38917: Delta = 69'sb000000000000000000111111111111111111111000000000000000000000000000000;
		32299: Delta = 69'sb111111111111111110111111111111111111111000000000000000000000000000000;
		21871: Delta = 69'sb000000000000000010000000000000000000001000000000000000000000000000000;
		8635: Delta = 69'sb111111111111111110000000000000000000001000000000000000000000000000000;
		42226: Delta = 69'sb000000000000000001111111111111111111111000000000000000000000000000000;
		28990: Delta = 69'sb111111111111111101111111111111111111111000000000000000000000000000000;
		28489: Delta = 69'sb000000000000000100000000000000000000001000000000000000000000000000000;
		2017: Delta = 69'sb111111111111111100000000000000000000001000000000000000000000000000000;
		48844: Delta = 69'sb000000000000000011111111111111111111111000000000000000000000000000000;
		22372: Delta = 69'sb111111111111111011111111111111111111111000000000000000000000000000000;
		41725: Delta = 69'sb000000000000001000000000000000000000001000000000000000000000000000000;
		39642: Delta = 69'sb111111111111111000000000000000000000001000000000000000000000000000000;
		11219: Delta = 69'sb000000000000000111111111111111111111111000000000000000000000000000000;
		9136: Delta = 69'sb111111111111110111111111111111111111111000000000000000000000000000000;
		17336: Delta = 69'sb000000000000010000000000000000000000001000000000000000000000000000000;
		13170: Delta = 69'sb111111111111110000000000000000000000001000000000000000000000000000000;
		37691: Delta = 69'sb000000000000001111111111111111111111111000000000000000000000000000000;
		33525: Delta = 69'sb111111111111101111111111111111111111111000000000000000000000000000000;
		19419: Delta = 69'sb000000000000100000000000000000000000001000000000000000000000000000000;
		11087: Delta = 69'sb111111111111100000000000000000000000001000000000000000000000000000000;
		39774: Delta = 69'sb000000000000011111111111111111111111111000000000000000000000000000000;
		31442: Delta = 69'sb111111111111011111111111111111111111111000000000000000000000000000000;
		23585: Delta = 69'sb000000000001000000000000000000000000001000000000000000000000000000000;
		6921: Delta = 69'sb111111111111000000000000000000000000001000000000000000000000000000000;
		43940: Delta = 69'sb000000000000111111111111111111111111111000000000000000000000000000000;
		27276: Delta = 69'sb111111111110111111111111111111111111111000000000000000000000000000000;
		31917: Delta = 69'sb000000000010000000000000000000000000001000000000000000000000000000000;
		49450: Delta = 69'sb111111111110000000000000000000000000001000000000000000000000000000000;
		1411: Delta = 69'sb000000000001111111111111111111111111111000000000000000000000000000000;
		18944: Delta = 69'sb111111111101111111111111111111111111111000000000000000000000000000000;
		48581: Delta = 69'sb000000000100000000000000000000000000001000000000000000000000000000000;
		32786: Delta = 69'sb111111111100000000000000000000000000001000000000000000000000000000000;
		18075: Delta = 69'sb000000000011111111111111111111111111111000000000000000000000000000000;
		2280: Delta = 69'sb111111111011111111111111111111111111111000000000000000000000000000000;
		31048: Delta = 69'sb000000001000000000000000000000000000001000000000000000000000000000000;
		50319: Delta = 69'sb111111111000000000000000000000000000001000000000000000000000000000000;
		542: Delta = 69'sb000000000111111111111111111111111111111000000000000000000000000000000;
		19813: Delta = 69'sb111111110111111111111111111111111111111000000000000000000000000000000;
		46843: Delta = 69'sb000000010000000000000000000000000000001000000000000000000000000000000;
		34524: Delta = 69'sb111111110000000000000000000000000000001000000000000000000000000000000;
		16337: Delta = 69'sb000000001111111111111111111111111111111000000000000000000000000000000;
		4018: Delta = 69'sb111111101111111111111111111111111111111000000000000000000000000000000;
		27572: Delta = 69'sb000000100000000000000000000000000000001000000000000000000000000000000;
		2934: Delta = 69'sb111111100000000000000000000000000000001000000000000000000000000000000;
		47927: Delta = 69'sb000000011111111111111111111111111111111000000000000000000000000000000;
		23289: Delta = 69'sb111111011111111111111111111111111111111000000000000000000000000000000;
		39891: Delta = 69'sb000001000000000000000000000000000000001000000000000000000000000000000;
		41476: Delta = 69'sb111111000000000000000000000000000000001000000000000000000000000000000;
		9385: Delta = 69'sb000000111111111111111111111111111111111000000000000000000000000000000;
		10970: Delta = 69'sb111110111111111111111111111111111111111000000000000000000000000000000;
		13668: Delta = 69'sb000010000000000000000000000000000000001000000000000000000000000000000;
		16838: Delta = 69'sb111110000000000000000000000000000000001000000000000000000000000000000;
		34023: Delta = 69'sb000001111111111111111111111111111111111000000000000000000000000000000;
		37193: Delta = 69'sb111101111111111111111111111111111111111000000000000000000000000000000;
		12083: Delta = 69'sb000100000000000000000000000000000000001000000000000000000000000000000;
		18423: Delta = 69'sb111100000000000000000000000000000000001000000000000000000000000000000;
		32438: Delta = 69'sb000011111111111111111111111111111111111000000000000000000000000000000;
		38778: Delta = 69'sb111011111111111111111111111111111111111000000000000000000000000000000;
		8913: Delta = 69'sb001000000000000000000000000000000000001000000000000000000000000000000;
		21593: Delta = 69'sb111000000000000000000000000000000000001000000000000000000000000000000;
		29268: Delta = 69'sb000111111111111111111111111111111111111000000000000000000000000000000;
		41948: Delta = 69'sb110111111111111111111111111111111111111000000000000000000000000000000;
		2573: Delta = 69'sb010000000000000000000000000000000000001000000000000000000000000000000;
		27933: Delta = 69'sb110000000000000000000000000000000000001000000000000000000000000000000;
		22928: Delta = 69'sb001111111111111111111111111111111111111000000000000000000000000000000;
		48288: Delta = 69'sb101111111111111111111111111111111111111000000000000000000000000000000;
		40657: Delta = 69'sb000000000000000000000000000000000000110000000000000000000000000000000;
		10204: Delta = 69'sb111111111111111111111111111111111111010000000000000000000000000000000;
		50808: Delta = 69'sb000000000000000000000000000000000001010000000000000000000000000000000;
		53: Delta = 69'sb111111111111111111111111111111111110110000000000000000000000000000000;
		20249: Delta = 69'sb000000000000000000000000000000000010010000000000000000000000000000000;
		40763: Delta = 69'sb111111111111111111111111111111111110010000000000000000000000000000000;
		10098: Delta = 69'sb000000000000000000000000000000000001110000000000000000000000000000000;
		30612: Delta = 69'sb111111111111111111111111111111111101110000000000000000000000000000000;
		9992: Delta = 69'sb000000000000000000000000000000000100010000000000000000000000000000000;
		159: Delta = 69'sb111111111111111111111111111111111100010000000000000000000000000000000;
		50702: Delta = 69'sb000000000000000000000000000000000011110000000000000000000000000000000;
		40869: Delta = 69'sb111111111111111111111111111111111011110000000000000000000000000000000;
		40339: Delta = 69'sb000000000000000000000000000000001000010000000000000000000000000000000;
		20673: Delta = 69'sb111111111111111111111111111111111000010000000000000000000000000000000;
		30188: Delta = 69'sb000000000000000000000000000000000111110000000000000000000000000000000;
		10522: Delta = 69'sb111111111111111111111111111111110111110000000000000000000000000000000;
		50172: Delta = 69'sb000000000000000000000000000000010000010000000000000000000000000000000;
		10840: Delta = 69'sb111111111111111111111111111111110000010000000000000000000000000000000;
		40021: Delta = 69'sb000000000000000000000000000000001111110000000000000000000000000000000;
		689: Delta = 69'sb111111111111111111111111111111101111110000000000000000000000000000000;
		18977: Delta = 69'sb000000000000000000000000000000100000010000000000000000000000000000000;
		42035: Delta = 69'sb111111111111111111111111111111100000010000000000000000000000000000000;
		8826: Delta = 69'sb000000000000000000000000000000011111110000000000000000000000000000000;
		31884: Delta = 69'sb111111111111111111111111111111011111110000000000000000000000000000000;
		7448: Delta = 69'sb000000000000000000000000000001000000010000000000000000000000000000000;
		2703: Delta = 69'sb111111111111111111111111111111000000010000000000000000000000000000000;
		48158: Delta = 69'sb000000000000000000000000000000111111110000000000000000000000000000000;
		43413: Delta = 69'sb111111111111111111111111111110111111110000000000000000000000000000000;
		35251: Delta = 69'sb000000000000000000000000000010000000010000000000000000000000000000000;
		25761: Delta = 69'sb111111111111111111111111111110000000010000000000000000000000000000000;
		25100: Delta = 69'sb000000000000000000000000000001111111110000000000000000000000000000000;
		15610: Delta = 69'sb111111111111111111111111111101111111110000000000000000000000000000000;
		39996: Delta = 69'sb000000000000000000000000000100000000010000000000000000000000000000000;
		21016: Delta = 69'sb111111111111111111111111111100000000010000000000000000000000000000000;
		29845: Delta = 69'sb000000000000000000000000000011111111110000000000000000000000000000000;
		10865: Delta = 69'sb111111111111111111111111111011111111110000000000000000000000000000000;
		49486: Delta = 69'sb000000000000000000000000001000000000010000000000000000000000000000000;
		11526: Delta = 69'sb111111111111111111111111111000000000010000000000000000000000000000000;
		39335: Delta = 69'sb000000000000000000000000000111111111110000000000000000000000000000000;
		1375: Delta = 69'sb111111111111111111111111110111111111110000000000000000000000000000000;
		17605: Delta = 69'sb000000000000000000000000010000000000010000000000000000000000000000000;
		43407: Delta = 69'sb111111111111111111111111110000000000010000000000000000000000000000000;
		7454: Delta = 69'sb000000000000000000000000001111111111110000000000000000000000000000000;
		33256: Delta = 69'sb111111111111111111111111101111111111110000000000000000000000000000000;
		4704: Delta = 69'sb000000000000000000000000100000000000010000000000000000000000000000000;
		5447: Delta = 69'sb111111111111111111111111100000000000010000000000000000000000000000000;
		45414: Delta = 69'sb000000000000000000000000011111111111110000000000000000000000000000000;
		46157: Delta = 69'sb111111111111111111111111011111111111110000000000000000000000000000000;
		29763: Delta = 69'sb000000000000000000000001000000000000010000000000000000000000000000000;
		31249: Delta = 69'sb111111111111111111111111000000000000010000000000000000000000000000000;
		19612: Delta = 69'sb000000000000000000000000111111111111110000000000000000000000000000000;
		21098: Delta = 69'sb111111111111111111111110111111111111110000000000000000000000000000000;
		29020: Delta = 69'sb000000000000000000000010000000000000010000000000000000000000000000000;
		31992: Delta = 69'sb111111111111111111111110000000000000010000000000000000000000000000000;
		18869: Delta = 69'sb000000000000000000000001111111111111110000000000000000000000000000000;
		21841: Delta = 69'sb111111111111111111111101111111111111110000000000000000000000000000000;
		27534: Delta = 69'sb000000000000000000000100000000000000010000000000000000000000000000000;
		33478: Delta = 69'sb111111111111111111111100000000000000010000000000000000000000000000000;
		17383: Delta = 69'sb000000000000000000000011111111111111110000000000000000000000000000000;
		23327: Delta = 69'sb111111111111111111111011111111111111110000000000000000000000000000000;
		24562: Delta = 69'sb000000000000000000001000000000000000010000000000000000000000000000000;
		36450: Delta = 69'sb111111111111111111111000000000000000010000000000000000000000000000000;
		14411: Delta = 69'sb000000000000000000000111111111111111110000000000000000000000000000000;
		26299: Delta = 69'sb111111111111111111110111111111111111110000000000000000000000000000000;
		18618: Delta = 69'sb000000000000000000010000000000000000010000000000000000000000000000000;
		42394: Delta = 69'sb111111111111111111110000000000000000010000000000000000000000000000000;
		8467: Delta = 69'sb000000000000000000001111111111111111110000000000000000000000000000000;
		32243: Delta = 69'sb111111111111111111101111111111111111110000000000000000000000000000000;
		6730: Delta = 69'sb000000000000000000100000000000000000010000000000000000000000000000000;
		3421: Delta = 69'sb111111111111111111100000000000000000010000000000000000000000000000000;
		47440: Delta = 69'sb000000000000000000011111111111111111110000000000000000000000000000000;
		44131: Delta = 69'sb111111111111111111011111111111111111110000000000000000000000000000000;
		33815: Delta = 69'sb000000000000000001000000000000000000010000000000000000000000000000000;
		27197: Delta = 69'sb111111111111111111000000000000000000010000000000000000000000000000000;
		23664: Delta = 69'sb000000000000000000111111111111111111110000000000000000000000000000000;
		17046: Delta = 69'sb111111111111111110111111111111111111110000000000000000000000000000000;
		37124: Delta = 69'sb000000000000000010000000000000000000010000000000000000000000000000000;
		23888: Delta = 69'sb111111111111111110000000000000000000010000000000000000000000000000000;
		26973: Delta = 69'sb000000000000000001111111111111111111110000000000000000000000000000000;
		13737: Delta = 69'sb111111111111111101111111111111111111110000000000000000000000000000000;
		43742: Delta = 69'sb000000000000000100000000000000000000010000000000000000000000000000000;
		17270: Delta = 69'sb111111111111111100000000000000000000010000000000000000000000000000000;
		33591: Delta = 69'sb000000000000000011111111111111111111110000000000000000000000000000000;
		7119: Delta = 69'sb111111111111111011111111111111111111110000000000000000000000000000000;
		6117: Delta = 69'sb000000000000001000000000000000000000010000000000000000000000000000000;
		4034: Delta = 69'sb111111111111111000000000000000000000010000000000000000000000000000000;
		46827: Delta = 69'sb000000000000000111111111111111111111110000000000000000000000000000000;
		44744: Delta = 69'sb111111111111110111111111111111111111110000000000000000000000000000000;
		32589: Delta = 69'sb000000000000010000000000000000000000010000000000000000000000000000000;
		28423: Delta = 69'sb111111111111110000000000000000000000010000000000000000000000000000000;
		22438: Delta = 69'sb000000000000001111111111111111111111110000000000000000000000000000000;
		18272: Delta = 69'sb111111111111101111111111111111111111110000000000000000000000000000000;
		34672: Delta = 69'sb000000000000100000000000000000000000010000000000000000000000000000000;
		26340: Delta = 69'sb111111111111100000000000000000000000010000000000000000000000000000000;
		24521: Delta = 69'sb000000000000011111111111111111111111110000000000000000000000000000000;
		16189: Delta = 69'sb111111111111011111111111111111111111110000000000000000000000000000000;
		38838: Delta = 69'sb000000000001000000000000000000000000010000000000000000000000000000000;
		22174: Delta = 69'sb111111111111000000000000000000000000010000000000000000000000000000000;
		28687: Delta = 69'sb000000000000111111111111111111111111110000000000000000000000000000000;
		12023: Delta = 69'sb111111111110111111111111111111111111110000000000000000000000000000000;
		47170: Delta = 69'sb000000000010000000000000000000000000010000000000000000000000000000000;
		13842: Delta = 69'sb111111111110000000000000000000000000010000000000000000000000000000000;
		37019: Delta = 69'sb000000000001111111111111111111111111110000000000000000000000000000000;
		3691: Delta = 69'sb111111111101111111111111111111111111110000000000000000000000000000000;
		12973: Delta = 69'sb000000000100000000000000000000000000010000000000000000000000000000000;
		48039: Delta = 69'sb111111111100000000000000000000000000010000000000000000000000000000000;
		2822: Delta = 69'sb000000000011111111111111111111111111110000000000000000000000000000000;
		37888: Delta = 69'sb111111111011111111111111111111111111110000000000000000000000000000000;
		46301: Delta = 69'sb000000001000000000000000000000000000010000000000000000000000000000000;
		14711: Delta = 69'sb111111111000000000000000000000000000010000000000000000000000000000000;
		36150: Delta = 69'sb000000000111111111111111111111111111110000000000000000000000000000000;
		4560: Delta = 69'sb111111110111111111111111111111111111110000000000000000000000000000000;
		11235: Delta = 69'sb000000010000000000000000000000000000010000000000000000000000000000000;
		49777: Delta = 69'sb111111110000000000000000000000000000010000000000000000000000000000000;
		1084: Delta = 69'sb000000001111111111111111111111111111110000000000000000000000000000000;
		39626: Delta = 69'sb111111101111111111111111111111111111110000000000000000000000000000000;
		42825: Delta = 69'sb000000100000000000000000000000000000010000000000000000000000000000000;
		18187: Delta = 69'sb111111100000000000000000000000000000010000000000000000000000000000000;
		32674: Delta = 69'sb000000011111111111111111111111111111110000000000000000000000000000000;
		8036: Delta = 69'sb111111011111111111111111111111111111110000000000000000000000000000000;
		4283: Delta = 69'sb000001000000000000000000000000000000010000000000000000000000000000000;
		5868: Delta = 69'sb111111000000000000000000000000000000010000000000000000000000000000000;
		44993: Delta = 69'sb000000111111111111111111111111111111110000000000000000000000000000000;
		46578: Delta = 69'sb111110111111111111111111111111111111110000000000000000000000000000000;
		28921: Delta = 69'sb000010000000000000000000000000000000010000000000000000000000000000000;
		32091: Delta = 69'sb111110000000000000000000000000000000010000000000000000000000000000000;
		18770: Delta = 69'sb000001111111111111111111111111111111110000000000000000000000000000000;
		21940: Delta = 69'sb111101111111111111111111111111111111110000000000000000000000000000000;
		27336: Delta = 69'sb000100000000000000000000000000000000010000000000000000000000000000000;
		33676: Delta = 69'sb111100000000000000000000000000000000010000000000000000000000000000000;
		17185: Delta = 69'sb000011111111111111111111111111111111110000000000000000000000000000000;
		23525: Delta = 69'sb111011111111111111111111111111111111110000000000000000000000000000000;
		24166: Delta = 69'sb001000000000000000000000000000000000010000000000000000000000000000000;
		36846: Delta = 69'sb111000000000000000000000000000000000010000000000000000000000000000000;
		14015: Delta = 69'sb000111111111111111111111111111111111110000000000000000000000000000000;
		26695: Delta = 69'sb110111111111111111111111111111111111110000000000000000000000000000000;
		17826: Delta = 69'sb010000000000000000000000000000000000010000000000000000000000000000000;
		43186: Delta = 69'sb110000000000000000000000000000000000010000000000000000000000000000000;
		7675: Delta = 69'sb001111111111111111111111111111111111110000000000000000000000000000000;
		33035: Delta = 69'sb101111111111111111111111111111111111110000000000000000000000000000000;
		30453: Delta = 69'sb000000000000000000000000000000000001100000000000000000000000000000000;
		20408: Delta = 69'sb111111111111111111111111111111111110100000000000000000000000000000000;
		50755: Delta = 69'sb000000000000000000000000000000000010100000000000000000000000000000000;
		106: Delta = 69'sb111111111111111111111111111111111101100000000000000000000000000000000;
		40498: Delta = 69'sb000000000000000000000000000000000100100000000000000000000000000000000;
		30665: Delta = 69'sb111111111111111111111111111111111100100000000000000000000000000000000;
		20196: Delta = 69'sb000000000000000000000000000000000011100000000000000000000000000000000;
		10363: Delta = 69'sb111111111111111111111111111111111011100000000000000000000000000000000;
		19984: Delta = 69'sb000000000000000000000000000000001000100000000000000000000000000000000;
		318: Delta = 69'sb111111111111111111111111111111111000100000000000000000000000000000000;
		50543: Delta = 69'sb000000000000000000000000000000000111100000000000000000000000000000000;
		30877: Delta = 69'sb111111111111111111111111111111110111100000000000000000000000000000000;
		29817: Delta = 69'sb000000000000000000000000000000010000100000000000000000000000000000000;
		41346: Delta = 69'sb111111111111111111111111111111110000100000000000000000000000000000000;
		9515: Delta = 69'sb000000000000000000000000000000001111100000000000000000000000000000000;
		21044: Delta = 69'sb111111111111111111111111111111101111100000000000000000000000000000000;
		49483: Delta = 69'sb000000000000000000000000000000100000100000000000000000000000000000000;
		21680: Delta = 69'sb111111111111111111111111111111100000100000000000000000000000000000000;
		29181: Delta = 69'sb000000000000000000000000000000011111100000000000000000000000000000000;
		1378: Delta = 69'sb111111111111111111111111111111011111100000000000000000000000000000000;
		37954: Delta = 69'sb000000000000000000000000000001000000100000000000000000000000000000000;
		33209: Delta = 69'sb111111111111111111111111111111000000100000000000000000000000000000000;
		17652: Delta = 69'sb000000000000000000000000000000111111100000000000000000000000000000000;
		12907: Delta = 69'sb111111111111111111111111111110111111100000000000000000000000000000000;
		14896: Delta = 69'sb000000000000000000000000000010000000100000000000000000000000000000000;
		5406: Delta = 69'sb111111111111111111111111111110000000100000000000000000000000000000000;
		45455: Delta = 69'sb000000000000000000000000000001111111100000000000000000000000000000000;
		35965: Delta = 69'sb111111111111111111111111111101111111100000000000000000000000000000000;
		19641: Delta = 69'sb000000000000000000000000000100000000100000000000000000000000000000000;
		661: Delta = 69'sb111111111111111111111111111100000000100000000000000000000000000000000;
		50200: Delta = 69'sb000000000000000000000000000011111111100000000000000000000000000000000;
		31220: Delta = 69'sb111111111111111111111111111011111111100000000000000000000000000000000;
		29131: Delta = 69'sb000000000000000000000000001000000000100000000000000000000000000000000;
		42032: Delta = 69'sb111111111111111111111111111000000000100000000000000000000000000000000;
		8829: Delta = 69'sb000000000000000000000000000111111111100000000000000000000000000000000;
		21730: Delta = 69'sb111111111111111111111111110111111111100000000000000000000000000000000;
		48111: Delta = 69'sb000000000000000000000000010000000000100000000000000000000000000000000;
		23052: Delta = 69'sb111111111111111111111111110000000000100000000000000000000000000000000;
		27809: Delta = 69'sb000000000000000000000000001111111111100000000000000000000000000000000;
		2750: Delta = 69'sb111111111111111111111111101111111111100000000000000000000000000000000;
		35210: Delta = 69'sb000000000000000000000000100000000000100000000000000000000000000000000;
		35953: Delta = 69'sb111111111111111111111111100000000000100000000000000000000000000000000;
		14908: Delta = 69'sb000000000000000000000000011111111111100000000000000000000000000000000;
		15651: Delta = 69'sb111111111111111111111111011111111111100000000000000000000000000000000;
		9408: Delta = 69'sb000000000000000000000001000000000000100000000000000000000000000000000;
		10894: Delta = 69'sb111111111111111111111111000000000000100000000000000000000000000000000;
		39967: Delta = 69'sb000000000000000000000000111111111111100000000000000000000000000000000;
		41453: Delta = 69'sb111111111111111111111110111111111111100000000000000000000000000000000;
		8665: Delta = 69'sb000000000000000000000010000000000000100000000000000000000000000000000;
		11637: Delta = 69'sb111111111111111111111110000000000000100000000000000000000000000000000;
		39224: Delta = 69'sb000000000000000000000001111111111111100000000000000000000000000000000;
		42196: Delta = 69'sb111111111111111111111101111111111111100000000000000000000000000000000;
		7179: Delta = 69'sb000000000000000000000100000000000000100000000000000000000000000000000;
		13123: Delta = 69'sb111111111111111111111100000000000000100000000000000000000000000000000;
		37738: Delta = 69'sb000000000000000000000011111111111111100000000000000000000000000000000;
		43682: Delta = 69'sb111111111111111111111011111111111111100000000000000000000000000000000;
		4207: Delta = 69'sb000000000000000000001000000000000000100000000000000000000000000000000;
		16095: Delta = 69'sb111111111111111111111000000000000000100000000000000000000000000000000;
		34766: Delta = 69'sb000000000000000000000111111111111111100000000000000000000000000000000;
		46654: Delta = 69'sb111111111111111111110111111111111111100000000000000000000000000000000;
		49124: Delta = 69'sb000000000000000000010000000000000000100000000000000000000000000000000;
		22039: Delta = 69'sb111111111111111111110000000000000000100000000000000000000000000000000;
		28822: Delta = 69'sb000000000000000000001111111111111111100000000000000000000000000000000;
		1737: Delta = 69'sb111111111111111111101111111111111111100000000000000000000000000000000;
		37236: Delta = 69'sb000000000000000000100000000000000000100000000000000000000000000000000;
		33927: Delta = 69'sb111111111111111111100000000000000000100000000000000000000000000000000;
		16934: Delta = 69'sb000000000000000000011111111111111111100000000000000000000000000000000;
		13625: Delta = 69'sb111111111111111111011111111111111111100000000000000000000000000000000;
		13460: Delta = 69'sb000000000000000001000000000000000000100000000000000000000000000000000;
		6842: Delta = 69'sb111111111111111111000000000000000000100000000000000000000000000000000;
		44019: Delta = 69'sb000000000000000000111111111111111111100000000000000000000000000000000;
		37401: Delta = 69'sb111111111111111110111111111111111111100000000000000000000000000000000;
		16769: Delta = 69'sb000000000000000010000000000000000000100000000000000000000000000000000;
		3533: Delta = 69'sb111111111111111110000000000000000000100000000000000000000000000000000;
		47328: Delta = 69'sb000000000000000001111111111111111111100000000000000000000000000000000;
		34092: Delta = 69'sb111111111111111101111111111111111111100000000000000000000000000000000;
		23387: Delta = 69'sb000000000000000100000000000000000000100000000000000000000000000000000;
		47776: Delta = 69'sb111111111111111100000000000000000000100000000000000000000000000000000;
		3085: Delta = 69'sb000000000000000011111111111111111111100000000000000000000000000000000;
		27474: Delta = 69'sb111111111111111011111111111111111111100000000000000000000000000000000;
		36623: Delta = 69'sb000000000000001000000000000000000000100000000000000000000000000000000;
		34540: Delta = 69'sb111111111111111000000000000000000000100000000000000000000000000000000;
		16321: Delta = 69'sb000000000000000111111111111111111111100000000000000000000000000000000;
		14238: Delta = 69'sb111111111111110111111111111111111111100000000000000000000000000000000;
		12234: Delta = 69'sb000000000000010000000000000000000000100000000000000000000000000000000;
		8068: Delta = 69'sb111111111111110000000000000000000000100000000000000000000000000000000;
		42793: Delta = 69'sb000000000000001111111111111111111111100000000000000000000000000000000;
		38627: Delta = 69'sb111111111111101111111111111111111111100000000000000000000000000000000;
		14317: Delta = 69'sb000000000000100000000000000000000000100000000000000000000000000000000;
		5985: Delta = 69'sb111111111111100000000000000000000000100000000000000000000000000000000;
		44876: Delta = 69'sb000000000000011111111111111111111111100000000000000000000000000000000;
		36544: Delta = 69'sb111111111111011111111111111111111111100000000000000000000000000000000;
		18483: Delta = 69'sb000000000001000000000000000000000000100000000000000000000000000000000;
		1819: Delta = 69'sb111111111111000000000000000000000000100000000000000000000000000000000;
		49042: Delta = 69'sb000000000000111111111111111111111111100000000000000000000000000000000;
		32378: Delta = 69'sb111111111110111111111111111111111111100000000000000000000000000000000;
		26815: Delta = 69'sb000000000010000000000000000000000000100000000000000000000000000000000;
		44348: Delta = 69'sb111111111110000000000000000000000000100000000000000000000000000000000;
		6513: Delta = 69'sb000000000001111111111111111111111111100000000000000000000000000000000;
		24046: Delta = 69'sb111111111101111111111111111111111111100000000000000000000000000000000;
		43479: Delta = 69'sb000000000100000000000000000000000000100000000000000000000000000000000;
		27684: Delta = 69'sb111111111100000000000000000000000000100000000000000000000000000000000;
		23177: Delta = 69'sb000000000011111111111111111111111111100000000000000000000000000000000;
		7382: Delta = 69'sb111111111011111111111111111111111111100000000000000000000000000000000;
		25946: Delta = 69'sb000000001000000000000000000000000000100000000000000000000000000000000;
		45217: Delta = 69'sb111111111000000000000000000000000000100000000000000000000000000000000;
		5644: Delta = 69'sb000000000111111111111111111111111111100000000000000000000000000000000;
		24915: Delta = 69'sb111111110111111111111111111111111111100000000000000000000000000000000;
		41741: Delta = 69'sb000000010000000000000000000000000000100000000000000000000000000000000;
		29422: Delta = 69'sb111111110000000000000000000000000000100000000000000000000000000000000;
		21439: Delta = 69'sb000000001111111111111111111111111111100000000000000000000000000000000;
		9120: Delta = 69'sb111111101111111111111111111111111111100000000000000000000000000000000;
		22470: Delta = 69'sb000000100000000000000000000000000000100000000000000000000000000000000;
		48693: Delta = 69'sb111111100000000000000000000000000000100000000000000000000000000000000;
		2168: Delta = 69'sb000000011111111111111111111111111111100000000000000000000000000000000;
		28391: Delta = 69'sb111111011111111111111111111111111111100000000000000000000000000000000;
		34789: Delta = 69'sb000001000000000000000000000000000000100000000000000000000000000000000;
		36374: Delta = 69'sb111111000000000000000000000000000000100000000000000000000000000000000;
		14487: Delta = 69'sb000000111111111111111111111111111111100000000000000000000000000000000;
		16072: Delta = 69'sb111110111111111111111111111111111111100000000000000000000000000000000;
		8566: Delta = 69'sb000010000000000000000000000000000000100000000000000000000000000000000;
		11736: Delta = 69'sb111110000000000000000000000000000000100000000000000000000000000000000;
		39125: Delta = 69'sb000001111111111111111111111111111111100000000000000000000000000000000;
		42295: Delta = 69'sb111101111111111111111111111111111111100000000000000000000000000000000;
		6981: Delta = 69'sb000100000000000000000000000000000000100000000000000000000000000000000;
		13321: Delta = 69'sb111100000000000000000000000000000000100000000000000000000000000000000;
		37540: Delta = 69'sb000011111111111111111111111111111111100000000000000000000000000000000;
		43880: Delta = 69'sb111011111111111111111111111111111111100000000000000000000000000000000;
		3811: Delta = 69'sb001000000000000000000000000000000000100000000000000000000000000000000;
		16491: Delta = 69'sb111000000000000000000000000000000000100000000000000000000000000000000;
		34370: Delta = 69'sb000111111111111111111111111111111111100000000000000000000000000000000;
		47050: Delta = 69'sb110111111111111111111111111111111111100000000000000000000000000000000;
		48332: Delta = 69'sb010000000000000000000000000000000000100000000000000000000000000000000;
		22831: Delta = 69'sb110000000000000000000000000000000000100000000000000000000000000000000;
		28030: Delta = 69'sb001111111111111111111111111111111111100000000000000000000000000000000;
		2529: Delta = 69'sb101111111111111111111111111111111111100000000000000000000000000000000;
		10045: Delta = 69'sb000000000000000000000000000000000011000000000000000000000000000000000;
		40816: Delta = 69'sb111111111111111111111111111111111101000000000000000000000000000000000;
		50649: Delta = 69'sb000000000000000000000000000000000101000000000000000000000000000000000;
		212: Delta = 69'sb111111111111111111111111111111111011000000000000000000000000000000000;
		30135: Delta = 69'sb000000000000000000000000000000001001000000000000000000000000000000000;
		10469: Delta = 69'sb111111111111111111111111111111111001000000000000000000000000000000000;
		40392: Delta = 69'sb000000000000000000000000000000000111000000000000000000000000000000000;
		20726: Delta = 69'sb111111111111111111111111111111110111000000000000000000000000000000000;
		39968: Delta = 69'sb000000000000000000000000000000010001000000000000000000000000000000000;
		636: Delta = 69'sb111111111111111111111111111111110001000000000000000000000000000000000;
		50225: Delta = 69'sb000000000000000000000000000000001111000000000000000000000000000000000;
		10893: Delta = 69'sb111111111111111111111111111111101111000000000000000000000000000000000;
		8773: Delta = 69'sb000000000000000000000000000000100001000000000000000000000000000000000;
		31831: Delta = 69'sb111111111111111111111111111111100001000000000000000000000000000000000;
		19030: Delta = 69'sb000000000000000000000000000000011111000000000000000000000000000000000;
		42088: Delta = 69'sb111111111111111111111111111111011111000000000000000000000000000000000;
		48105: Delta = 69'sb000000000000000000000000000001000001000000000000000000000000000000000;
		43360: Delta = 69'sb111111111111111111111111111111000001000000000000000000000000000000000;
		7501: Delta = 69'sb000000000000000000000000000000111111000000000000000000000000000000000;
		2756: Delta = 69'sb111111111111111111111111111110111111000000000000000000000000000000000;
		25047: Delta = 69'sb000000000000000000000000000010000001000000000000000000000000000000000;
		15557: Delta = 69'sb111111111111111111111111111110000001000000000000000000000000000000000;
		35304: Delta = 69'sb000000000000000000000000000001111111000000000000000000000000000000000;
		25814: Delta = 69'sb111111111111111111111111111101111111000000000000000000000000000000000;
		29792: Delta = 69'sb000000000000000000000000000100000001000000000000000000000000000000000;
		10812: Delta = 69'sb111111111111111111111111111100000001000000000000000000000000000000000;
		40049: Delta = 69'sb000000000000000000000000000011111111000000000000000000000000000000000;
		21069: Delta = 69'sb111111111111111111111111111011111111000000000000000000000000000000000;
		39282: Delta = 69'sb000000000000000000000000001000000001000000000000000000000000000000000;
		1322: Delta = 69'sb111111111111111111111111111000000001000000000000000000000000000000000;
		49539: Delta = 69'sb000000000000000000000000000111111111000000000000000000000000000000000;
		11579: Delta = 69'sb111111111111111111111111110111111111000000000000000000000000000000000;
		7401: Delta = 69'sb000000000000000000000000010000000001000000000000000000000000000000000;
		33203: Delta = 69'sb111111111111111111111111110000000001000000000000000000000000000000000;
		17658: Delta = 69'sb000000000000000000000000001111111111000000000000000000000000000000000;
		43460: Delta = 69'sb111111111111111111111111101111111111000000000000000000000000000000000;
		45361: Delta = 69'sb000000000000000000000000100000000001000000000000000000000000000000000;
		46104: Delta = 69'sb111111111111111111111111100000000001000000000000000000000000000000000;
		4757: Delta = 69'sb000000000000000000000000011111111111000000000000000000000000000000000;
		5500: Delta = 69'sb111111111111111111111111011111111111000000000000000000000000000000000;
		19559: Delta = 69'sb000000000000000000000001000000000001000000000000000000000000000000000;
		21045: Delta = 69'sb111111111111111111111111000000000001000000000000000000000000000000000;
		29816: Delta = 69'sb000000000000000000000000111111111111000000000000000000000000000000000;
		31302: Delta = 69'sb111111111111111111111110111111111111000000000000000000000000000000000;
		18816: Delta = 69'sb000000000000000000000010000000000001000000000000000000000000000000000;
		21788: Delta = 69'sb111111111111111111111110000000000001000000000000000000000000000000000;
		29073: Delta = 69'sb000000000000000000000001111111111111000000000000000000000000000000000;
		32045: Delta = 69'sb111111111111111111111101111111111111000000000000000000000000000000000;
		17330: Delta = 69'sb000000000000000000000100000000000001000000000000000000000000000000000;
		23274: Delta = 69'sb111111111111111111111100000000000001000000000000000000000000000000000;
		27587: Delta = 69'sb000000000000000000000011111111111111000000000000000000000000000000000;
		33531: Delta = 69'sb111111111111111111111011111111111111000000000000000000000000000000000;
		14358: Delta = 69'sb000000000000000000001000000000000001000000000000000000000000000000000;
		26246: Delta = 69'sb111111111111111111111000000000000001000000000000000000000000000000000;
		24615: Delta = 69'sb000000000000000000000111111111111111000000000000000000000000000000000;
		36503: Delta = 69'sb111111111111111111110111111111111111000000000000000000000000000000000;
		8414: Delta = 69'sb000000000000000000010000000000000001000000000000000000000000000000000;
		32190: Delta = 69'sb111111111111111111110000000000000001000000000000000000000000000000000;
		18671: Delta = 69'sb000000000000000000001111111111111111000000000000000000000000000000000;
		42447: Delta = 69'sb111111111111111111101111111111111111000000000000000000000000000000000;
		47387: Delta = 69'sb000000000000000000100000000000000001000000000000000000000000000000000;
		44078: Delta = 69'sb111111111111111111100000000000000001000000000000000000000000000000000;
		6783: Delta = 69'sb000000000000000000011111111111111111000000000000000000000000000000000;
		3474: Delta = 69'sb111111111111111111011111111111111111000000000000000000000000000000000;
		23611: Delta = 69'sb000000000000000001000000000000000001000000000000000000000000000000000;
		16993: Delta = 69'sb111111111111111111000000000000000001000000000000000000000000000000000;
		33868: Delta = 69'sb000000000000000000111111111111111111000000000000000000000000000000000;
		27250: Delta = 69'sb111111111111111110111111111111111111000000000000000000000000000000000;
		26920: Delta = 69'sb000000000000000010000000000000000001000000000000000000000000000000000;
		13684: Delta = 69'sb111111111111111110000000000000000001000000000000000000000000000000000;
		37177: Delta = 69'sb000000000000000001111111111111111111000000000000000000000000000000000;
		23941: Delta = 69'sb111111111111111101111111111111111111000000000000000000000000000000000;
		33538: Delta = 69'sb000000000000000100000000000000000001000000000000000000000000000000000;
		7066: Delta = 69'sb111111111111111100000000000000000001000000000000000000000000000000000;
		43795: Delta = 69'sb000000000000000011111111111111111111000000000000000000000000000000000;
		17323: Delta = 69'sb111111111111111011111111111111111111000000000000000000000000000000000;
		46774: Delta = 69'sb000000000000001000000000000000000001000000000000000000000000000000000;
		44691: Delta = 69'sb111111111111111000000000000000000001000000000000000000000000000000000;
		6170: Delta = 69'sb000000000000000111111111111111111111000000000000000000000000000000000;
		4087: Delta = 69'sb111111111111110111111111111111111111000000000000000000000000000000000;
		22385: Delta = 69'sb000000000000010000000000000000000001000000000000000000000000000000000;
		18219: Delta = 69'sb111111111111110000000000000000000001000000000000000000000000000000000;
		32642: Delta = 69'sb000000000000001111111111111111111111000000000000000000000000000000000;
		28476: Delta = 69'sb111111111111101111111111111111111111000000000000000000000000000000000;
		24468: Delta = 69'sb000000000000100000000000000000000001000000000000000000000000000000000;
		16136: Delta = 69'sb111111111111100000000000000000000001000000000000000000000000000000000;
		34725: Delta = 69'sb000000000000011111111111111111111111000000000000000000000000000000000;
		26393: Delta = 69'sb111111111111011111111111111111111111000000000000000000000000000000000;
		28634: Delta = 69'sb000000000001000000000000000000000001000000000000000000000000000000000;
		11970: Delta = 69'sb111111111111000000000000000000000001000000000000000000000000000000000;
		38891: Delta = 69'sb000000000000111111111111111111111111000000000000000000000000000000000;
		22227: Delta = 69'sb111111111110111111111111111111111111000000000000000000000000000000000;
		36966: Delta = 69'sb000000000010000000000000000000000001000000000000000000000000000000000;
		3638: Delta = 69'sb111111111110000000000000000000000001000000000000000000000000000000000;
		47223: Delta = 69'sb000000000001111111111111111111111111000000000000000000000000000000000;
		13895: Delta = 69'sb111111111101111111111111111111111111000000000000000000000000000000000;
		2769: Delta = 69'sb000000000100000000000000000000000001000000000000000000000000000000000;
		37835: Delta = 69'sb111111111100000000000000000000000001000000000000000000000000000000000;
		13026: Delta = 69'sb000000000011111111111111111111111111000000000000000000000000000000000;
		48092: Delta = 69'sb111111111011111111111111111111111111000000000000000000000000000000000;
		36097: Delta = 69'sb000000001000000000000000000000000001000000000000000000000000000000000;
		4507: Delta = 69'sb111111111000000000000000000000000001000000000000000000000000000000000;
		46354: Delta = 69'sb000000000111111111111111111111111111000000000000000000000000000000000;
		14764: Delta = 69'sb111111110111111111111111111111111111000000000000000000000000000000000;
		1031: Delta = 69'sb000000010000000000000000000000000001000000000000000000000000000000000;
		39573: Delta = 69'sb111111110000000000000000000000000001000000000000000000000000000000000;
		11288: Delta = 69'sb000000001111111111111111111111111111000000000000000000000000000000000;
		49830: Delta = 69'sb111111101111111111111111111111111111000000000000000000000000000000000;
		32621: Delta = 69'sb000000100000000000000000000000000001000000000000000000000000000000000;
		7983: Delta = 69'sb111111100000000000000000000000000001000000000000000000000000000000000;
		42878: Delta = 69'sb000000011111111111111111111111111111000000000000000000000000000000000;
		18240: Delta = 69'sb111111011111111111111111111111111111000000000000000000000000000000000;
		44940: Delta = 69'sb000001000000000000000000000000000001000000000000000000000000000000000;
		46525: Delta = 69'sb111111000000000000000000000000000001000000000000000000000000000000000;
		4336: Delta = 69'sb000000111111111111111111111111111111000000000000000000000000000000000;
		5921: Delta = 69'sb111110111111111111111111111111111111000000000000000000000000000000000;
		18717: Delta = 69'sb000010000000000000000000000000000001000000000000000000000000000000000;
		21887: Delta = 69'sb111110000000000000000000000000000001000000000000000000000000000000000;
		28974: Delta = 69'sb000001111111111111111111111111111111000000000000000000000000000000000;
		32144: Delta = 69'sb111101111111111111111111111111111111000000000000000000000000000000000;
		17132: Delta = 69'sb000100000000000000000000000000000001000000000000000000000000000000000;
		23472: Delta = 69'sb111100000000000000000000000000000001000000000000000000000000000000000;
		27389: Delta = 69'sb000011111111111111111111111111111111000000000000000000000000000000000;
		33729: Delta = 69'sb111011111111111111111111111111111111000000000000000000000000000000000;
		13962: Delta = 69'sb001000000000000000000000000000000001000000000000000000000000000000000;
		26642: Delta = 69'sb111000000000000000000000000000000001000000000000000000000000000000000;
		24219: Delta = 69'sb000111111111111111111111111111111111000000000000000000000000000000000;
		36899: Delta = 69'sb110111111111111111111111111111111111000000000000000000000000000000000;
		7622: Delta = 69'sb010000000000000000000000000000000001000000000000000000000000000000000;
		32982: Delta = 69'sb110000000000000000000000000000000001000000000000000000000000000000000;
		17879: Delta = 69'sb001111111111111111111111111111111111000000000000000000000000000000000;
		43239: Delta = 69'sb101111111111111111111111111111111111000000000000000000000000000000000;
		20090: Delta = 69'sb000000000000000000000000000000000110000000000000000000000000000000000;
		30771: Delta = 69'sb111111111111111111111111111111111010000000000000000000000000000000000;
		50437: Delta = 69'sb000000000000000000000000000000001010000000000000000000000000000000000;
		424: Delta = 69'sb111111111111111111111111111111110110000000000000000000000000000000000;
		9409: Delta = 69'sb000000000000000000000000000000010010000000000000000000000000000000000;
		20938: Delta = 69'sb111111111111111111111111111111110010000000000000000000000000000000000;
		29923: Delta = 69'sb000000000000000000000000000000001110000000000000000000000000000000000;
		41452: Delta = 69'sb111111111111111111111111111111101110000000000000000000000000000000000;
		29075: Delta = 69'sb000000000000000000000000000000100010000000000000000000000000000000000;
		1272: Delta = 69'sb111111111111111111111111111111100010000000000000000000000000000000000;
		49589: Delta = 69'sb000000000000000000000000000000011110000000000000000000000000000000000;
		21786: Delta = 69'sb111111111111111111111111111111011110000000000000000000000000000000000;
		17546: Delta = 69'sb000000000000000000000000000001000010000000000000000000000000000000000;
		12801: Delta = 69'sb111111111111111111111111111111000010000000000000000000000000000000000;
		38060: Delta = 69'sb000000000000000000000000000000111110000000000000000000000000000000000;
		33315: Delta = 69'sb111111111111111111111111111110111110000000000000000000000000000000000;
		45349: Delta = 69'sb000000000000000000000000000010000010000000000000000000000000000000000;
		35859: Delta = 69'sb111111111111111111111111111110000010000000000000000000000000000000000;
		15002: Delta = 69'sb000000000000000000000000000001111110000000000000000000000000000000000;
		5512: Delta = 69'sb111111111111111111111111111101111110000000000000000000000000000000000;
		50094: Delta = 69'sb000000000000000000000000000100000010000000000000000000000000000000000;
		31114: Delta = 69'sb111111111111111111111111111100000010000000000000000000000000000000000;
		19747: Delta = 69'sb000000000000000000000000000011111110000000000000000000000000000000000;
		767: Delta = 69'sb111111111111111111111111111011111110000000000000000000000000000000000;
		8723: Delta = 69'sb000000000000000000000000001000000010000000000000000000000000000000000;
		21624: Delta = 69'sb111111111111111111111111111000000010000000000000000000000000000000000;
		29237: Delta = 69'sb000000000000000000000000000111111110000000000000000000000000000000000;
		42138: Delta = 69'sb111111111111111111111111110111111110000000000000000000000000000000000;
		27703: Delta = 69'sb000000000000000000000000010000000010000000000000000000000000000000000;
		2644: Delta = 69'sb111111111111111111111111110000000010000000000000000000000000000000000;
		48217: Delta = 69'sb000000000000000000000000001111111110000000000000000000000000000000000;
		23158: Delta = 69'sb111111111111111111111111101111111110000000000000000000000000000000000;
		14802: Delta = 69'sb000000000000000000000000100000000010000000000000000000000000000000000;
		15545: Delta = 69'sb111111111111111111111111100000000010000000000000000000000000000000000;
		35316: Delta = 69'sb000000000000000000000000011111111110000000000000000000000000000000000;
		36059: Delta = 69'sb111111111111111111111111011111111110000000000000000000000000000000000;
		39861: Delta = 69'sb000000000000000000000001000000000010000000000000000000000000000000000;
		41347: Delta = 69'sb111111111111111111111111000000000010000000000000000000000000000000000;
		9514: Delta = 69'sb000000000000000000000000111111111110000000000000000000000000000000000;
		11000: Delta = 69'sb111111111111111111111110111111111110000000000000000000000000000000000;
		39118: Delta = 69'sb000000000000000000000010000000000010000000000000000000000000000000000;
		42090: Delta = 69'sb111111111111111111111110000000000010000000000000000000000000000000000;
		8771: Delta = 69'sb000000000000000000000001111111111110000000000000000000000000000000000;
		11743: Delta = 69'sb111111111111111111111101111111111110000000000000000000000000000000000;
		37632: Delta = 69'sb000000000000000000000100000000000010000000000000000000000000000000000;
		43576: Delta = 69'sb111111111111111111111100000000000010000000000000000000000000000000000;
		7285: Delta = 69'sb000000000000000000000011111111111110000000000000000000000000000000000;
		13229: Delta = 69'sb111111111111111111111011111111111110000000000000000000000000000000000;
		34660: Delta = 69'sb000000000000000000001000000000000010000000000000000000000000000000000;
		46548: Delta = 69'sb111111111111111111111000000000000010000000000000000000000000000000000;
		4313: Delta = 69'sb000000000000000000000111111111111110000000000000000000000000000000000;
		16201: Delta = 69'sb111111111111111111110111111111111110000000000000000000000000000000000;
		28716: Delta = 69'sb000000000000000000010000000000000010000000000000000000000000000000000;
		1631: Delta = 69'sb111111111111111111110000000000000010000000000000000000000000000000000;
		49230: Delta = 69'sb000000000000000000001111111111111110000000000000000000000000000000000;
		22145: Delta = 69'sb111111111111111111101111111111111110000000000000000000000000000000000;
		16828: Delta = 69'sb000000000000000000100000000000000010000000000000000000000000000000000;
		13519: Delta = 69'sb111111111111111111100000000000000010000000000000000000000000000000000;
		37342: Delta = 69'sb000000000000000000011111111111111110000000000000000000000000000000000;
		34033: Delta = 69'sb111111111111111111011111111111111110000000000000000000000000000000000;
		43913: Delta = 69'sb000000000000000001000000000000000010000000000000000000000000000000000;
		37295: Delta = 69'sb111111111111111111000000000000000010000000000000000000000000000000000;
		13566: Delta = 69'sb000000000000000000111111111111111110000000000000000000000000000000000;
		6948: Delta = 69'sb111111111111111110111111111111111110000000000000000000000000000000000;
		47222: Delta = 69'sb000000000000000010000000000000000010000000000000000000000000000000000;
		33986: Delta = 69'sb111111111111111110000000000000000010000000000000000000000000000000000;
		16875: Delta = 69'sb000000000000000001111111111111111110000000000000000000000000000000000;
		3639: Delta = 69'sb111111111111111101111111111111111110000000000000000000000000000000000;
		2979: Delta = 69'sb000000000000000100000000000000000010000000000000000000000000000000000;
		27368: Delta = 69'sb111111111111111100000000000000000010000000000000000000000000000000000;
		23493: Delta = 69'sb000000000000000011111111111111111110000000000000000000000000000000000;
		47882: Delta = 69'sb111111111111111011111111111111111110000000000000000000000000000000000;
		16215: Delta = 69'sb000000000000001000000000000000000010000000000000000000000000000000000;
		14132: Delta = 69'sb111111111111111000000000000000000010000000000000000000000000000000000;
		36729: Delta = 69'sb000000000000000111111111111111111110000000000000000000000000000000000;
		34646: Delta = 69'sb111111111111110111111111111111111110000000000000000000000000000000000;
		42687: Delta = 69'sb000000000000010000000000000000000010000000000000000000000000000000000;
		38521: Delta = 69'sb111111111111110000000000000000000010000000000000000000000000000000000;
		12340: Delta = 69'sb000000000000001111111111111111111110000000000000000000000000000000000;
		8174: Delta = 69'sb111111111111101111111111111111111110000000000000000000000000000000000;
		44770: Delta = 69'sb000000000000100000000000000000000010000000000000000000000000000000000;
		36438: Delta = 69'sb111111111111100000000000000000000010000000000000000000000000000000000;
		14423: Delta = 69'sb000000000000011111111111111111111110000000000000000000000000000000000;
		6091: Delta = 69'sb111111111111011111111111111111111110000000000000000000000000000000000;
		48936: Delta = 69'sb000000000001000000000000000000000010000000000000000000000000000000000;
		32272: Delta = 69'sb111111111111000000000000000000000010000000000000000000000000000000000;
		18589: Delta = 69'sb000000000000111111111111111111111110000000000000000000000000000000000;
		1925: Delta = 69'sb111111111110111111111111111111111110000000000000000000000000000000000;
		6407: Delta = 69'sb000000000010000000000000000000000010000000000000000000000000000000000;
		23940: Delta = 69'sb111111111110000000000000000000000010000000000000000000000000000000000;
		26921: Delta = 69'sb000000000001111111111111111111111110000000000000000000000000000000000;
		44454: Delta = 69'sb111111111101111111111111111111111110000000000000000000000000000000000;
		23071: Delta = 69'sb000000000100000000000000000000000010000000000000000000000000000000000;
		7276: Delta = 69'sb111111111100000000000000000000000010000000000000000000000000000000000;
		43585: Delta = 69'sb000000000011111111111111111111111110000000000000000000000000000000000;
		27790: Delta = 69'sb111111111011111111111111111111111110000000000000000000000000000000000;
		5538: Delta = 69'sb000000001000000000000000000000000010000000000000000000000000000000000;
		24809: Delta = 69'sb111111111000000000000000000000000010000000000000000000000000000000000;
		26052: Delta = 69'sb000000000111111111111111111111111110000000000000000000000000000000000;
		45323: Delta = 69'sb111111110111111111111111111111111110000000000000000000000000000000000;
		21333: Delta = 69'sb000000010000000000000000000000000010000000000000000000000000000000000;
		9014: Delta = 69'sb111111110000000000000000000000000010000000000000000000000000000000000;
		41847: Delta = 69'sb000000001111111111111111111111111110000000000000000000000000000000000;
		29528: Delta = 69'sb111111101111111111111111111111111110000000000000000000000000000000000;
		2062: Delta = 69'sb000000100000000000000000000000000010000000000000000000000000000000000;
		28285: Delta = 69'sb111111100000000000000000000000000010000000000000000000000000000000000;
		22576: Delta = 69'sb000000011111111111111111111111111110000000000000000000000000000000000;
		48799: Delta = 69'sb111111011111111111111111111111111110000000000000000000000000000000000;
		14381: Delta = 69'sb000001000000000000000000000000000010000000000000000000000000000000000;
		15966: Delta = 69'sb111111000000000000000000000000000010000000000000000000000000000000000;
		34895: Delta = 69'sb000000111111111111111111111111111110000000000000000000000000000000000;
		36480: Delta = 69'sb111110111111111111111111111111111110000000000000000000000000000000000;
		39019: Delta = 69'sb000010000000000000000000000000000010000000000000000000000000000000000;
		42189: Delta = 69'sb111110000000000000000000000000000010000000000000000000000000000000000;
		8672: Delta = 69'sb000001111111111111111111111111111110000000000000000000000000000000000;
		11842: Delta = 69'sb111101111111111111111111111111111110000000000000000000000000000000000;
		37434: Delta = 69'sb000100000000000000000000000000000010000000000000000000000000000000000;
		43774: Delta = 69'sb111100000000000000000000000000000010000000000000000000000000000000000;
		7087: Delta = 69'sb000011111111111111111111111111111110000000000000000000000000000000000;
		13427: Delta = 69'sb111011111111111111111111111111111110000000000000000000000000000000000;
		34264: Delta = 69'sb001000000000000000000000000000000010000000000000000000000000000000000;
		46944: Delta = 69'sb111000000000000000000000000000000010000000000000000000000000000000000;
		3917: Delta = 69'sb000111111111111111111111111111111110000000000000000000000000000000000;
		16597: Delta = 69'sb110111111111111111111111111111111110000000000000000000000000000000000;
		27924: Delta = 69'sb010000000000000000000000000000000010000000000000000000000000000000000;
		2423: Delta = 69'sb110000000000000000000000000000000010000000000000000000000000000000000;
		48438: Delta = 69'sb001111111111111111111111111111111110000000000000000000000000000000000;
		22937: Delta = 69'sb101111111111111111111111111111111110000000000000000000000000000000000;
		40180: Delta = 69'sb000000000000000000000000000000001100000000000000000000000000000000000;
		10681: Delta = 69'sb111111111111111111111111111111110100000000000000000000000000000000000;
		50013: Delta = 69'sb000000000000000000000000000000010100000000000000000000000000000000000;
		848: Delta = 69'sb111111111111111111111111111111101100000000000000000000000000000000000;
		18818: Delta = 69'sb000000000000000000000000000000100100000000000000000000000000000000000;
		41876: Delta = 69'sb111111111111111111111111111111100100000000000000000000000000000000000;
		8985: Delta = 69'sb000000000000000000000000000000011100000000000000000000000000000000000;
		32043: Delta = 69'sb111111111111111111111111111111011100000000000000000000000000000000000;
		7289: Delta = 69'sb000000000000000000000000000001000100000000000000000000000000000000000;
		2544: Delta = 69'sb111111111111111111111111111111000100000000000000000000000000000000000;
		48317: Delta = 69'sb000000000000000000000000000000111100000000000000000000000000000000000;
		43572: Delta = 69'sb111111111111111111111111111110111100000000000000000000000000000000000;
		35092: Delta = 69'sb000000000000000000000000000010000100000000000000000000000000000000000;
		25602: Delta = 69'sb111111111111111111111111111110000100000000000000000000000000000000000;
		25259: Delta = 69'sb000000000000000000000000000001111100000000000000000000000000000000000;
		15769: Delta = 69'sb111111111111111111111111111101111100000000000000000000000000000000000;
		39837: Delta = 69'sb000000000000000000000000000100000100000000000000000000000000000000000;
		20857: Delta = 69'sb111111111111111111111111111100000100000000000000000000000000000000000;
		30004: Delta = 69'sb000000000000000000000000000011111100000000000000000000000000000000000;
		11024: Delta = 69'sb111111111111111111111111111011111100000000000000000000000000000000000;
		49327: Delta = 69'sb000000000000000000000000001000000100000000000000000000000000000000000;
		11367: Delta = 69'sb111111111111111111111111111000000100000000000000000000000000000000000;
		39494: Delta = 69'sb000000000000000000000000000111111100000000000000000000000000000000000;
		1534: Delta = 69'sb111111111111111111111111110111111100000000000000000000000000000000000;
		17446: Delta = 69'sb000000000000000000000000010000000100000000000000000000000000000000000;
		43248: Delta = 69'sb111111111111111111111111110000000100000000000000000000000000000000000;
		7613: Delta = 69'sb000000000000000000000000001111111100000000000000000000000000000000000;
		33415: Delta = 69'sb111111111111111111111111101111111100000000000000000000000000000000000;
		4545: Delta = 69'sb000000000000000000000000100000000100000000000000000000000000000000000;
		5288: Delta = 69'sb111111111111111111111111100000000100000000000000000000000000000000000;
		45573: Delta = 69'sb000000000000000000000000011111111100000000000000000000000000000000000;
		46316: Delta = 69'sb111111111111111111111111011111111100000000000000000000000000000000000;
		29604: Delta = 69'sb000000000000000000000001000000000100000000000000000000000000000000000;
		31090: Delta = 69'sb111111111111111111111111000000000100000000000000000000000000000000000;
		19771: Delta = 69'sb000000000000000000000000111111111100000000000000000000000000000000000;
		21257: Delta = 69'sb111111111111111111111110111111111100000000000000000000000000000000000;
		28861: Delta = 69'sb000000000000000000000010000000000100000000000000000000000000000000000;
		31833: Delta = 69'sb111111111111111111111110000000000100000000000000000000000000000000000;
		19028: Delta = 69'sb000000000000000000000001111111111100000000000000000000000000000000000;
		22000: Delta = 69'sb111111111111111111111101111111111100000000000000000000000000000000000;
		27375: Delta = 69'sb000000000000000000000100000000000100000000000000000000000000000000000;
		33319: Delta = 69'sb111111111111111111111100000000000100000000000000000000000000000000000;
		17542: Delta = 69'sb000000000000000000000011111111111100000000000000000000000000000000000;
		23486: Delta = 69'sb111111111111111111111011111111111100000000000000000000000000000000000;
		24403: Delta = 69'sb000000000000000000001000000000000100000000000000000000000000000000000;
		36291: Delta = 69'sb111111111111111111111000000000000100000000000000000000000000000000000;
		14570: Delta = 69'sb000000000000000000000111111111111100000000000000000000000000000000000;
		26458: Delta = 69'sb111111111111111111110111111111111100000000000000000000000000000000000;
		18459: Delta = 69'sb000000000000000000010000000000000100000000000000000000000000000000000;
		42235: Delta = 69'sb111111111111111111110000000000000100000000000000000000000000000000000;
		8626: Delta = 69'sb000000000000000000001111111111111100000000000000000000000000000000000;
		32402: Delta = 69'sb111111111111111111101111111111111100000000000000000000000000000000000;
		6571: Delta = 69'sb000000000000000000100000000000000100000000000000000000000000000000000;
		3262: Delta = 69'sb111111111111111111100000000000000100000000000000000000000000000000000;
		47599: Delta = 69'sb000000000000000000011111111111111100000000000000000000000000000000000;
		44290: Delta = 69'sb111111111111111111011111111111111100000000000000000000000000000000000;
		33656: Delta = 69'sb000000000000000001000000000000000100000000000000000000000000000000000;
		27038: Delta = 69'sb111111111111111111000000000000000100000000000000000000000000000000000;
		23823: Delta = 69'sb000000000000000000111111111111111100000000000000000000000000000000000;
		17205: Delta = 69'sb111111111111111110111111111111111100000000000000000000000000000000000;
		36965: Delta = 69'sb000000000000000010000000000000000100000000000000000000000000000000000;
		23729: Delta = 69'sb111111111111111110000000000000000100000000000000000000000000000000000;
		27132: Delta = 69'sb000000000000000001111111111111111100000000000000000000000000000000000;
		13896: Delta = 69'sb111111111111111101111111111111111100000000000000000000000000000000000;
		43583: Delta = 69'sb000000000000000100000000000000000100000000000000000000000000000000000;
		17111: Delta = 69'sb111111111111111100000000000000000100000000000000000000000000000000000;
		33750: Delta = 69'sb000000000000000011111111111111111100000000000000000000000000000000000;
		7278: Delta = 69'sb111111111111111011111111111111111100000000000000000000000000000000000;
		5958: Delta = 69'sb000000000000001000000000000000000100000000000000000000000000000000000;
		3875: Delta = 69'sb111111111111111000000000000000000100000000000000000000000000000000000;
		46986: Delta = 69'sb000000000000000111111111111111111100000000000000000000000000000000000;
		44903: Delta = 69'sb111111111111110111111111111111111100000000000000000000000000000000000;
		32430: Delta = 69'sb000000000000010000000000000000000100000000000000000000000000000000000;
		28264: Delta = 69'sb111111111111110000000000000000000100000000000000000000000000000000000;
		22597: Delta = 69'sb000000000000001111111111111111111100000000000000000000000000000000000;
		18431: Delta = 69'sb111111111111101111111111111111111100000000000000000000000000000000000;
		34513: Delta = 69'sb000000000000100000000000000000000100000000000000000000000000000000000;
		26181: Delta = 69'sb111111111111100000000000000000000100000000000000000000000000000000000;
		24680: Delta = 69'sb000000000000011111111111111111111100000000000000000000000000000000000;
		16348: Delta = 69'sb111111111111011111111111111111111100000000000000000000000000000000000;
		38679: Delta = 69'sb000000000001000000000000000000000100000000000000000000000000000000000;
		22015: Delta = 69'sb111111111111000000000000000000000100000000000000000000000000000000000;
		28846: Delta = 69'sb000000000000111111111111111111111100000000000000000000000000000000000;
		12182: Delta = 69'sb111111111110111111111111111111111100000000000000000000000000000000000;
		47011: Delta = 69'sb000000000010000000000000000000000100000000000000000000000000000000000;
		13683: Delta = 69'sb111111111110000000000000000000000100000000000000000000000000000000000;
		37178: Delta = 69'sb000000000001111111111111111111111100000000000000000000000000000000000;
		3850: Delta = 69'sb111111111101111111111111111111111100000000000000000000000000000000000;
		12814: Delta = 69'sb000000000100000000000000000000000100000000000000000000000000000000000;
		47880: Delta = 69'sb111111111100000000000000000000000100000000000000000000000000000000000;
		2981: Delta = 69'sb000000000011111111111111111111111100000000000000000000000000000000000;
		38047: Delta = 69'sb111111111011111111111111111111111100000000000000000000000000000000000;
		46142: Delta = 69'sb000000001000000000000000000000000100000000000000000000000000000000000;
		14552: Delta = 69'sb111111111000000000000000000000000100000000000000000000000000000000000;
		36309: Delta = 69'sb000000000111111111111111111111111100000000000000000000000000000000000;
		4719: Delta = 69'sb111111110111111111111111111111111100000000000000000000000000000000000;
		11076: Delta = 69'sb000000010000000000000000000000000100000000000000000000000000000000000;
		49618: Delta = 69'sb111111110000000000000000000000000100000000000000000000000000000000000;
		1243: Delta = 69'sb000000001111111111111111111111111100000000000000000000000000000000000;
		39785: Delta = 69'sb111111101111111111111111111111111100000000000000000000000000000000000;
		42666: Delta = 69'sb000000100000000000000000000000000100000000000000000000000000000000000;
		18028: Delta = 69'sb111111100000000000000000000000000100000000000000000000000000000000000;
		32833: Delta = 69'sb000000011111111111111111111111111100000000000000000000000000000000000;
		8195: Delta = 69'sb111111011111111111111111111111111100000000000000000000000000000000000;
		4124: Delta = 69'sb000001000000000000000000000000000100000000000000000000000000000000000;
		5709: Delta = 69'sb111111000000000000000000000000000100000000000000000000000000000000000;
		45152: Delta = 69'sb000000111111111111111111111111111100000000000000000000000000000000000;
		46737: Delta = 69'sb111110111111111111111111111111111100000000000000000000000000000000000;
		28762: Delta = 69'sb000010000000000000000000000000000100000000000000000000000000000000000;
		31932: Delta = 69'sb111110000000000000000000000000000100000000000000000000000000000000000;
		18929: Delta = 69'sb000001111111111111111111111111111100000000000000000000000000000000000;
		22099: Delta = 69'sb111101111111111111111111111111111100000000000000000000000000000000000;
		27177: Delta = 69'sb000100000000000000000000000000000100000000000000000000000000000000000;
		33517: Delta = 69'sb111100000000000000000000000000000100000000000000000000000000000000000;
		17344: Delta = 69'sb000011111111111111111111111111111100000000000000000000000000000000000;
		23684: Delta = 69'sb111011111111111111111111111111111100000000000000000000000000000000000;
		24007: Delta = 69'sb001000000000000000000000000000000100000000000000000000000000000000000;
		36687: Delta = 69'sb111000000000000000000000000000000100000000000000000000000000000000000;
		14174: Delta = 69'sb000111111111111111111111111111111100000000000000000000000000000000000;
		26854: Delta = 69'sb110111111111111111111111111111111100000000000000000000000000000000000;
		17667: Delta = 69'sb010000000000000000000000000000000100000000000000000000000000000000000;
		43027: Delta = 69'sb110000000000000000000000000000000100000000000000000000000000000000000;
		7834: Delta = 69'sb001111111111111111111111111111111100000000000000000000000000000000000;
		33194: Delta = 69'sb101111111111111111111111111111111100000000000000000000000000000000000;
		29499: Delta = 69'sb000000000000000000000000000000011000000000000000000000000000000000000;
		21362: Delta = 69'sb111111111111111111111111111111101000000000000000000000000000000000000;
		49165: Delta = 69'sb000000000000000000000000000000101000000000000000000000000000000000000;
		1696: Delta = 69'sb111111111111111111111111111111011000000000000000000000000000000000000;
		37636: Delta = 69'sb000000000000000000000000000001001000000000000000000000000000000000000;
		32891: Delta = 69'sb111111111111111111111111111111001000000000000000000000000000000000000;
		17970: Delta = 69'sb000000000000000000000000000000111000000000000000000000000000000000000;
		13225: Delta = 69'sb111111111111111111111111111110111000000000000000000000000000000000000;
		14578: Delta = 69'sb000000000000000000000000000010001000000000000000000000000000000000000;
		5088: Delta = 69'sb111111111111111111111111111110001000000000000000000000000000000000000;
		45773: Delta = 69'sb000000000000000000000000000001111000000000000000000000000000000000000;
		36283: Delta = 69'sb111111111111111111111111111101111000000000000000000000000000000000000;
		19323: Delta = 69'sb000000000000000000000000000100001000000000000000000000000000000000000;
		343: Delta = 69'sb111111111111111111111111111100001000000000000000000000000000000000000;
		50518: Delta = 69'sb000000000000000000000000000011111000000000000000000000000000000000000;
		31538: Delta = 69'sb111111111111111111111111111011111000000000000000000000000000000000000;
		28813: Delta = 69'sb000000000000000000000000001000001000000000000000000000000000000000000;
		41714: Delta = 69'sb111111111111111111111111111000001000000000000000000000000000000000000;
		9147: Delta = 69'sb000000000000000000000000000111111000000000000000000000000000000000000;
		22048: Delta = 69'sb111111111111111111111111110111111000000000000000000000000000000000000;
		47793: Delta = 69'sb000000000000000000000000010000001000000000000000000000000000000000000;
		22734: Delta = 69'sb111111111111111111111111110000001000000000000000000000000000000000000;
		28127: Delta = 69'sb000000000000000000000000001111111000000000000000000000000000000000000;
		3068: Delta = 69'sb111111111111111111111111101111111000000000000000000000000000000000000;
		34892: Delta = 69'sb000000000000000000000000100000001000000000000000000000000000000000000;
		35635: Delta = 69'sb111111111111111111111111100000001000000000000000000000000000000000000;
		15226: Delta = 69'sb000000000000000000000000011111111000000000000000000000000000000000000;
		15969: Delta = 69'sb111111111111111111111111011111111000000000000000000000000000000000000;
		9090: Delta = 69'sb000000000000000000000001000000001000000000000000000000000000000000000;
		10576: Delta = 69'sb111111111111111111111111000000001000000000000000000000000000000000000;
		40285: Delta = 69'sb000000000000000000000000111111111000000000000000000000000000000000000;
		41771: Delta = 69'sb111111111111111111111110111111111000000000000000000000000000000000000;
		8347: Delta = 69'sb000000000000000000000010000000001000000000000000000000000000000000000;
		11319: Delta = 69'sb111111111111111111111110000000001000000000000000000000000000000000000;
		39542: Delta = 69'sb000000000000000000000001111111111000000000000000000000000000000000000;
		42514: Delta = 69'sb111111111111111111111101111111111000000000000000000000000000000000000;
		6861: Delta = 69'sb000000000000000000000100000000001000000000000000000000000000000000000;
		12805: Delta = 69'sb111111111111111111111100000000001000000000000000000000000000000000000;
		38056: Delta = 69'sb000000000000000000000011111111111000000000000000000000000000000000000;
		44000: Delta = 69'sb111111111111111111111011111111111000000000000000000000000000000000000;
		3889: Delta = 69'sb000000000000000000001000000000001000000000000000000000000000000000000;
		15777: Delta = 69'sb111111111111111111111000000000001000000000000000000000000000000000000;
		35084: Delta = 69'sb000000000000000000000111111111111000000000000000000000000000000000000;
		46972: Delta = 69'sb111111111111111111110111111111111000000000000000000000000000000000000;
		48806: Delta = 69'sb000000000000000000010000000000001000000000000000000000000000000000000;
		21721: Delta = 69'sb111111111111111111110000000000001000000000000000000000000000000000000;
		29140: Delta = 69'sb000000000000000000001111111111111000000000000000000000000000000000000;
		2055: Delta = 69'sb111111111111111111101111111111111000000000000000000000000000000000000;
		36918: Delta = 69'sb000000000000000000100000000000001000000000000000000000000000000000000;
		33609: Delta = 69'sb111111111111111111100000000000001000000000000000000000000000000000000;
		17252: Delta = 69'sb000000000000000000011111111111111000000000000000000000000000000000000;
		13943: Delta = 69'sb111111111111111111011111111111111000000000000000000000000000000000000;
		13142: Delta = 69'sb000000000000000001000000000000001000000000000000000000000000000000000;
		6524: Delta = 69'sb111111111111111111000000000000001000000000000000000000000000000000000;
		44337: Delta = 69'sb000000000000000000111111111111111000000000000000000000000000000000000;
		37719: Delta = 69'sb111111111111111110111111111111111000000000000000000000000000000000000;
		16451: Delta = 69'sb000000000000000010000000000000001000000000000000000000000000000000000;
		3215: Delta = 69'sb111111111111111110000000000000001000000000000000000000000000000000000;
		47646: Delta = 69'sb000000000000000001111111111111111000000000000000000000000000000000000;
		34410: Delta = 69'sb111111111111111101111111111111111000000000000000000000000000000000000;
		23069: Delta = 69'sb000000000000000100000000000000001000000000000000000000000000000000000;
		47458: Delta = 69'sb111111111111111100000000000000001000000000000000000000000000000000000;
		3403: Delta = 69'sb000000000000000011111111111111111000000000000000000000000000000000000;
		27792: Delta = 69'sb111111111111111011111111111111111000000000000000000000000000000000000;
		36305: Delta = 69'sb000000000000001000000000000000001000000000000000000000000000000000000;
		34222: Delta = 69'sb111111111111111000000000000000001000000000000000000000000000000000000;
		16639: Delta = 69'sb000000000000000111111111111111111000000000000000000000000000000000000;
		14556: Delta = 69'sb111111111111110111111111111111111000000000000000000000000000000000000;
		11916: Delta = 69'sb000000000000010000000000000000001000000000000000000000000000000000000;
		7750: Delta = 69'sb111111111111110000000000000000001000000000000000000000000000000000000;
		43111: Delta = 69'sb000000000000001111111111111111111000000000000000000000000000000000000;
		38945: Delta = 69'sb111111111111101111111111111111111000000000000000000000000000000000000;
		13999: Delta = 69'sb000000000000100000000000000000001000000000000000000000000000000000000;
		5667: Delta = 69'sb111111111111100000000000000000001000000000000000000000000000000000000;
		45194: Delta = 69'sb000000000000011111111111111111111000000000000000000000000000000000000;
		36862: Delta = 69'sb111111111111011111111111111111111000000000000000000000000000000000000;
		18165: Delta = 69'sb000000000001000000000000000000001000000000000000000000000000000000000;
		1501: Delta = 69'sb111111111111000000000000000000001000000000000000000000000000000000000;
		49360: Delta = 69'sb000000000000111111111111111111111000000000000000000000000000000000000;
		32696: Delta = 69'sb111111111110111111111111111111111000000000000000000000000000000000000;
		26497: Delta = 69'sb000000000010000000000000000000001000000000000000000000000000000000000;
		44030: Delta = 69'sb111111111110000000000000000000001000000000000000000000000000000000000;
		6831: Delta = 69'sb000000000001111111111111111111111000000000000000000000000000000000000;
		24364: Delta = 69'sb111111111101111111111111111111111000000000000000000000000000000000000;
		43161: Delta = 69'sb000000000100000000000000000000001000000000000000000000000000000000000;
		27366: Delta = 69'sb111111111100000000000000000000001000000000000000000000000000000000000;
		23495: Delta = 69'sb000000000011111111111111111111111000000000000000000000000000000000000;
		7700: Delta = 69'sb111111111011111111111111111111111000000000000000000000000000000000000;
		25628: Delta = 69'sb000000001000000000000000000000001000000000000000000000000000000000000;
		44899: Delta = 69'sb111111111000000000000000000000001000000000000000000000000000000000000;
		5962: Delta = 69'sb000000000111111111111111111111111000000000000000000000000000000000000;
		25233: Delta = 69'sb111111110111111111111111111111111000000000000000000000000000000000000;
		41423: Delta = 69'sb000000010000000000000000000000001000000000000000000000000000000000000;
		29104: Delta = 69'sb111111110000000000000000000000001000000000000000000000000000000000000;
		21757: Delta = 69'sb000000001111111111111111111111111000000000000000000000000000000000000;
		9438: Delta = 69'sb111111101111111111111111111111111000000000000000000000000000000000000;
		22152: Delta = 69'sb000000100000000000000000000000001000000000000000000000000000000000000;
		48375: Delta = 69'sb111111100000000000000000000000001000000000000000000000000000000000000;
		2486: Delta = 69'sb000000011111111111111111111111111000000000000000000000000000000000000;
		28709: Delta = 69'sb111111011111111111111111111111111000000000000000000000000000000000000;
		34471: Delta = 69'sb000001000000000000000000000000001000000000000000000000000000000000000;
		36056: Delta = 69'sb111111000000000000000000000000001000000000000000000000000000000000000;
		14805: Delta = 69'sb000000111111111111111111111111111000000000000000000000000000000000000;
		16390: Delta = 69'sb111110111111111111111111111111111000000000000000000000000000000000000;
		8248: Delta = 69'sb000010000000000000000000000000001000000000000000000000000000000000000;
		11418: Delta = 69'sb111110000000000000000000000000001000000000000000000000000000000000000;
		39443: Delta = 69'sb000001111111111111111111111111111000000000000000000000000000000000000;
		42613: Delta = 69'sb111101111111111111111111111111111000000000000000000000000000000000000;
		6663: Delta = 69'sb000100000000000000000000000000001000000000000000000000000000000000000;
		13003: Delta = 69'sb111100000000000000000000000000001000000000000000000000000000000000000;
		37858: Delta = 69'sb000011111111111111111111111111111000000000000000000000000000000000000;
		44198: Delta = 69'sb111011111111111111111111111111111000000000000000000000000000000000000;
		3493: Delta = 69'sb001000000000000000000000000000001000000000000000000000000000000000000;
		16173: Delta = 69'sb111000000000000000000000000000001000000000000000000000000000000000000;
		34688: Delta = 69'sb000111111111111111111111111111111000000000000000000000000000000000000;
		47368: Delta = 69'sb110111111111111111111111111111111000000000000000000000000000000000000;
		48014: Delta = 69'sb010000000000000000000000000000001000000000000000000000000000000000000;
		22513: Delta = 69'sb110000000000000000000000000000001000000000000000000000000000000000000;
		28348: Delta = 69'sb001111111111111111111111111111111000000000000000000000000000000000000;
		2847: Delta = 69'sb101111111111111111111111111111111000000000000000000000000000000000000;
		8137: Delta = 69'sb000000000000000000000000000000110000000000000000000000000000000000000;
		42724: Delta = 69'sb111111111111111111111111111111010000000000000000000000000000000000000;
		47469: Delta = 69'sb000000000000000000000000000001010000000000000000000000000000000000000;
		3392: Delta = 69'sb111111111111111111111111111110110000000000000000000000000000000000000;
		24411: Delta = 69'sb000000000000000000000000000010010000000000000000000000000000000000000;
		14921: Delta = 69'sb111111111111111111111111111110010000000000000000000000000000000000000;
		35940: Delta = 69'sb000000000000000000000000000001110000000000000000000000000000000000000;
		26450: Delta = 69'sb111111111111111111111111111101110000000000000000000000000000000000000;
		29156: Delta = 69'sb000000000000000000000000000100010000000000000000000000000000000000000;
		10176: Delta = 69'sb111111111111111111111111111100010000000000000000000000000000000000000;
		40685: Delta = 69'sb000000000000000000000000000011110000000000000000000000000000000000000;
		21705: Delta = 69'sb111111111111111111111111111011110000000000000000000000000000000000000;
		38646: Delta = 69'sb000000000000000000000000001000010000000000000000000000000000000000000;
		686: Delta = 69'sb111111111111111111111111111000010000000000000000000000000000000000000;
		50175: Delta = 69'sb000000000000000000000000000111110000000000000000000000000000000000000;
		12215: Delta = 69'sb111111111111111111111111110111110000000000000000000000000000000000000;
		6765: Delta = 69'sb000000000000000000000000010000010000000000000000000000000000000000000;
		32567: Delta = 69'sb111111111111111111111111110000010000000000000000000000000000000000000;
		18294: Delta = 69'sb000000000000000000000000001111110000000000000000000000000000000000000;
		44096: Delta = 69'sb111111111111111111111111101111110000000000000000000000000000000000000;
		44725: Delta = 69'sb000000000000000000000000100000010000000000000000000000000000000000000;
		45468: Delta = 69'sb111111111111111111111111100000010000000000000000000000000000000000000;
		5393: Delta = 69'sb000000000000000000000000011111110000000000000000000000000000000000000;
		6136: Delta = 69'sb111111111111111111111111011111110000000000000000000000000000000000000;
		18923: Delta = 69'sb000000000000000000000001000000010000000000000000000000000000000000000;
		20409: Delta = 69'sb111111111111111111111111000000010000000000000000000000000000000000000;
		30452: Delta = 69'sb000000000000000000000000111111110000000000000000000000000000000000000;
		31938: Delta = 69'sb111111111111111111111110111111110000000000000000000000000000000000000;
		18180: Delta = 69'sb000000000000000000000010000000010000000000000000000000000000000000000;
		21152: Delta = 69'sb111111111111111111111110000000010000000000000000000000000000000000000;
		29709: Delta = 69'sb000000000000000000000001111111110000000000000000000000000000000000000;
		32681: Delta = 69'sb111111111111111111111101111111110000000000000000000000000000000000000;
		16694: Delta = 69'sb000000000000000000000100000000010000000000000000000000000000000000000;
		22638: Delta = 69'sb111111111111111111111100000000010000000000000000000000000000000000000;
		28223: Delta = 69'sb000000000000000000000011111111110000000000000000000000000000000000000;
		34167: Delta = 69'sb111111111111111111111011111111110000000000000000000000000000000000000;
		13722: Delta = 69'sb000000000000000000001000000000010000000000000000000000000000000000000;
		25610: Delta = 69'sb111111111111111111111000000000010000000000000000000000000000000000000;
		25251: Delta = 69'sb000000000000000000000111111111110000000000000000000000000000000000000;
		37139: Delta = 69'sb111111111111111111110111111111110000000000000000000000000000000000000;
		7778: Delta = 69'sb000000000000000000010000000000010000000000000000000000000000000000000;
		31554: Delta = 69'sb111111111111111111110000000000010000000000000000000000000000000000000;
		19307: Delta = 69'sb000000000000000000001111111111110000000000000000000000000000000000000;
		43083: Delta = 69'sb111111111111111111101111111111110000000000000000000000000000000000000;
		46751: Delta = 69'sb000000000000000000100000000000010000000000000000000000000000000000000;
		43442: Delta = 69'sb111111111111111111100000000000010000000000000000000000000000000000000;
		7419: Delta = 69'sb000000000000000000011111111111110000000000000000000000000000000000000;
		4110: Delta = 69'sb111111111111111111011111111111110000000000000000000000000000000000000;
		22975: Delta = 69'sb000000000000000001000000000000010000000000000000000000000000000000000;
		16357: Delta = 69'sb111111111111111111000000000000010000000000000000000000000000000000000;
		34504: Delta = 69'sb000000000000000000111111111111110000000000000000000000000000000000000;
		27886: Delta = 69'sb111111111111111110111111111111110000000000000000000000000000000000000;
		26284: Delta = 69'sb000000000000000010000000000000010000000000000000000000000000000000000;
		13048: Delta = 69'sb111111111111111110000000000000010000000000000000000000000000000000000;
		37813: Delta = 69'sb000000000000000001111111111111110000000000000000000000000000000000000;
		24577: Delta = 69'sb111111111111111101111111111111110000000000000000000000000000000000000;
		32902: Delta = 69'sb000000000000000100000000000000010000000000000000000000000000000000000;
		6430: Delta = 69'sb111111111111111100000000000000010000000000000000000000000000000000000;
		44431: Delta = 69'sb000000000000000011111111111111110000000000000000000000000000000000000;
		17959: Delta = 69'sb111111111111111011111111111111110000000000000000000000000000000000000;
		46138: Delta = 69'sb000000000000001000000000000000010000000000000000000000000000000000000;
		44055: Delta = 69'sb111111111111111000000000000000010000000000000000000000000000000000000;
		6806: Delta = 69'sb000000000000000111111111111111110000000000000000000000000000000000000;
		4723: Delta = 69'sb111111111111110111111111111111110000000000000000000000000000000000000;
		21749: Delta = 69'sb000000000000010000000000000000010000000000000000000000000000000000000;
		17583: Delta = 69'sb111111111111110000000000000000010000000000000000000000000000000000000;
		33278: Delta = 69'sb000000000000001111111111111111110000000000000000000000000000000000000;
		29112: Delta = 69'sb111111111111101111111111111111110000000000000000000000000000000000000;
		23832: Delta = 69'sb000000000000100000000000000000010000000000000000000000000000000000000;
		15500: Delta = 69'sb111111111111100000000000000000010000000000000000000000000000000000000;
		35361: Delta = 69'sb000000000000011111111111111111110000000000000000000000000000000000000;
		27029: Delta = 69'sb111111111111011111111111111111110000000000000000000000000000000000000;
		27998: Delta = 69'sb000000000001000000000000000000010000000000000000000000000000000000000;
		11334: Delta = 69'sb111111111111000000000000000000010000000000000000000000000000000000000;
		39527: Delta = 69'sb000000000000111111111111111111110000000000000000000000000000000000000;
		22863: Delta = 69'sb111111111110111111111111111111110000000000000000000000000000000000000;
		36330: Delta = 69'sb000000000010000000000000000000010000000000000000000000000000000000000;
		3002: Delta = 69'sb111111111110000000000000000000010000000000000000000000000000000000000;
		47859: Delta = 69'sb000000000001111111111111111111110000000000000000000000000000000000000;
		14531: Delta = 69'sb111111111101111111111111111111110000000000000000000000000000000000000;
		2133: Delta = 69'sb000000000100000000000000000000010000000000000000000000000000000000000;
		37199: Delta = 69'sb111111111100000000000000000000010000000000000000000000000000000000000;
		13662: Delta = 69'sb000000000011111111111111111111110000000000000000000000000000000000000;
		48728: Delta = 69'sb111111111011111111111111111111110000000000000000000000000000000000000;
		35461: Delta = 69'sb000000001000000000000000000000010000000000000000000000000000000000000;
		3871: Delta = 69'sb111111111000000000000000000000010000000000000000000000000000000000000;
		46990: Delta = 69'sb000000000111111111111111111111110000000000000000000000000000000000000;
		15400: Delta = 69'sb111111110111111111111111111111110000000000000000000000000000000000000;
		395: Delta = 69'sb000000010000000000000000000000010000000000000000000000000000000000000;
		38937: Delta = 69'sb111111110000000000000000000000010000000000000000000000000000000000000;
		11924: Delta = 69'sb000000001111111111111111111111110000000000000000000000000000000000000;
		50466: Delta = 69'sb111111101111111111111111111111110000000000000000000000000000000000000;
		31985: Delta = 69'sb000000100000000000000000000000010000000000000000000000000000000000000;
		7347: Delta = 69'sb111111100000000000000000000000010000000000000000000000000000000000000;
		43514: Delta = 69'sb000000011111111111111111111111110000000000000000000000000000000000000;
		18876: Delta = 69'sb111111011111111111111111111111110000000000000000000000000000000000000;
		44304: Delta = 69'sb000001000000000000000000000000010000000000000000000000000000000000000;
		45889: Delta = 69'sb111111000000000000000000000000010000000000000000000000000000000000000;
		4972: Delta = 69'sb000000111111111111111111111111110000000000000000000000000000000000000;
		6557: Delta = 69'sb111110111111111111111111111111110000000000000000000000000000000000000;
		18081: Delta = 69'sb000010000000000000000000000000010000000000000000000000000000000000000;
		21251: Delta = 69'sb111110000000000000000000000000010000000000000000000000000000000000000;
		29610: Delta = 69'sb000001111111111111111111111111110000000000000000000000000000000000000;
		32780: Delta = 69'sb111101111111111111111111111111110000000000000000000000000000000000000;
		16496: Delta = 69'sb000100000000000000000000000000010000000000000000000000000000000000000;
		22836: Delta = 69'sb111100000000000000000000000000010000000000000000000000000000000000000;
		28025: Delta = 69'sb000011111111111111111111111111110000000000000000000000000000000000000;
		34365: Delta = 69'sb111011111111111111111111111111110000000000000000000000000000000000000;
		13326: Delta = 69'sb001000000000000000000000000000010000000000000000000000000000000000000;
		26006: Delta = 69'sb111000000000000000000000000000010000000000000000000000000000000000000;
		24855: Delta = 69'sb000111111111111111111111111111110000000000000000000000000000000000000;
		37535: Delta = 69'sb110111111111111111111111111111110000000000000000000000000000000000000;
		6986: Delta = 69'sb010000000000000000000000000000010000000000000000000000000000000000000;
		32346: Delta = 69'sb110000000000000000000000000000010000000000000000000000000000000000000;
		18515: Delta = 69'sb001111111111111111111111111111110000000000000000000000000000000000000;
		43875: Delta = 69'sb101111111111111111111111111111110000000000000000000000000000000000000;
		16274: Delta = 69'sb000000000000000000000000000001100000000000000000000000000000000000000;
		34587: Delta = 69'sb111111111111111111111111111110100000000000000000000000000000000000000;
		44077: Delta = 69'sb000000000000000000000000000010100000000000000000000000000000000000000;
		6784: Delta = 69'sb111111111111111111111111111101100000000000000000000000000000000000000;
		48822: Delta = 69'sb000000000000000000000000000100100000000000000000000000000000000000000;
		29842: Delta = 69'sb111111111111111111111111111100100000000000000000000000000000000000000;
		21019: Delta = 69'sb000000000000000000000000000011100000000000000000000000000000000000000;
		2039: Delta = 69'sb111111111111111111111111111011100000000000000000000000000000000000000;
		7451: Delta = 69'sb000000000000000000000000001000100000000000000000000000000000000000000;
		20352: Delta = 69'sb111111111111111111111111111000100000000000000000000000000000000000000;
		30509: Delta = 69'sb000000000000000000000000000111100000000000000000000000000000000000000;
		43410: Delta = 69'sb111111111111111111111111110111100000000000000000000000000000000000000;
		26431: Delta = 69'sb000000000000000000000000010000100000000000000000000000000000000000000;
		1372: Delta = 69'sb111111111111111111111111110000100000000000000000000000000000000000000;
		49489: Delta = 69'sb000000000000000000000000001111100000000000000000000000000000000000000;
		24430: Delta = 69'sb111111111111111111111111101111100000000000000000000000000000000000000;
		13530: Delta = 69'sb000000000000000000000000100000100000000000000000000000000000000000000;
		14273: Delta = 69'sb111111111111111111111111100000100000000000000000000000000000000000000;
		36588: Delta = 69'sb000000000000000000000000011111100000000000000000000000000000000000000;
		37331: Delta = 69'sb111111111111111111111111011111100000000000000000000000000000000000000;
		38589: Delta = 69'sb000000000000000000000001000000100000000000000000000000000000000000000;
		40075: Delta = 69'sb111111111111111111111111000000100000000000000000000000000000000000000;
		10786: Delta = 69'sb000000000000000000000000111111100000000000000000000000000000000000000;
		12272: Delta = 69'sb111111111111111111111110111111100000000000000000000000000000000000000;
		37846: Delta = 69'sb000000000000000000000010000000100000000000000000000000000000000000000;
		40818: Delta = 69'sb111111111111111111111110000000100000000000000000000000000000000000000;
		10043: Delta = 69'sb000000000000000000000001111111100000000000000000000000000000000000000;
		13015: Delta = 69'sb111111111111111111111101111111100000000000000000000000000000000000000;
		36360: Delta = 69'sb000000000000000000000100000000100000000000000000000000000000000000000;
		42304: Delta = 69'sb111111111111111111111100000000100000000000000000000000000000000000000;
		8557: Delta = 69'sb000000000000000000000011111111100000000000000000000000000000000000000;
		14501: Delta = 69'sb111111111111111111111011111111100000000000000000000000000000000000000;
		33388: Delta = 69'sb000000000000000000001000000000100000000000000000000000000000000000000;
		45276: Delta = 69'sb111111111111111111111000000000100000000000000000000000000000000000000;
		5585: Delta = 69'sb000000000000000000000111111111100000000000000000000000000000000000000;
		17473: Delta = 69'sb111111111111111111110111111111100000000000000000000000000000000000000;
		27444: Delta = 69'sb000000000000000000010000000000100000000000000000000000000000000000000;
		359: Delta = 69'sb111111111111111111110000000000100000000000000000000000000000000000000;
		50502: Delta = 69'sb000000000000000000001111111111100000000000000000000000000000000000000;
		23417: Delta = 69'sb111111111111111111101111111111100000000000000000000000000000000000000;
		15556: Delta = 69'sb000000000000000000100000000000100000000000000000000000000000000000000;
		12247: Delta = 69'sb111111111111111111100000000000100000000000000000000000000000000000000;
		38614: Delta = 69'sb000000000000000000011111111111100000000000000000000000000000000000000;
		35305: Delta = 69'sb111111111111111111011111111111100000000000000000000000000000000000000;
		42641: Delta = 69'sb000000000000000001000000000000100000000000000000000000000000000000000;
		36023: Delta = 69'sb111111111111111111000000000000100000000000000000000000000000000000000;
		14838: Delta = 69'sb000000000000000000111111111111100000000000000000000000000000000000000;
		8220: Delta = 69'sb111111111111111110111111111111100000000000000000000000000000000000000;
		45950: Delta = 69'sb000000000000000010000000000000100000000000000000000000000000000000000;
		32714: Delta = 69'sb111111111111111110000000000000100000000000000000000000000000000000000;
		18147: Delta = 69'sb000000000000000001111111111111100000000000000000000000000000000000000;
		4911: Delta = 69'sb111111111111111101111111111111100000000000000000000000000000000000000;
		1707: Delta = 69'sb000000000000000100000000000000100000000000000000000000000000000000000;
		26096: Delta = 69'sb111111111111111100000000000000100000000000000000000000000000000000000;
		24765: Delta = 69'sb000000000000000011111111111111100000000000000000000000000000000000000;
		49154: Delta = 69'sb111111111111111011111111111111100000000000000000000000000000000000000;
		14943: Delta = 69'sb000000000000001000000000000000100000000000000000000000000000000000000;
		12860: Delta = 69'sb111111111111111000000000000000100000000000000000000000000000000000000;
		38001: Delta = 69'sb000000000000000111111111111111100000000000000000000000000000000000000;
		35918: Delta = 69'sb111111111111110111111111111111100000000000000000000000000000000000000;
		41415: Delta = 69'sb000000000000010000000000000000100000000000000000000000000000000000000;
		37249: Delta = 69'sb111111111111110000000000000000100000000000000000000000000000000000000;
		13612: Delta = 69'sb000000000000001111111111111111100000000000000000000000000000000000000;
		9446: Delta = 69'sb111111111111101111111111111111100000000000000000000000000000000000000;
		43498: Delta = 69'sb000000000000100000000000000000100000000000000000000000000000000000000;
		35166: Delta = 69'sb111111111111100000000000000000100000000000000000000000000000000000000;
		15695: Delta = 69'sb000000000000011111111111111111100000000000000000000000000000000000000;
		7363: Delta = 69'sb111111111111011111111111111111100000000000000000000000000000000000000;
		47664: Delta = 69'sb000000000001000000000000000000100000000000000000000000000000000000000;
		31000: Delta = 69'sb111111111111000000000000000000100000000000000000000000000000000000000;
		19861: Delta = 69'sb000000000000111111111111111111100000000000000000000000000000000000000;
		3197: Delta = 69'sb111111111110111111111111111111100000000000000000000000000000000000000;
		5135: Delta = 69'sb000000000010000000000000000000100000000000000000000000000000000000000;
		22668: Delta = 69'sb111111111110000000000000000000100000000000000000000000000000000000000;
		28193: Delta = 69'sb000000000001111111111111111111100000000000000000000000000000000000000;
		45726: Delta = 69'sb111111111101111111111111111111100000000000000000000000000000000000000;
		21799: Delta = 69'sb000000000100000000000000000000100000000000000000000000000000000000000;
		6004: Delta = 69'sb111111111100000000000000000000100000000000000000000000000000000000000;
		44857: Delta = 69'sb000000000011111111111111111111100000000000000000000000000000000000000;
		29062: Delta = 69'sb111111111011111111111111111111100000000000000000000000000000000000000;
		4266: Delta = 69'sb000000001000000000000000000000100000000000000000000000000000000000000;
		23537: Delta = 69'sb111111111000000000000000000000100000000000000000000000000000000000000;
		27324: Delta = 69'sb000000000111111111111111111111100000000000000000000000000000000000000;
		46595: Delta = 69'sb111111110111111111111111111111100000000000000000000000000000000000000;
		20061: Delta = 69'sb000000010000000000000000000000100000000000000000000000000000000000000;
		7742: Delta = 69'sb111111110000000000000000000000100000000000000000000000000000000000000;
		43119: Delta = 69'sb000000001111111111111111111111100000000000000000000000000000000000000;
		30800: Delta = 69'sb111111101111111111111111111111100000000000000000000000000000000000000;
		790: Delta = 69'sb000000100000000000000000000000100000000000000000000000000000000000000;
		27013: Delta = 69'sb111111100000000000000000000000100000000000000000000000000000000000000;
		23848: Delta = 69'sb000000011111111111111111111111100000000000000000000000000000000000000;
		50071: Delta = 69'sb111111011111111111111111111111100000000000000000000000000000000000000;
		13109: Delta = 69'sb000001000000000000000000000000100000000000000000000000000000000000000;
		14694: Delta = 69'sb111111000000000000000000000000100000000000000000000000000000000000000;
		36167: Delta = 69'sb000000111111111111111111111111100000000000000000000000000000000000000;
		37752: Delta = 69'sb111110111111111111111111111111100000000000000000000000000000000000000;
		37747: Delta = 69'sb000010000000000000000000000000100000000000000000000000000000000000000;
		40917: Delta = 69'sb111110000000000000000000000000100000000000000000000000000000000000000;
		9944: Delta = 69'sb000001111111111111111111111111100000000000000000000000000000000000000;
		13114: Delta = 69'sb111101111111111111111111111111100000000000000000000000000000000000000;
		36162: Delta = 69'sb000100000000000000000000000000100000000000000000000000000000000000000;
		42502: Delta = 69'sb111100000000000000000000000000100000000000000000000000000000000000000;
		8359: Delta = 69'sb000011111111111111111111111111100000000000000000000000000000000000000;
		14699: Delta = 69'sb111011111111111111111111111111100000000000000000000000000000000000000;
		32992: Delta = 69'sb001000000000000000000000000000100000000000000000000000000000000000000;
		45672: Delta = 69'sb111000000000000000000000000000100000000000000000000000000000000000000;
		5189: Delta = 69'sb000111111111111111111111111111100000000000000000000000000000000000000;
		17869: Delta = 69'sb110111111111111111111111111111100000000000000000000000000000000000000;
		26652: Delta = 69'sb010000000000000000000000000000100000000000000000000000000000000000000;
		1151: Delta = 69'sb110000000000000000000000000000100000000000000000000000000000000000000;
		49710: Delta = 69'sb001111111111111111111111111111100000000000000000000000000000000000000;
		24209: Delta = 69'sb101111111111111111111111111111100000000000000000000000000000000000000;
		32548: Delta = 69'sb000000000000000000000000000011000000000000000000000000000000000000000;
		18313: Delta = 69'sb111111111111111111111111111101000000000000000000000000000000000000000;
		37293: Delta = 69'sb000000000000000000000000000101000000000000000000000000000000000000000;
		13568: Delta = 69'sb111111111111111111111111111011000000000000000000000000000000000000000;
		46783: Delta = 69'sb000000000000000000000000001001000000000000000000000000000000000000000;
		8823: Delta = 69'sb111111111111111111111111111001000000000000000000000000000000000000000;
		42038: Delta = 69'sb000000000000000000000000000111000000000000000000000000000000000000000;
		4078: Delta = 69'sb111111111111111111111111110111000000000000000000000000000000000000000;
		14902: Delta = 69'sb000000000000000000000000010001000000000000000000000000000000000000000;
		40704: Delta = 69'sb111111111111111111111111110001000000000000000000000000000000000000000;
		10157: Delta = 69'sb000000000000000000000000001111000000000000000000000000000000000000000;
		35959: Delta = 69'sb111111111111111111111111101111000000000000000000000000000000000000000;
		2001: Delta = 69'sb000000000000000000000000100001000000000000000000000000000000000000000;
		2744: Delta = 69'sb111111111111111111111111100001000000000000000000000000000000000000000;
		48117: Delta = 69'sb000000000000000000000000011111000000000000000000000000000000000000000;
		48860: Delta = 69'sb111111111111111111111111011111000000000000000000000000000000000000000;
		27060: Delta = 69'sb000000000000000000000001000001000000000000000000000000000000000000000;
		28546: Delta = 69'sb111111111111111111111111000001000000000000000000000000000000000000000;
		22315: Delta = 69'sb000000000000000000000000111111000000000000000000000000000000000000000;
		23801: Delta = 69'sb111111111111111111111110111111000000000000000000000000000000000000000;
		26317: Delta = 69'sb000000000000000000000010000001000000000000000000000000000000000000000;
		29289: Delta = 69'sb111111111111111111111110000001000000000000000000000000000000000000000;
		21572: Delta = 69'sb000000000000000000000001111111000000000000000000000000000000000000000;
		24544: Delta = 69'sb111111111111111111111101111111000000000000000000000000000000000000000;
		24831: Delta = 69'sb000000000000000000000100000001000000000000000000000000000000000000000;
		30775: Delta = 69'sb111111111111111111111100000001000000000000000000000000000000000000000;
		20086: Delta = 69'sb000000000000000000000011111111000000000000000000000000000000000000000;
		26030: Delta = 69'sb111111111111111111111011111111000000000000000000000000000000000000000;
		21859: Delta = 69'sb000000000000000000001000000001000000000000000000000000000000000000000;
		33747: Delta = 69'sb111111111111111111111000000001000000000000000000000000000000000000000;
		17114: Delta = 69'sb000000000000000000000111111111000000000000000000000000000000000000000;
		29002: Delta = 69'sb111111111111111111110111111111000000000000000000000000000000000000000;
		15915: Delta = 69'sb000000000000000000010000000001000000000000000000000000000000000000000;
		39691: Delta = 69'sb111111111111111111110000000001000000000000000000000000000000000000000;
		11170: Delta = 69'sb000000000000000000001111111111000000000000000000000000000000000000000;
		34946: Delta = 69'sb111111111111111111101111111111000000000000000000000000000000000000000;
		4027: Delta = 69'sb000000000000000000100000000001000000000000000000000000000000000000000;
		718: Delta = 69'sb111111111111111111100000000001000000000000000000000000000000000000000;
		50143: Delta = 69'sb000000000000000000011111111111000000000000000000000000000000000000000;
		46834: Delta = 69'sb111111111111111111011111111111000000000000000000000000000000000000000;
		31112: Delta = 69'sb000000000000000001000000000001000000000000000000000000000000000000000;
		24494: Delta = 69'sb111111111111111111000000000001000000000000000000000000000000000000000;
		26367: Delta = 69'sb000000000000000000111111111111000000000000000000000000000000000000000;
		19749: Delta = 69'sb111111111111111110111111111111000000000000000000000000000000000000000;
		34421: Delta = 69'sb000000000000000010000000000001000000000000000000000000000000000000000;
		21185: Delta = 69'sb111111111111111110000000000001000000000000000000000000000000000000000;
		29676: Delta = 69'sb000000000000000001111111111111000000000000000000000000000000000000000;
		16440: Delta = 69'sb111111111111111101111111111111000000000000000000000000000000000000000;
		41039: Delta = 69'sb000000000000000100000000000001000000000000000000000000000000000000000;
		14567: Delta = 69'sb111111111111111100000000000001000000000000000000000000000000000000000;
		36294: Delta = 69'sb000000000000000011111111111111000000000000000000000000000000000000000;
		9822: Delta = 69'sb111111111111111011111111111111000000000000000000000000000000000000000;
		3414: Delta = 69'sb000000000000001000000000000001000000000000000000000000000000000000000;
		1331: Delta = 69'sb111111111111111000000000000001000000000000000000000000000000000000000;
		49530: Delta = 69'sb000000000000000111111111111111000000000000000000000000000000000000000;
		47447: Delta = 69'sb111111111111110111111111111111000000000000000000000000000000000000000;
		29886: Delta = 69'sb000000000000010000000000000001000000000000000000000000000000000000000;
		25720: Delta = 69'sb111111111111110000000000000001000000000000000000000000000000000000000;
		25141: Delta = 69'sb000000000000001111111111111111000000000000000000000000000000000000000;
		20975: Delta = 69'sb111111111111101111111111111111000000000000000000000000000000000000000;
		31969: Delta = 69'sb000000000000100000000000000001000000000000000000000000000000000000000;
		23637: Delta = 69'sb111111111111100000000000000001000000000000000000000000000000000000000;
		27224: Delta = 69'sb000000000000011111111111111111000000000000000000000000000000000000000;
		18892: Delta = 69'sb111111111111011111111111111111000000000000000000000000000000000000000;
		36135: Delta = 69'sb000000000001000000000000000001000000000000000000000000000000000000000;
		19471: Delta = 69'sb111111111111000000000000000001000000000000000000000000000000000000000;
		31390: Delta = 69'sb000000000000111111111111111111000000000000000000000000000000000000000;
		14726: Delta = 69'sb111111111110111111111111111111000000000000000000000000000000000000000;
		44467: Delta = 69'sb000000000010000000000000000001000000000000000000000000000000000000000;
		11139: Delta = 69'sb111111111110000000000000000001000000000000000000000000000000000000000;
		39722: Delta = 69'sb000000000001111111111111111111000000000000000000000000000000000000000;
		6394: Delta = 69'sb111111111101111111111111111111000000000000000000000000000000000000000;
		10270: Delta = 69'sb000000000100000000000000000001000000000000000000000000000000000000000;
		45336: Delta = 69'sb111111111100000000000000000001000000000000000000000000000000000000000;
		5525: Delta = 69'sb000000000011111111111111111111000000000000000000000000000000000000000;
		40591: Delta = 69'sb111111111011111111111111111111000000000000000000000000000000000000000;
		43598: Delta = 69'sb000000001000000000000000000001000000000000000000000000000000000000000;
		12008: Delta = 69'sb111111111000000000000000000001000000000000000000000000000000000000000;
		38853: Delta = 69'sb000000000111111111111111111111000000000000000000000000000000000000000;
		7263: Delta = 69'sb111111110111111111111111111111000000000000000000000000000000000000000;
		8532: Delta = 69'sb000000010000000000000000000001000000000000000000000000000000000000000;
		47074: Delta = 69'sb111111110000000000000000000001000000000000000000000000000000000000000;
		3787: Delta = 69'sb000000001111111111111111111111000000000000000000000000000000000000000;
		42329: Delta = 69'sb111111101111111111111111111111000000000000000000000000000000000000000;
		40122: Delta = 69'sb000000100000000000000000000001000000000000000000000000000000000000000;
		15484: Delta = 69'sb111111100000000000000000000001000000000000000000000000000000000000000;
		35377: Delta = 69'sb000000011111111111111111111111000000000000000000000000000000000000000;
		10739: Delta = 69'sb111111011111111111111111111111000000000000000000000000000000000000000;
		1580: Delta = 69'sb000001000000000000000000000001000000000000000000000000000000000000000;
		3165: Delta = 69'sb111111000000000000000000000001000000000000000000000000000000000000000;
		47696: Delta = 69'sb000000111111111111111111111111000000000000000000000000000000000000000;
		49281: Delta = 69'sb111110111111111111111111111111000000000000000000000000000000000000000;
		26218: Delta = 69'sb000010000000000000000000000001000000000000000000000000000000000000000;
		29388: Delta = 69'sb111110000000000000000000000001000000000000000000000000000000000000000;
		21473: Delta = 69'sb000001111111111111111111111111000000000000000000000000000000000000000;
		24643: Delta = 69'sb111101111111111111111111111111000000000000000000000000000000000000000;
		24633: Delta = 69'sb000100000000000000000000000001000000000000000000000000000000000000000;
		30973: Delta = 69'sb111100000000000000000000000001000000000000000000000000000000000000000;
		19888: Delta = 69'sb000011111111111111111111111111000000000000000000000000000000000000000;
		26228: Delta = 69'sb111011111111111111111111111111000000000000000000000000000000000000000;
		21463: Delta = 69'sb001000000000000000000000000001000000000000000000000000000000000000000;
		34143: Delta = 69'sb111000000000000000000000000001000000000000000000000000000000000000000;
		16718: Delta = 69'sb000111111111111111111111111111000000000000000000000000000000000000000;
		29398: Delta = 69'sb110111111111111111111111111111000000000000000000000000000000000000000;
		15123: Delta = 69'sb010000000000000000000000000001000000000000000000000000000000000000000;
		40483: Delta = 69'sb110000000000000000000000000001000000000000000000000000000000000000000;
		10378: Delta = 69'sb001111111111111111111111111111000000000000000000000000000000000000000;
		35738: Delta = 69'sb101111111111111111111111111111000000000000000000000000000000000000000;
		14235: Delta = 69'sb000000000000000000000000000110000000000000000000000000000000000000000;
		36626: Delta = 69'sb111111111111111111111111111010000000000000000000000000000000000000000;
		23725: Delta = 69'sb000000000000000000000000001010000000000000000000000000000000000000000;
		27136: Delta = 69'sb111111111111111111111111110110000000000000000000000000000000000000000;
		42705: Delta = 69'sb000000000000000000000000010010000000000000000000000000000000000000000;
		17646: Delta = 69'sb111111111111111111111111110010000000000000000000000000000000000000000;
		33215: Delta = 69'sb000000000000000000000000001110000000000000000000000000000000000000000;
		8156: Delta = 69'sb111111111111111111111111101110000000000000000000000000000000000000000;
		29804: Delta = 69'sb000000000000000000000000100010000000000000000000000000000000000000000;
		30547: Delta = 69'sb111111111111111111111111100010000000000000000000000000000000000000000;
		20314: Delta = 69'sb000000000000000000000000011110000000000000000000000000000000000000000;
		21057: Delta = 69'sb111111111111111111111111011110000000000000000000000000000000000000000;
		4002: Delta = 69'sb000000000000000000000001000010000000000000000000000000000000000000000;
		5488: Delta = 69'sb111111111111111111111111000010000000000000000000000000000000000000000;
		45373: Delta = 69'sb000000000000000000000000111110000000000000000000000000000000000000000;
		46859: Delta = 69'sb111111111111111111111110111110000000000000000000000000000000000000000;
		3259: Delta = 69'sb000000000000000000000010000010000000000000000000000000000000000000000;
		6231: Delta = 69'sb111111111111111111111110000010000000000000000000000000000000000000000;
		44630: Delta = 69'sb000000000000000000000001111110000000000000000000000000000000000000000;
		47602: Delta = 69'sb111111111111111111111101111110000000000000000000000000000000000000000;
		1773: Delta = 69'sb000000000000000000000100000010000000000000000000000000000000000000000;
		7717: Delta = 69'sb111111111111111111111100000010000000000000000000000000000000000000000;
		43144: Delta = 69'sb000000000000000000000011111110000000000000000000000000000000000000000;
		49088: Delta = 69'sb111111111111111111111011111110000000000000000000000000000000000000000;
		49662: Delta = 69'sb000000000000000000001000000010000000000000000000000000000000000000000;
		10689: Delta = 69'sb111111111111111111111000000010000000000000000000000000000000000000000;
		40172: Delta = 69'sb000000000000000000000111111110000000000000000000000000000000000000000;
		1199: Delta = 69'sb111111111111111111110111111110000000000000000000000000000000000000000;
		43718: Delta = 69'sb000000000000000000010000000010000000000000000000000000000000000000000;
		16633: Delta = 69'sb111111111111111111110000000010000000000000000000000000000000000000000;
		34228: Delta = 69'sb000000000000000000001111111110000000000000000000000000000000000000000;
		7143: Delta = 69'sb111111111111111111101111111110000000000000000000000000000000000000000;
		31830: Delta = 69'sb000000000000000000100000000010000000000000000000000000000000000000000;
		28521: Delta = 69'sb111111111111111111100000000010000000000000000000000000000000000000000;
		22340: Delta = 69'sb000000000000000000011111111110000000000000000000000000000000000000000;
		19031: Delta = 69'sb111111111111111111011111111110000000000000000000000000000000000000000;
		8054: Delta = 69'sb000000000000000001000000000010000000000000000000000000000000000000000;
		1436: Delta = 69'sb111111111111111111000000000010000000000000000000000000000000000000000;
		49425: Delta = 69'sb000000000000000000111111111110000000000000000000000000000000000000000;
		42807: Delta = 69'sb111111111111111110111111111110000000000000000000000000000000000000000;
		11363: Delta = 69'sb000000000000000010000000000010000000000000000000000000000000000000000;
		48988: Delta = 69'sb111111111111111110000000000010000000000000000000000000000000000000000;
		1873: Delta = 69'sb000000000000000001111111111110000000000000000000000000000000000000000;
		39498: Delta = 69'sb111111111111111101111111111110000000000000000000000000000000000000000;
		17981: Delta = 69'sb000000000000000100000000000010000000000000000000000000000000000000000;
		42370: Delta = 69'sb111111111111111100000000000010000000000000000000000000000000000000000;
		8491: Delta = 69'sb000000000000000011111111111110000000000000000000000000000000000000000;
		32880: Delta = 69'sb111111111111111011111111111110000000000000000000000000000000000000000;
		31217: Delta = 69'sb000000000000001000000000000010000000000000000000000000000000000000000;
		29134: Delta = 69'sb111111111111111000000000000010000000000000000000000000000000000000000;
		21727: Delta = 69'sb000000000000000111111111111110000000000000000000000000000000000000000;
		19644: Delta = 69'sb111111111111110111111111111110000000000000000000000000000000000000000;
		6828: Delta = 69'sb000000000000010000000000000010000000000000000000000000000000000000000;
		2662: Delta = 69'sb111111111111110000000000000010000000000000000000000000000000000000000;
		48199: Delta = 69'sb000000000000001111111111111110000000000000000000000000000000000000000;
		44033: Delta = 69'sb111111111111101111111111111110000000000000000000000000000000000000000;
		8911: Delta = 69'sb000000000000100000000000000010000000000000000000000000000000000000000;
		579: Delta = 69'sb111111111111100000000000000010000000000000000000000000000000000000000;
		50282: Delta = 69'sb000000000000011111111111111110000000000000000000000000000000000000000;
		41950: Delta = 69'sb111111111111011111111111111110000000000000000000000000000000000000000;
		13077: Delta = 69'sb000000000001000000000000000010000000000000000000000000000000000000000;
		47274: Delta = 69'sb111111111111000000000000000010000000000000000000000000000000000000000;
		3587: Delta = 69'sb000000000000111111111111111110000000000000000000000000000000000000000;
		37784: Delta = 69'sb111111111110111111111111111110000000000000000000000000000000000000000;
		21409: Delta = 69'sb000000000010000000000000000010000000000000000000000000000000000000000;
		38942: Delta = 69'sb111111111110000000000000000010000000000000000000000000000000000000000;
		11919: Delta = 69'sb000000000001111111111111111110000000000000000000000000000000000000000;
		29452: Delta = 69'sb111111111101111111111111111110000000000000000000000000000000000000000;
		38073: Delta = 69'sb000000000100000000000000000010000000000000000000000000000000000000000;
		22278: Delta = 69'sb111111111100000000000000000010000000000000000000000000000000000000000;
		28583: Delta = 69'sb000000000011111111111111111110000000000000000000000000000000000000000;
		12788: Delta = 69'sb111111111011111111111111111110000000000000000000000000000000000000000;
		20540: Delta = 69'sb000000001000000000000000000010000000000000000000000000000000000000000;
		39811: Delta = 69'sb111111111000000000000000000010000000000000000000000000000000000000000;
		11050: Delta = 69'sb000000000111111111111111111110000000000000000000000000000000000000000;
		30321: Delta = 69'sb111111110111111111111111111110000000000000000000000000000000000000000;
		36335: Delta = 69'sb000000010000000000000000000010000000000000000000000000000000000000000;
		24016: Delta = 69'sb111111110000000000000000000010000000000000000000000000000000000000000;
		26845: Delta = 69'sb000000001111111111111111111110000000000000000000000000000000000000000;
		14526: Delta = 69'sb111111101111111111111111111110000000000000000000000000000000000000000;
		17064: Delta = 69'sb000000100000000000000000000010000000000000000000000000000000000000000;
		43287: Delta = 69'sb111111100000000000000000000010000000000000000000000000000000000000000;
		7574: Delta = 69'sb000000011111111111111111111110000000000000000000000000000000000000000;
		33797: Delta = 69'sb111111011111111111111111111110000000000000000000000000000000000000000;
		29383: Delta = 69'sb000001000000000000000000000010000000000000000000000000000000000000000;
		30968: Delta = 69'sb111111000000000000000000000010000000000000000000000000000000000000000;
		19893: Delta = 69'sb000000111111111111111111111110000000000000000000000000000000000000000;
		21478: Delta = 69'sb111110111111111111111111111110000000000000000000000000000000000000000;
		3160: Delta = 69'sb000010000000000000000000000010000000000000000000000000000000000000000;
		6330: Delta = 69'sb111110000000000000000000000010000000000000000000000000000000000000000;
		44531: Delta = 69'sb000001111111111111111111111110000000000000000000000000000000000000000;
		47701: Delta = 69'sb111101111111111111111111111110000000000000000000000000000000000000000;
		1575: Delta = 69'sb000100000000000000000000000010000000000000000000000000000000000000000;
		7915: Delta = 69'sb111100000000000000000000000010000000000000000000000000000000000000000;
		42946: Delta = 69'sb000011111111111111111111111110000000000000000000000000000000000000000;
		49286: Delta = 69'sb111011111111111111111111111110000000000000000000000000000000000000000;
		49266: Delta = 69'sb001000000000000000000000000010000000000000000000000000000000000000000;
		11085: Delta = 69'sb111000000000000000000000000010000000000000000000000000000000000000000;
		39776: Delta = 69'sb000111111111111111111111111110000000000000000000000000000000000000000;
		1595: Delta = 69'sb110111111111111111111111111110000000000000000000000000000000000000000;
		42926: Delta = 69'sb010000000000000000000000000010000000000000000000000000000000000000000;
		17425: Delta = 69'sb110000000000000000000000000010000000000000000000000000000000000000000;
		33436: Delta = 69'sb001111111111111111111111111110000000000000000000000000000000000000000;
		7935: Delta = 69'sb101111111111111111111111111110000000000000000000000000000000000000000;
		28470: Delta = 69'sb000000000000000000000000001100000000000000000000000000000000000000000;
		22391: Delta = 69'sb111111111111111111111111110100000000000000000000000000000000000000000;
		47450: Delta = 69'sb000000000000000000000000010100000000000000000000000000000000000000000;
		3411: Delta = 69'sb111111111111111111111111101100000000000000000000000000000000000000000;
		34549: Delta = 69'sb000000000000000000000000100100000000000000000000000000000000000000000;
		35292: Delta = 69'sb111111111111111111111111100100000000000000000000000000000000000000000;
		15569: Delta = 69'sb000000000000000000000000011100000000000000000000000000000000000000000;
		16312: Delta = 69'sb111111111111111111111111011100000000000000000000000000000000000000000;
		8747: Delta = 69'sb000000000000000000000001000100000000000000000000000000000000000000000;
		10233: Delta = 69'sb111111111111111111111111000100000000000000000000000000000000000000000;
		40628: Delta = 69'sb000000000000000000000000111100000000000000000000000000000000000000000;
		42114: Delta = 69'sb111111111111111111111110111100000000000000000000000000000000000000000;
		8004: Delta = 69'sb000000000000000000000010000100000000000000000000000000000000000000000;
		10976: Delta = 69'sb111111111111111111111110000100000000000000000000000000000000000000000;
		39885: Delta = 69'sb000000000000000000000001111100000000000000000000000000000000000000000;
		42857: Delta = 69'sb111111111111111111111101111100000000000000000000000000000000000000000;
		6518: Delta = 69'sb000000000000000000000100000100000000000000000000000000000000000000000;
		12462: Delta = 69'sb111111111111111111111100000100000000000000000000000000000000000000000;
		38399: Delta = 69'sb000000000000000000000011111100000000000000000000000000000000000000000;
		44343: Delta = 69'sb111111111111111111111011111100000000000000000000000000000000000000000;
		3546: Delta = 69'sb000000000000000000001000000100000000000000000000000000000000000000000;
		15434: Delta = 69'sb111111111111111111111000000100000000000000000000000000000000000000000;
		35427: Delta = 69'sb000000000000000000000111111100000000000000000000000000000000000000000;
		47315: Delta = 69'sb111111111111111111110111111100000000000000000000000000000000000000000;
		48463: Delta = 69'sb000000000000000000010000000100000000000000000000000000000000000000000;
		21378: Delta = 69'sb111111111111111111110000000100000000000000000000000000000000000000000;
		29483: Delta = 69'sb000000000000000000001111111100000000000000000000000000000000000000000;
		2398: Delta = 69'sb111111111111111111101111111100000000000000000000000000000000000000000;
		36575: Delta = 69'sb000000000000000000100000000100000000000000000000000000000000000000000;
		33266: Delta = 69'sb111111111111111111100000000100000000000000000000000000000000000000000;
		17595: Delta = 69'sb000000000000000000011111111100000000000000000000000000000000000000000;
		14286: Delta = 69'sb111111111111111111011111111100000000000000000000000000000000000000000;
		12799: Delta = 69'sb000000000000000001000000000100000000000000000000000000000000000000000;
		6181: Delta = 69'sb111111111111111111000000000100000000000000000000000000000000000000000;
		44680: Delta = 69'sb000000000000000000111111111100000000000000000000000000000000000000000;
		38062: Delta = 69'sb111111111111111110111111111100000000000000000000000000000000000000000;
		16108: Delta = 69'sb000000000000000010000000000100000000000000000000000000000000000000000;
		2872: Delta = 69'sb111111111111111110000000000100000000000000000000000000000000000000000;
		47989: Delta = 69'sb000000000000000001111111111100000000000000000000000000000000000000000;
		34753: Delta = 69'sb111111111111111101111111111100000000000000000000000000000000000000000;
		22726: Delta = 69'sb000000000000000100000000000100000000000000000000000000000000000000000;
		47115: Delta = 69'sb111111111111111100000000000100000000000000000000000000000000000000000;
		3746: Delta = 69'sb000000000000000011111111111100000000000000000000000000000000000000000;
		28135: Delta = 69'sb111111111111111011111111111100000000000000000000000000000000000000000;
		35962: Delta = 69'sb000000000000001000000000000100000000000000000000000000000000000000000;
		33879: Delta = 69'sb111111111111111000000000000100000000000000000000000000000000000000000;
		16982: Delta = 69'sb000000000000000111111111111100000000000000000000000000000000000000000;
		14899: Delta = 69'sb111111111111110111111111111100000000000000000000000000000000000000000;
		11573: Delta = 69'sb000000000000010000000000000100000000000000000000000000000000000000000;
		7407: Delta = 69'sb111111111111110000000000000100000000000000000000000000000000000000000;
		43454: Delta = 69'sb000000000000001111111111111100000000000000000000000000000000000000000;
		39288: Delta = 69'sb111111111111101111111111111100000000000000000000000000000000000000000;
		13656: Delta = 69'sb000000000000100000000000000100000000000000000000000000000000000000000;
		5324: Delta = 69'sb111111111111100000000000000100000000000000000000000000000000000000000;
		45537: Delta = 69'sb000000000000011111111111111100000000000000000000000000000000000000000;
		37205: Delta = 69'sb111111111111011111111111111100000000000000000000000000000000000000000;
		17822: Delta = 69'sb000000000001000000000000000100000000000000000000000000000000000000000;
		1158: Delta = 69'sb111111111111000000000000000100000000000000000000000000000000000000000;
		49703: Delta = 69'sb000000000000111111111111111100000000000000000000000000000000000000000;
		33039: Delta = 69'sb111111111110111111111111111100000000000000000000000000000000000000000;
		26154: Delta = 69'sb000000000010000000000000000100000000000000000000000000000000000000000;
		43687: Delta = 69'sb111111111110000000000000000100000000000000000000000000000000000000000;
		7174: Delta = 69'sb000000000001111111111111111100000000000000000000000000000000000000000;
		24707: Delta = 69'sb111111111101111111111111111100000000000000000000000000000000000000000;
		42818: Delta = 69'sb000000000100000000000000000100000000000000000000000000000000000000000;
		27023: Delta = 69'sb111111111100000000000000000100000000000000000000000000000000000000000;
		23838: Delta = 69'sb000000000011111111111111111100000000000000000000000000000000000000000;
		8043: Delta = 69'sb111111111011111111111111111100000000000000000000000000000000000000000;
		25285: Delta = 69'sb000000001000000000000000000100000000000000000000000000000000000000000;
		44556: Delta = 69'sb111111111000000000000000000100000000000000000000000000000000000000000;
		6305: Delta = 69'sb000000000111111111111111111100000000000000000000000000000000000000000;
		25576: Delta = 69'sb111111110111111111111111111100000000000000000000000000000000000000000;
		41080: Delta = 69'sb000000010000000000000000000100000000000000000000000000000000000000000;
		28761: Delta = 69'sb111111110000000000000000000100000000000000000000000000000000000000000;
		22100: Delta = 69'sb000000001111111111111111111100000000000000000000000000000000000000000;
		9781: Delta = 69'sb111111101111111111111111111100000000000000000000000000000000000000000;
		21809: Delta = 69'sb000000100000000000000000000100000000000000000000000000000000000000000;
		48032: Delta = 69'sb111111100000000000000000000100000000000000000000000000000000000000000;
		2829: Delta = 69'sb000000011111111111111111111100000000000000000000000000000000000000000;
		29052: Delta = 69'sb111111011111111111111111111100000000000000000000000000000000000000000;
		34128: Delta = 69'sb000001000000000000000000000100000000000000000000000000000000000000000;
		35713: Delta = 69'sb111111000000000000000000000100000000000000000000000000000000000000000;
		15148: Delta = 69'sb000000111111111111111111111100000000000000000000000000000000000000000;
		16733: Delta = 69'sb111110111111111111111111111100000000000000000000000000000000000000000;
		7905: Delta = 69'sb000010000000000000000000000100000000000000000000000000000000000000000;
		11075: Delta = 69'sb111110000000000000000000000100000000000000000000000000000000000000000;
		39786: Delta = 69'sb000001111111111111111111111100000000000000000000000000000000000000000;
		42956: Delta = 69'sb111101111111111111111111111100000000000000000000000000000000000000000;
		6320: Delta = 69'sb000100000000000000000000000100000000000000000000000000000000000000000;
		12660: Delta = 69'sb111100000000000000000000000100000000000000000000000000000000000000000;
		38201: Delta = 69'sb000011111111111111111111111100000000000000000000000000000000000000000;
		44541: Delta = 69'sb111011111111111111111111111100000000000000000000000000000000000000000;
		3150: Delta = 69'sb001000000000000000000000000100000000000000000000000000000000000000000;
		15830: Delta = 69'sb111000000000000000000000000100000000000000000000000000000000000000000;
		35031: Delta = 69'sb000111111111111111111111111100000000000000000000000000000000000000000;
		47711: Delta = 69'sb110111111111111111111111111100000000000000000000000000000000000000000;
		47671: Delta = 69'sb010000000000000000000000000100000000000000000000000000000000000000000;
		22170: Delta = 69'sb110000000000000000000000000100000000000000000000000000000000000000000;
		28691: Delta = 69'sb001111111111111111111111111100000000000000000000000000000000000000000;
		3190: Delta = 69'sb101111111111111111111111111100000000000000000000000000000000000000000;
		6079: Delta = 69'sb000000000000000000000000011000000000000000000000000000000000000000000;
		44782: Delta = 69'sb111111111111111111111111101000000000000000000000000000000000000000000;
		44039: Delta = 69'sb000000000000000000000000101000000000000000000000000000000000000000000;
		6822: Delta = 69'sb111111111111111111111111011000000000000000000000000000000000000000000;
		18237: Delta = 69'sb000000000000000000000001001000000000000000000000000000000000000000000;
		19723: Delta = 69'sb111111111111111111111111001000000000000000000000000000000000000000000;
		31138: Delta = 69'sb000000000000000000000000111000000000000000000000000000000000000000000;
		32624: Delta = 69'sb111111111111111111111110111000000000000000000000000000000000000000000;
		17494: Delta = 69'sb000000000000000000000010001000000000000000000000000000000000000000000;
		20466: Delta = 69'sb111111111111111111111110001000000000000000000000000000000000000000000;
		30395: Delta = 69'sb000000000000000000000001111000000000000000000000000000000000000000000;
		33367: Delta = 69'sb111111111111111111111101111000000000000000000000000000000000000000000;
		16008: Delta = 69'sb000000000000000000000100001000000000000000000000000000000000000000000;
		21952: Delta = 69'sb111111111111111111111100001000000000000000000000000000000000000000000;
		28909: Delta = 69'sb000000000000000000000011111000000000000000000000000000000000000000000;
		34853: Delta = 69'sb111111111111111111111011111000000000000000000000000000000000000000000;
		13036: Delta = 69'sb000000000000000000001000001000000000000000000000000000000000000000000;
		24924: Delta = 69'sb111111111111111111111000001000000000000000000000000000000000000000000;
		25937: Delta = 69'sb000000000000000000000111111000000000000000000000000000000000000000000;
		37825: Delta = 69'sb111111111111111111110111111000000000000000000000000000000000000000000;
		7092: Delta = 69'sb000000000000000000010000001000000000000000000000000000000000000000000;
		30868: Delta = 69'sb111111111111111111110000001000000000000000000000000000000000000000000;
		19993: Delta = 69'sb000000000000000000001111111000000000000000000000000000000000000000000;
		43769: Delta = 69'sb111111111111111111101111111000000000000000000000000000000000000000000;
		46065: Delta = 69'sb000000000000000000100000001000000000000000000000000000000000000000000;
		42756: Delta = 69'sb111111111111111111100000001000000000000000000000000000000000000000000;
		8105: Delta = 69'sb000000000000000000011111111000000000000000000000000000000000000000000;
		4796: Delta = 69'sb111111111111111111011111111000000000000000000000000000000000000000000;
		22289: Delta = 69'sb000000000000000001000000001000000000000000000000000000000000000000000;
		15671: Delta = 69'sb111111111111111111000000001000000000000000000000000000000000000000000;
		35190: Delta = 69'sb000000000000000000111111111000000000000000000000000000000000000000000;
		28572: Delta = 69'sb111111111111111110111111111000000000000000000000000000000000000000000;
		25598: Delta = 69'sb000000000000000010000000001000000000000000000000000000000000000000000;
		12362: Delta = 69'sb111111111111111110000000001000000000000000000000000000000000000000000;
		38499: Delta = 69'sb000000000000000001111111111000000000000000000000000000000000000000000;
		25263: Delta = 69'sb111111111111111101111111111000000000000000000000000000000000000000000;
		32216: Delta = 69'sb000000000000000100000000001000000000000000000000000000000000000000000;
		5744: Delta = 69'sb111111111111111100000000001000000000000000000000000000000000000000000;
		45117: Delta = 69'sb000000000000000011111111111000000000000000000000000000000000000000000;
		18645: Delta = 69'sb111111111111111011111111111000000000000000000000000000000000000000000;
		45452: Delta = 69'sb000000000000001000000000001000000000000000000000000000000000000000000;
		43369: Delta = 69'sb111111111111111000000000001000000000000000000000000000000000000000000;
		7492: Delta = 69'sb000000000000000111111111111000000000000000000000000000000000000000000;
		5409: Delta = 69'sb111111111111110111111111111000000000000000000000000000000000000000000;
		21063: Delta = 69'sb000000000000010000000000001000000000000000000000000000000000000000000;
		16897: Delta = 69'sb111111111111110000000000001000000000000000000000000000000000000000000;
		33964: Delta = 69'sb000000000000001111111111111000000000000000000000000000000000000000000;
		29798: Delta = 69'sb111111111111101111111111111000000000000000000000000000000000000000000;
		23146: Delta = 69'sb000000000000100000000000001000000000000000000000000000000000000000000;
		14814: Delta = 69'sb111111111111100000000000001000000000000000000000000000000000000000000;
		36047: Delta = 69'sb000000000000011111111111111000000000000000000000000000000000000000000;
		27715: Delta = 69'sb111111111111011111111111111000000000000000000000000000000000000000000;
		27312: Delta = 69'sb000000000001000000000000001000000000000000000000000000000000000000000;
		10648: Delta = 69'sb111111111111000000000000001000000000000000000000000000000000000000000;
		40213: Delta = 69'sb000000000000111111111111111000000000000000000000000000000000000000000;
		23549: Delta = 69'sb111111111110111111111111111000000000000000000000000000000000000000000;
		35644: Delta = 69'sb000000000010000000000000001000000000000000000000000000000000000000000;
		2316: Delta = 69'sb111111111110000000000000001000000000000000000000000000000000000000000;
		48545: Delta = 69'sb000000000001111111111111111000000000000000000000000000000000000000000;
		15217: Delta = 69'sb111111111101111111111111111000000000000000000000000000000000000000000;
		1447: Delta = 69'sb000000000100000000000000001000000000000000000000000000000000000000000;
		36513: Delta = 69'sb111111111100000000000000001000000000000000000000000000000000000000000;
		14348: Delta = 69'sb000000000011111111111111111000000000000000000000000000000000000000000;
		49414: Delta = 69'sb111111111011111111111111111000000000000000000000000000000000000000000;
		34775: Delta = 69'sb000000001000000000000000001000000000000000000000000000000000000000000;
		3185: Delta = 69'sb111111111000000000000000001000000000000000000000000000000000000000000;
		47676: Delta = 69'sb000000000111111111111111111000000000000000000000000000000000000000000;
		16086: Delta = 69'sb111111110111111111111111111000000000000000000000000000000000000000000;
		50570: Delta = 69'sb000000010000000000000000001000000000000000000000000000000000000000000;
		38251: Delta = 69'sb111111110000000000000000001000000000000000000000000000000000000000000;
		12610: Delta = 69'sb000000001111111111111111111000000000000000000000000000000000000000000;
		291: Delta = 69'sb111111101111111111111111111000000000000000000000000000000000000000000;
		31299: Delta = 69'sb000000100000000000000000001000000000000000000000000000000000000000000;
		6661: Delta = 69'sb111111100000000000000000001000000000000000000000000000000000000000000;
		44200: Delta = 69'sb000000011111111111111111111000000000000000000000000000000000000000000;
		19562: Delta = 69'sb111111011111111111111111111000000000000000000000000000000000000000000;
		43618: Delta = 69'sb000001000000000000000000001000000000000000000000000000000000000000000;
		45203: Delta = 69'sb111111000000000000000000001000000000000000000000000000000000000000000;
		5658: Delta = 69'sb000000111111111111111111111000000000000000000000000000000000000000000;
		7243: Delta = 69'sb111110111111111111111111111000000000000000000000000000000000000000000;
		17395: Delta = 69'sb000010000000000000000000001000000000000000000000000000000000000000000;
		20565: Delta = 69'sb111110000000000000000000001000000000000000000000000000000000000000000;
		30296: Delta = 69'sb000001111111111111111111111000000000000000000000000000000000000000000;
		33466: Delta = 69'sb111101111111111111111111111000000000000000000000000000000000000000000;
		15810: Delta = 69'sb000100000000000000000000001000000000000000000000000000000000000000000;
		22150: Delta = 69'sb111100000000000000000000001000000000000000000000000000000000000000000;
		28711: Delta = 69'sb000011111111111111111111111000000000000000000000000000000000000000000;
		35051: Delta = 69'sb111011111111111111111111111000000000000000000000000000000000000000000;
		12640: Delta = 69'sb001000000000000000000000001000000000000000000000000000000000000000000;
		25320: Delta = 69'sb111000000000000000000000001000000000000000000000000000000000000000000;
		25541: Delta = 69'sb000111111111111111111111111000000000000000000000000000000000000000000;
		38221: Delta = 69'sb110111111111111111111111111000000000000000000000000000000000000000000;
		6300: Delta = 69'sb010000000000000000000000001000000000000000000000000000000000000000000;
		31660: Delta = 69'sb110000000000000000000000001000000000000000000000000000000000000000000;
		19201: Delta = 69'sb001111111111111111111111111000000000000000000000000000000000000000000;
		44561: Delta = 69'sb101111111111111111111111111000000000000000000000000000000000000000000;
		12158: Delta = 69'sb000000000000000000000000110000000000000000000000000000000000000000000;
		38703: Delta = 69'sb111111111111111111111111010000000000000000000000000000000000000000000;
		37217: Delta = 69'sb000000000000000000000001010000000000000000000000000000000000000000000;
		13644: Delta = 69'sb111111111111111111111110110000000000000000000000000000000000000000000;
		36474: Delta = 69'sb000000000000000000000010010000000000000000000000000000000000000000000;
		39446: Delta = 69'sb111111111111111111111110010000000000000000000000000000000000000000000;
		11415: Delta = 69'sb000000000000000000000001110000000000000000000000000000000000000000000;
		14387: Delta = 69'sb111111111111111111111101110000000000000000000000000000000000000000000;
		34988: Delta = 69'sb000000000000000000000100010000000000000000000000000000000000000000000;
		40932: Delta = 69'sb111111111111111111111100010000000000000000000000000000000000000000000;
		9929: Delta = 69'sb000000000000000000000011110000000000000000000000000000000000000000000;
		15873: Delta = 69'sb111111111111111111111011110000000000000000000000000000000000000000000;
		32016: Delta = 69'sb000000000000000000001000010000000000000000000000000000000000000000000;
		43904: Delta = 69'sb111111111111111111111000010000000000000000000000000000000000000000000;
		6957: Delta = 69'sb000000000000000000000111110000000000000000000000000000000000000000000;
		18845: Delta = 69'sb111111111111111111110111110000000000000000000000000000000000000000000;
		26072: Delta = 69'sb000000000000000000010000010000000000000000000000000000000000000000000;
		49848: Delta = 69'sb111111111111111111110000010000000000000000000000000000000000000000000;
		1013: Delta = 69'sb000000000000000000001111110000000000000000000000000000000000000000000;
		24789: Delta = 69'sb111111111111111111101111110000000000000000000000000000000000000000000;
		14184: Delta = 69'sb000000000000000000100000010000000000000000000000000000000000000000000;
		10875: Delta = 69'sb111111111111111111100000010000000000000000000000000000000000000000000;
		39986: Delta = 69'sb000000000000000000011111110000000000000000000000000000000000000000000;
		36677: Delta = 69'sb111111111111111111011111110000000000000000000000000000000000000000000;
		41269: Delta = 69'sb000000000000000001000000010000000000000000000000000000000000000000000;
		34651: Delta = 69'sb111111111111111111000000010000000000000000000000000000000000000000000;
		16210: Delta = 69'sb000000000000000000111111110000000000000000000000000000000000000000000;
		9592: Delta = 69'sb111111111111111110111111110000000000000000000000000000000000000000000;
		44578: Delta = 69'sb000000000000000010000000010000000000000000000000000000000000000000000;
		31342: Delta = 69'sb111111111111111110000000010000000000000000000000000000000000000000000;
		19519: Delta = 69'sb000000000000000001111111110000000000000000000000000000000000000000000;
		6283: Delta = 69'sb111111111111111101111111110000000000000000000000000000000000000000000;
		335: Delta = 69'sb000000000000000100000000010000000000000000000000000000000000000000000;
		24724: Delta = 69'sb111111111111111100000000010000000000000000000000000000000000000000000;
		26137: Delta = 69'sb000000000000000011111111110000000000000000000000000000000000000000000;
		50526: Delta = 69'sb111111111111111011111111110000000000000000000000000000000000000000000;
		13571: Delta = 69'sb000000000000001000000000010000000000000000000000000000000000000000000;
		11488: Delta = 69'sb111111111111111000000000010000000000000000000000000000000000000000000;
		39373: Delta = 69'sb000000000000000111111111110000000000000000000000000000000000000000000;
		37290: Delta = 69'sb111111111111110111111111110000000000000000000000000000000000000000000;
		40043: Delta = 69'sb000000000000010000000000010000000000000000000000000000000000000000000;
		35877: Delta = 69'sb111111111111110000000000010000000000000000000000000000000000000000000;
		14984: Delta = 69'sb000000000000001111111111110000000000000000000000000000000000000000000;
		10818: Delta = 69'sb111111111111101111111111110000000000000000000000000000000000000000000;
		42126: Delta = 69'sb000000000000100000000000010000000000000000000000000000000000000000000;
		33794: Delta = 69'sb111111111111100000000000010000000000000000000000000000000000000000000;
		17067: Delta = 69'sb000000000000011111111111110000000000000000000000000000000000000000000;
		8735: Delta = 69'sb111111111111011111111111110000000000000000000000000000000000000000000;
		46292: Delta = 69'sb000000000001000000000000010000000000000000000000000000000000000000000;
		29628: Delta = 69'sb111111111111000000000000010000000000000000000000000000000000000000000;
		21233: Delta = 69'sb000000000000111111111111110000000000000000000000000000000000000000000;
		4569: Delta = 69'sb111111111110111111111111110000000000000000000000000000000000000000000;
		3763: Delta = 69'sb000000000010000000000000010000000000000000000000000000000000000000000;
		21296: Delta = 69'sb111111111110000000000000010000000000000000000000000000000000000000000;
		29565: Delta = 69'sb000000000001111111111111110000000000000000000000000000000000000000000;
		47098: Delta = 69'sb111111111101111111111111110000000000000000000000000000000000000000000;
		20427: Delta = 69'sb000000000100000000000000010000000000000000000000000000000000000000000;
		4632: Delta = 69'sb111111111100000000000000010000000000000000000000000000000000000000000;
		46229: Delta = 69'sb000000000011111111111111110000000000000000000000000000000000000000000;
		30434: Delta = 69'sb111111111011111111111111110000000000000000000000000000000000000000000;
		2894: Delta = 69'sb000000001000000000000000010000000000000000000000000000000000000000000;
		22165: Delta = 69'sb111111111000000000000000010000000000000000000000000000000000000000000;
		28696: Delta = 69'sb000000000111111111111111110000000000000000000000000000000000000000000;
		47967: Delta = 69'sb111111110111111111111111110000000000000000000000000000000000000000000;
		18689: Delta = 69'sb000000010000000000000000010000000000000000000000000000000000000000000;
		6370: Delta = 69'sb111111110000000000000000010000000000000000000000000000000000000000000;
		44491: Delta = 69'sb000000001111111111111111110000000000000000000000000000000000000000000;
		32172: Delta = 69'sb111111101111111111111111110000000000000000000000000000000000000000000;
		50279: Delta = 69'sb000000100000000000000000010000000000000000000000000000000000000000000;
		25641: Delta = 69'sb111111100000000000000000010000000000000000000000000000000000000000000;
		25220: Delta = 69'sb000000011111111111111111110000000000000000000000000000000000000000000;
		582: Delta = 69'sb111111011111111111111111110000000000000000000000000000000000000000000;
		11737: Delta = 69'sb000001000000000000000000010000000000000000000000000000000000000000000;
		13322: Delta = 69'sb111111000000000000000000010000000000000000000000000000000000000000000;
		37539: Delta = 69'sb000000111111111111111111110000000000000000000000000000000000000000000;
		39124: Delta = 69'sb111110111111111111111111110000000000000000000000000000000000000000000;
		36375: Delta = 69'sb000010000000000000000000010000000000000000000000000000000000000000000;
		39545: Delta = 69'sb111110000000000000000000010000000000000000000000000000000000000000000;
		11316: Delta = 69'sb000001111111111111111111110000000000000000000000000000000000000000000;
		14486: Delta = 69'sb111101111111111111111111110000000000000000000000000000000000000000000;
		34790: Delta = 69'sb000100000000000000000000010000000000000000000000000000000000000000000;
		41130: Delta = 69'sb111100000000000000000000010000000000000000000000000000000000000000000;
		9731: Delta = 69'sb000011111111111111111111110000000000000000000000000000000000000000000;
		16071: Delta = 69'sb111011111111111111111111110000000000000000000000000000000000000000000;
		31620: Delta = 69'sb001000000000000000000000010000000000000000000000000000000000000000000;
		44300: Delta = 69'sb111000000000000000000000010000000000000000000000000000000000000000000;
		6561: Delta = 69'sb000111111111111111111111110000000000000000000000000000000000000000000;
		19241: Delta = 69'sb110111111111111111111111110000000000000000000000000000000000000000000;
		25280: Delta = 69'sb010000000000000000000000010000000000000000000000000000000000000000000;
		50640: Delta = 69'sb110000000000000000000000010000000000000000000000000000000000000000000;
		221: Delta = 69'sb001111111111111111111111110000000000000000000000000000000000000000000;
		25581: Delta = 69'sb101111111111111111111111110000000000000000000000000000000000000000000;
		24316: Delta = 69'sb000000000000000000000001100000000000000000000000000000000000000000000;
		26545: Delta = 69'sb111111111111111111111110100000000000000000000000000000000000000000000;
		23573: Delta = 69'sb000000000000000000000010100000000000000000000000000000000000000000000;
		27288: Delta = 69'sb111111111111111111111101100000000000000000000000000000000000000000000;
		22087: Delta = 69'sb000000000000000000000100100000000000000000000000000000000000000000000;
		28031: Delta = 69'sb111111111111111111111100100000000000000000000000000000000000000000000;
		22830: Delta = 69'sb000000000000000000000011100000000000000000000000000000000000000000000;
		28774: Delta = 69'sb111111111111111111111011100000000000000000000000000000000000000000000;
		19115: Delta = 69'sb000000000000000000001000100000000000000000000000000000000000000000000;
		31003: Delta = 69'sb111111111111111111111000100000000000000000000000000000000000000000000;
		19858: Delta = 69'sb000000000000000000000111100000000000000000000000000000000000000000000;
		31746: Delta = 69'sb111111111111111111110111100000000000000000000000000000000000000000000;
		13171: Delta = 69'sb000000000000000000010000100000000000000000000000000000000000000000000;
		36947: Delta = 69'sb111111111111111111110000100000000000000000000000000000000000000000000;
		13914: Delta = 69'sb000000000000000000001111100000000000000000000000000000000000000000000;
		37690: Delta = 69'sb111111111111111111101111100000000000000000000000000000000000000000000;
		1283: Delta = 69'sb000000000000000000100000100000000000000000000000000000000000000000000;
		48835: Delta = 69'sb111111111111111111100000100000000000000000000000000000000000000000000;
		2026: Delta = 69'sb000000000000000000011111100000000000000000000000000000000000000000000;
		49578: Delta = 69'sb111111111111111111011111100000000000000000000000000000000000000000000;
		28368: Delta = 69'sb000000000000000001000000100000000000000000000000000000000000000000000;
		21750: Delta = 69'sb111111111111111111000000100000000000000000000000000000000000000000000;
		29111: Delta = 69'sb000000000000000000111111100000000000000000000000000000000000000000000;
		22493: Delta = 69'sb111111111111111110111111100000000000000000000000000000000000000000000;
		31677: Delta = 69'sb000000000000000010000000100000000000000000000000000000000000000000000;
		18441: Delta = 69'sb111111111111111110000000100000000000000000000000000000000000000000000;
		32420: Delta = 69'sb000000000000000001111111100000000000000000000000000000000000000000000;
		19184: Delta = 69'sb111111111111111101111111100000000000000000000000000000000000000000000;
		38295: Delta = 69'sb000000000000000100000000100000000000000000000000000000000000000000000;
		11823: Delta = 69'sb111111111111111100000000100000000000000000000000000000000000000000000;
		39038: Delta = 69'sb000000000000000011111111100000000000000000000000000000000000000000000;
		12566: Delta = 69'sb111111111111111011111111100000000000000000000000000000000000000000000;
		670: Delta = 69'sb000000000000001000000000100000000000000000000000000000000000000000000;
		49448: Delta = 69'sb111111111111111000000000100000000000000000000000000000000000000000000;
		1413: Delta = 69'sb000000000000000111111111100000000000000000000000000000000000000000000;
		50191: Delta = 69'sb111111111111110111111111100000000000000000000000000000000000000000000;
		27142: Delta = 69'sb000000000000010000000000100000000000000000000000000000000000000000000;
		22976: Delta = 69'sb111111111111110000000000100000000000000000000000000000000000000000000;
		27885: Delta = 69'sb000000000000001111111111100000000000000000000000000000000000000000000;
		23719: Delta = 69'sb111111111111101111111111100000000000000000000000000000000000000000000;
		29225: Delta = 69'sb000000000000100000000000100000000000000000000000000000000000000000000;
		20893: Delta = 69'sb111111111111100000000000100000000000000000000000000000000000000000000;
		29968: Delta = 69'sb000000000000011111111111100000000000000000000000000000000000000000000;
		21636: Delta = 69'sb111111111111011111111111100000000000000000000000000000000000000000000;
		33391: Delta = 69'sb000000000001000000000000100000000000000000000000000000000000000000000;
		16727: Delta = 69'sb111111111111000000000000100000000000000000000000000000000000000000000;
		34134: Delta = 69'sb000000000000111111111111100000000000000000000000000000000000000000000;
		17470: Delta = 69'sb111111111110111111111111100000000000000000000000000000000000000000000;
		41723: Delta = 69'sb000000000010000000000000100000000000000000000000000000000000000000000;
		8395: Delta = 69'sb111111111110000000000000100000000000000000000000000000000000000000000;
		42466: Delta = 69'sb000000000001111111111111100000000000000000000000000000000000000000000;
		9138: Delta = 69'sb111111111101111111111111100000000000000000000000000000000000000000000;
		7526: Delta = 69'sb000000000100000000000000100000000000000000000000000000000000000000000;
		42592: Delta = 69'sb111111111100000000000000100000000000000000000000000000000000000000000;
		8269: Delta = 69'sb000000000011111111111111100000000000000000000000000000000000000000000;
		43335: Delta = 69'sb111111111011111111111111100000000000000000000000000000000000000000000;
		40854: Delta = 69'sb000000001000000000000000100000000000000000000000000000000000000000000;
		9264: Delta = 69'sb111111111000000000000000100000000000000000000000000000000000000000000;
		41597: Delta = 69'sb000000000111111111111111100000000000000000000000000000000000000000000;
		10007: Delta = 69'sb111111110111111111111111100000000000000000000000000000000000000000000;
		5788: Delta = 69'sb000000010000000000000000100000000000000000000000000000000000000000000;
		44330: Delta = 69'sb111111110000000000000000100000000000000000000000000000000000000000000;
		6531: Delta = 69'sb000000001111111111111111100000000000000000000000000000000000000000000;
		45073: Delta = 69'sb111111101111111111111111100000000000000000000000000000000000000000000;
		37378: Delta = 69'sb000000100000000000000000100000000000000000000000000000000000000000000;
		12740: Delta = 69'sb111111100000000000000000100000000000000000000000000000000000000000000;
		38121: Delta = 69'sb000000011111111111111111100000000000000000000000000000000000000000000;
		13483: Delta = 69'sb111111011111111111111111100000000000000000000000000000000000000000000;
		49697: Delta = 69'sb000001000000000000000000100000000000000000000000000000000000000000000;
		421: Delta = 69'sb111111000000000000000000100000000000000000000000000000000000000000000;
		50440: Delta = 69'sb000000111111111111111111100000000000000000000000000000000000000000000;
		1164: Delta = 69'sb111110111111111111111111100000000000000000000000000000000000000000000;
		23474: Delta = 69'sb000010000000000000000000100000000000000000000000000000000000000000000;
		26644: Delta = 69'sb111110000000000000000000100000000000000000000000000000000000000000000;
		24217: Delta = 69'sb000001111111111111111111100000000000000000000000000000000000000000000;
		27387: Delta = 69'sb111101111111111111111111100000000000000000000000000000000000000000000;
		21889: Delta = 69'sb000100000000000000000000100000000000000000000000000000000000000000000;
		28229: Delta = 69'sb111100000000000000000000100000000000000000000000000000000000000000000;
		22632: Delta = 69'sb000011111111111111111111100000000000000000000000000000000000000000000;
		28972: Delta = 69'sb111011111111111111111111100000000000000000000000000000000000000000000;
		18719: Delta = 69'sb001000000000000000000000100000000000000000000000000000000000000000000;
		31399: Delta = 69'sb111000000000000000000000100000000000000000000000000000000000000000000;
		19462: Delta = 69'sb000111111111111111111111100000000000000000000000000000000000000000000;
		32142: Delta = 69'sb110111111111111111111111100000000000000000000000000000000000000000000;
		12379: Delta = 69'sb010000000000000000000000100000000000000000000000000000000000000000000;
		37739: Delta = 69'sb110000000000000000000000100000000000000000000000000000000000000000000;
		13122: Delta = 69'sb001111111111111111111111100000000000000000000000000000000000000000000;
		38482: Delta = 69'sb101111111111111111111111100000000000000000000000000000000000000000000;
		48632: Delta = 69'sb000000000000000000000011000000000000000000000000000000000000000000000;
		2229: Delta = 69'sb111111111111111111111101000000000000000000000000000000000000000000000;
		47146: Delta = 69'sb000000000000000000000101000000000000000000000000000000000000000000000;
		3715: Delta = 69'sb111111111111111111111011000000000000000000000000000000000000000000000;
		44174: Delta = 69'sb000000000000000000001001000000000000000000000000000000000000000000000;
		5201: Delta = 69'sb111111111111111111111001000000000000000000000000000000000000000000000;
		45660: Delta = 69'sb000000000000000000000111000000000000000000000000000000000000000000000;
		6687: Delta = 69'sb111111111111111111110111000000000000000000000000000000000000000000000;
		38230: Delta = 69'sb000000000000000000010001000000000000000000000000000000000000000000000;
		11145: Delta = 69'sb111111111111111111110001000000000000000000000000000000000000000000000;
		39716: Delta = 69'sb000000000000000000001111000000000000000000000000000000000000000000000;
		12631: Delta = 69'sb111111111111111111101111000000000000000000000000000000000000000000000;
		26342: Delta = 69'sb000000000000000000100001000000000000000000000000000000000000000000000;
		23033: Delta = 69'sb111111111111111111100001000000000000000000000000000000000000000000000;
		27828: Delta = 69'sb000000000000000000011111000000000000000000000000000000000000000000000;
		24519: Delta = 69'sb111111111111111111011111000000000000000000000000000000000000000000000;
		2566: Delta = 69'sb000000000000000001000001000000000000000000000000000000000000000000000;
		46809: Delta = 69'sb111111111111111111000001000000000000000000000000000000000000000000000;
		4052: Delta = 69'sb000000000000000000111111000000000000000000000000000000000000000000000;
		48295: Delta = 69'sb111111111111111110111111000000000000000000000000000000000000000000000;
		5875: Delta = 69'sb000000000000000010000001000000000000000000000000000000000000000000000;
		43500: Delta = 69'sb111111111111111110000001000000000000000000000000000000000000000000000;
		7361: Delta = 69'sb000000000000000001111111000000000000000000000000000000000000000000000;
		44986: Delta = 69'sb111111111111111101111111000000000000000000000000000000000000000000000;
		12493: Delta = 69'sb000000000000000100000001000000000000000000000000000000000000000000000;
		36882: Delta = 69'sb111111111111111100000001000000000000000000000000000000000000000000000;
		13979: Delta = 69'sb000000000000000011111111000000000000000000000000000000000000000000000;
		38368: Delta = 69'sb111111111111111011111111000000000000000000000000000000000000000000000;
		25729: Delta = 69'sb000000000000001000000001000000000000000000000000000000000000000000000;
		23646: Delta = 69'sb111111111111111000000001000000000000000000000000000000000000000000000;
		27215: Delta = 69'sb000000000000000111111111000000000000000000000000000000000000000000000;
		25132: Delta = 69'sb111111111111110111111111000000000000000000000000000000000000000000000;
		1340: Delta = 69'sb000000000000010000000001000000000000000000000000000000000000000000000;
		48035: Delta = 69'sb111111111111110000000001000000000000000000000000000000000000000000000;
		2826: Delta = 69'sb000000000000001111111111000000000000000000000000000000000000000000000;
		49521: Delta = 69'sb111111111111101111111111000000000000000000000000000000000000000000000;
		3423: Delta = 69'sb000000000000100000000001000000000000000000000000000000000000000000000;
		45952: Delta = 69'sb111111111111100000000001000000000000000000000000000000000000000000000;
		4909: Delta = 69'sb000000000000011111111111000000000000000000000000000000000000000000000;
		47438: Delta = 69'sb111111111111011111111111000000000000000000000000000000000000000000000;
		7589: Delta = 69'sb000000000001000000000001000000000000000000000000000000000000000000000;
		41786: Delta = 69'sb111111111111000000000001000000000000000000000000000000000000000000000;
		9075: Delta = 69'sb000000000000111111111111000000000000000000000000000000000000000000000;
		43272: Delta = 69'sb111111111110111111111111000000000000000000000000000000000000000000000;
		15921: Delta = 69'sb000000000010000000000001000000000000000000000000000000000000000000000;
		33454: Delta = 69'sb111111111110000000000001000000000000000000000000000000000000000000000;
		17407: Delta = 69'sb000000000001111111111111000000000000000000000000000000000000000000000;
		34940: Delta = 69'sb111111111101111111111111000000000000000000000000000000000000000000000;
		32585: Delta = 69'sb000000000100000000000001000000000000000000000000000000000000000000000;
		16790: Delta = 69'sb111111111100000000000001000000000000000000000000000000000000000000000;
		34071: Delta = 69'sb000000000011111111111111000000000000000000000000000000000000000000000;
		18276: Delta = 69'sb111111111011111111111111000000000000000000000000000000000000000000000;
		15052: Delta = 69'sb000000001000000000000001000000000000000000000000000000000000000000000;
		34323: Delta = 69'sb111111111000000000000001000000000000000000000000000000000000000000000;
		16538: Delta = 69'sb000000000111111111111111000000000000000000000000000000000000000000000;
		35809: Delta = 69'sb111111110111111111111111000000000000000000000000000000000000000000000;
		30847: Delta = 69'sb000000010000000000000001000000000000000000000000000000000000000000000;
		18528: Delta = 69'sb111111110000000000000001000000000000000000000000000000000000000000000;
		32333: Delta = 69'sb000000001111111111111111000000000000000000000000000000000000000000000;
		20014: Delta = 69'sb111111101111111111111111000000000000000000000000000000000000000000000;
		11576: Delta = 69'sb000000100000000000000001000000000000000000000000000000000000000000000;
		37799: Delta = 69'sb111111100000000000000001000000000000000000000000000000000000000000000;
		13062: Delta = 69'sb000000011111111111111111000000000000000000000000000000000000000000000;
		39285: Delta = 69'sb111111011111111111111111000000000000000000000000000000000000000000000;
		23895: Delta = 69'sb000001000000000000000001000000000000000000000000000000000000000000000;
		25480: Delta = 69'sb111111000000000000000001000000000000000000000000000000000000000000000;
		25381: Delta = 69'sb000000111111111111111111000000000000000000000000000000000000000000000;
		26966: Delta = 69'sb111110111111111111111111000000000000000000000000000000000000000000000;
		48533: Delta = 69'sb000010000000000000000001000000000000000000000000000000000000000000000;
		842: Delta = 69'sb111110000000000000000001000000000000000000000000000000000000000000000;
		50019: Delta = 69'sb000001111111111111111111000000000000000000000000000000000000000000000;
		2328: Delta = 69'sb111101111111111111111111000000000000000000000000000000000000000000000;
		46948: Delta = 69'sb000100000000000000000001000000000000000000000000000000000000000000000;
		2427: Delta = 69'sb111100000000000000000001000000000000000000000000000000000000000000000;
		48434: Delta = 69'sb000011111111111111111111000000000000000000000000000000000000000000000;
		3913: Delta = 69'sb111011111111111111111111000000000000000000000000000000000000000000000;
		43778: Delta = 69'sb001000000000000000000001000000000000000000000000000000000000000000000;
		5597: Delta = 69'sb111000000000000000000001000000000000000000000000000000000000000000000;
		45264: Delta = 69'sb000111111111111111111111000000000000000000000000000000000000000000000;
		7083: Delta = 69'sb110111111111111111111111000000000000000000000000000000000000000000000;
		37438: Delta = 69'sb010000000000000000000001000000000000000000000000000000000000000000000;
		11937: Delta = 69'sb110000000000000000000001000000000000000000000000000000000000000000000;
		38924: Delta = 69'sb001111111111111111111111000000000000000000000000000000000000000000000;
		13423: Delta = 69'sb101111111111111111111111000000000000000000000000000000000000000000000;
		46403: Delta = 69'sb000000000000000000000110000000000000000000000000000000000000000000000;
		4458: Delta = 69'sb111111111111111111111010000000000000000000000000000000000000000000000;
		43431: Delta = 69'sb000000000000000000001010000000000000000000000000000000000000000000000;
		7430: Delta = 69'sb111111111111111111110110000000000000000000000000000000000000000000000;
		37487: Delta = 69'sb000000000000000000010010000000000000000000000000000000000000000000000;
		10402: Delta = 69'sb111111111111111111110010000000000000000000000000000000000000000000000;
		40459: Delta = 69'sb000000000000000000001110000000000000000000000000000000000000000000000;
		13374: Delta = 69'sb111111111111111111101110000000000000000000000000000000000000000000000;
		25599: Delta = 69'sb000000000000000000100010000000000000000000000000000000000000000000000;
		22290: Delta = 69'sb111111111111111111100010000000000000000000000000000000000000000000000;
		28571: Delta = 69'sb000000000000000000011110000000000000000000000000000000000000000000000;
		25262: Delta = 69'sb111111111111111111011110000000000000000000000000000000000000000000000;
		1823: Delta = 69'sb000000000000000001000010000000000000000000000000000000000000000000000;
		46066: Delta = 69'sb111111111111111111000010000000000000000000000000000000000000000000000;
		4795: Delta = 69'sb000000000000000000111110000000000000000000000000000000000000000000000;
		49038: Delta = 69'sb111111111111111110111110000000000000000000000000000000000000000000000;
		5132: Delta = 69'sb000000000000000010000010000000000000000000000000000000000000000000000;
		42757: Delta = 69'sb111111111111111110000010000000000000000000000000000000000000000000000;
		8104: Delta = 69'sb000000000000000001111110000000000000000000000000000000000000000000000;
		45729: Delta = 69'sb111111111111111101111110000000000000000000000000000000000000000000000;
		11750: Delta = 69'sb000000000000000100000010000000000000000000000000000000000000000000000;
		36139: Delta = 69'sb111111111111111100000010000000000000000000000000000000000000000000000;
		14722: Delta = 69'sb000000000000000011111110000000000000000000000000000000000000000000000;
		39111: Delta = 69'sb111111111111111011111110000000000000000000000000000000000000000000000;
		24986: Delta = 69'sb000000000000001000000010000000000000000000000000000000000000000000000;
		22903: Delta = 69'sb111111111111111000000010000000000000000000000000000000000000000000000;
		27958: Delta = 69'sb000000000000000111111110000000000000000000000000000000000000000000000;
		25875: Delta = 69'sb111111111111110111111110000000000000000000000000000000000000000000000;
		597: Delta = 69'sb000000000000010000000010000000000000000000000000000000000000000000000;
		47292: Delta = 69'sb111111111111110000000010000000000000000000000000000000000000000000000;
		3569: Delta = 69'sb000000000000001111111110000000000000000000000000000000000000000000000;
		50264: Delta = 69'sb111111111111101111111110000000000000000000000000000000000000000000000;
		2680: Delta = 69'sb000000000000100000000010000000000000000000000000000000000000000000000;
		45209: Delta = 69'sb111111111111100000000010000000000000000000000000000000000000000000000;
		5652: Delta = 69'sb000000000000011111111110000000000000000000000000000000000000000000000;
		48181: Delta = 69'sb111111111111011111111110000000000000000000000000000000000000000000000;
		6846: Delta = 69'sb000000000001000000000010000000000000000000000000000000000000000000000;
		41043: Delta = 69'sb111111111111000000000010000000000000000000000000000000000000000000000;
		9818: Delta = 69'sb000000000000111111111110000000000000000000000000000000000000000000000;
		44015: Delta = 69'sb111111111110111111111110000000000000000000000000000000000000000000000;
		15178: Delta = 69'sb000000000010000000000010000000000000000000000000000000000000000000000;
		32711: Delta = 69'sb111111111110000000000010000000000000000000000000000000000000000000000;
		18150: Delta = 69'sb000000000001111111111110000000000000000000000000000000000000000000000;
		35683: Delta = 69'sb111111111101111111111110000000000000000000000000000000000000000000000;
		31842: Delta = 69'sb000000000100000000000010000000000000000000000000000000000000000000000;
		16047: Delta = 69'sb111111111100000000000010000000000000000000000000000000000000000000000;
		34814: Delta = 69'sb000000000011111111111110000000000000000000000000000000000000000000000;
		19019: Delta = 69'sb111111111011111111111110000000000000000000000000000000000000000000000;
		14309: Delta = 69'sb000000001000000000000010000000000000000000000000000000000000000000000;
		33580: Delta = 69'sb111111111000000000000010000000000000000000000000000000000000000000000;
		17281: Delta = 69'sb000000000111111111111110000000000000000000000000000000000000000000000;
		36552: Delta = 69'sb111111110111111111111110000000000000000000000000000000000000000000000;
		30104: Delta = 69'sb000000010000000000000010000000000000000000000000000000000000000000000;
		17785: Delta = 69'sb111111110000000000000010000000000000000000000000000000000000000000000;
		33076: Delta = 69'sb000000001111111111111110000000000000000000000000000000000000000000000;
		20757: Delta = 69'sb111111101111111111111110000000000000000000000000000000000000000000000;
		10833: Delta = 69'sb000000100000000000000010000000000000000000000000000000000000000000000;
		37056: Delta = 69'sb111111100000000000000010000000000000000000000000000000000000000000000;
		13805: Delta = 69'sb000000011111111111111110000000000000000000000000000000000000000000000;
		40028: Delta = 69'sb111111011111111111111110000000000000000000000000000000000000000000000;
		23152: Delta = 69'sb000001000000000000000010000000000000000000000000000000000000000000000;
		24737: Delta = 69'sb111111000000000000000010000000000000000000000000000000000000000000000;
		26124: Delta = 69'sb000000111111111111111110000000000000000000000000000000000000000000000;
		27709: Delta = 69'sb111110111111111111111110000000000000000000000000000000000000000000000;
		47790: Delta = 69'sb000010000000000000000010000000000000000000000000000000000000000000000;
		99: Delta = 69'sb111110000000000000000010000000000000000000000000000000000000000000000;
		50762: Delta = 69'sb000001111111111111111110000000000000000000000000000000000000000000000;
		3071: Delta = 69'sb111101111111111111111110000000000000000000000000000000000000000000000;
		46205: Delta = 69'sb000100000000000000000010000000000000000000000000000000000000000000000;
		1684: Delta = 69'sb111100000000000000000010000000000000000000000000000000000000000000000;
		49177: Delta = 69'sb000011111111111111111110000000000000000000000000000000000000000000000;
		4656: Delta = 69'sb111011111111111111111110000000000000000000000000000000000000000000000;
		43035: Delta = 69'sb001000000000000000000010000000000000000000000000000000000000000000000;
		4854: Delta = 69'sb111000000000000000000010000000000000000000000000000000000000000000000;
		46007: Delta = 69'sb000111111111111111111110000000000000000000000000000000000000000000000;
		7826: Delta = 69'sb110111111111111111111110000000000000000000000000000000000000000000000;
		36695: Delta = 69'sb010000000000000000000010000000000000000000000000000000000000000000000;
		11194: Delta = 69'sb110000000000000000000010000000000000000000000000000000000000000000000;
		39667: Delta = 69'sb001111111111111111111110000000000000000000000000000000000000000000000;
		14166: Delta = 69'sb101111111111111111111110000000000000000000000000000000000000000000000;
		41945: Delta = 69'sb000000000000000000001100000000000000000000000000000000000000000000000;
		8916: Delta = 69'sb111111111111111111110100000000000000000000000000000000000000000000000;
		36001: Delta = 69'sb000000000000000000010100000000000000000000000000000000000000000000000;
		14860: Delta = 69'sb111111111111111111101100000000000000000000000000000000000000000000000;
		24113: Delta = 69'sb000000000000000000100100000000000000000000000000000000000000000000000;
		20804: Delta = 69'sb111111111111111111100100000000000000000000000000000000000000000000000;
		30057: Delta = 69'sb000000000000000000011100000000000000000000000000000000000000000000000;
		26748: Delta = 69'sb111111111111111111011100000000000000000000000000000000000000000000000;
		337: Delta = 69'sb000000000000000001000100000000000000000000000000000000000000000000000;
		44580: Delta = 69'sb111111111111111111000100000000000000000000000000000000000000000000000;
		6281: Delta = 69'sb000000000000000000111100000000000000000000000000000000000000000000000;
		50524: Delta = 69'sb111111111111111110111100000000000000000000000000000000000000000000000;
		3646: Delta = 69'sb000000000000000010000100000000000000000000000000000000000000000000000;
		41271: Delta = 69'sb111111111111111110000100000000000000000000000000000000000000000000000;
		9590: Delta = 69'sb000000000000000001111100000000000000000000000000000000000000000000000;
		47215: Delta = 69'sb111111111111111101111100000000000000000000000000000000000000000000000;
		10264: Delta = 69'sb000000000000000100000100000000000000000000000000000000000000000000000;
		34653: Delta = 69'sb111111111111111100000100000000000000000000000000000000000000000000000;
		16208: Delta = 69'sb000000000000000011111100000000000000000000000000000000000000000000000;
		40597: Delta = 69'sb111111111111111011111100000000000000000000000000000000000000000000000;
		23500: Delta = 69'sb000000000000001000000100000000000000000000000000000000000000000000000;
		21417: Delta = 69'sb111111111111111000000100000000000000000000000000000000000000000000000;
		29444: Delta = 69'sb000000000000000111111100000000000000000000000000000000000000000000000;
		27361: Delta = 69'sb111111111111110111111100000000000000000000000000000000000000000000000;
		49972: Delta = 69'sb000000000000010000000100000000000000000000000000000000000000000000000;
		45806: Delta = 69'sb111111111111110000000100000000000000000000000000000000000000000000000;
		5055: Delta = 69'sb000000000000001111111100000000000000000000000000000000000000000000000;
		889: Delta = 69'sb111111111111101111111100000000000000000000000000000000000000000000000;
		1194: Delta = 69'sb000000000000100000000100000000000000000000000000000000000000000000000;
		43723: Delta = 69'sb111111111111100000000100000000000000000000000000000000000000000000000;
		7138: Delta = 69'sb000000000000011111111100000000000000000000000000000000000000000000000;
		49667: Delta = 69'sb111111111111011111111100000000000000000000000000000000000000000000000;
		5360: Delta = 69'sb000000000001000000000100000000000000000000000000000000000000000000000;
		39557: Delta = 69'sb111111111111000000000100000000000000000000000000000000000000000000000;
		11304: Delta = 69'sb000000000000111111111100000000000000000000000000000000000000000000000;
		45501: Delta = 69'sb111111111110111111111100000000000000000000000000000000000000000000000;
		13692: Delta = 69'sb000000000010000000000100000000000000000000000000000000000000000000000;
		31225: Delta = 69'sb111111111110000000000100000000000000000000000000000000000000000000000;
		19636: Delta = 69'sb000000000001111111111100000000000000000000000000000000000000000000000;
		37169: Delta = 69'sb111111111101111111111100000000000000000000000000000000000000000000000;
		30356: Delta = 69'sb000000000100000000000100000000000000000000000000000000000000000000000;
		14561: Delta = 69'sb111111111100000000000100000000000000000000000000000000000000000000000;
		36300: Delta = 69'sb000000000011111111111100000000000000000000000000000000000000000000000;
		20505: Delta = 69'sb111111111011111111111100000000000000000000000000000000000000000000000;
		12823: Delta = 69'sb000000001000000000000100000000000000000000000000000000000000000000000;
		32094: Delta = 69'sb111111111000000000000100000000000000000000000000000000000000000000000;
		18767: Delta = 69'sb000000000111111111111100000000000000000000000000000000000000000000000;
		38038: Delta = 69'sb111111110111111111111100000000000000000000000000000000000000000000000;
		28618: Delta = 69'sb000000010000000000000100000000000000000000000000000000000000000000000;
		16299: Delta = 69'sb111111110000000000000100000000000000000000000000000000000000000000000;
		34562: Delta = 69'sb000000001111111111111100000000000000000000000000000000000000000000000;
		22243: Delta = 69'sb111111101111111111111100000000000000000000000000000000000000000000000;
		9347: Delta = 69'sb000000100000000000000100000000000000000000000000000000000000000000000;
		35570: Delta = 69'sb111111100000000000000100000000000000000000000000000000000000000000000;
		15291: Delta = 69'sb000000011111111111111100000000000000000000000000000000000000000000000;
		41514: Delta = 69'sb111111011111111111111100000000000000000000000000000000000000000000000;
		21666: Delta = 69'sb000001000000000000000100000000000000000000000000000000000000000000000;
		23251: Delta = 69'sb111111000000000000000100000000000000000000000000000000000000000000000;
		27610: Delta = 69'sb000000111111111111111100000000000000000000000000000000000000000000000;
		29195: Delta = 69'sb111110111111111111111100000000000000000000000000000000000000000000000;
		46304: Delta = 69'sb000010000000000000000100000000000000000000000000000000000000000000000;
		49474: Delta = 69'sb111110000000000000000100000000000000000000000000000000000000000000000;
		1387: Delta = 69'sb000001111111111111111100000000000000000000000000000000000000000000000;
		4557: Delta = 69'sb111101111111111111111100000000000000000000000000000000000000000000000;
		44719: Delta = 69'sb000100000000000000000100000000000000000000000000000000000000000000000;
		198: Delta = 69'sb111100000000000000000100000000000000000000000000000000000000000000000;
		50663: Delta = 69'sb000011111111111111111100000000000000000000000000000000000000000000000;
		6142: Delta = 69'sb111011111111111111111100000000000000000000000000000000000000000000000;
		41549: Delta = 69'sb001000000000000000000100000000000000000000000000000000000000000000000;
		3368: Delta = 69'sb111000000000000000000100000000000000000000000000000000000000000000000;
		47493: Delta = 69'sb000111111111111111111100000000000000000000000000000000000000000000000;
		9312: Delta = 69'sb110111111111111111111100000000000000000000000000000000000000000000000;
		35209: Delta = 69'sb010000000000000000000100000000000000000000000000000000000000000000000;
		9708: Delta = 69'sb110000000000000000000100000000000000000000000000000000000000000000000;
		41153: Delta = 69'sb001111111111111111111100000000000000000000000000000000000000000000000;
		15652: Delta = 69'sb101111111111111111111100000000000000000000000000000000000000000000000;
		33029: Delta = 69'sb000000000000000000011000000000000000000000000000000000000000000000000;
		17832: Delta = 69'sb111111111111111111101000000000000000000000000000000000000000000000000;
		21141: Delta = 69'sb000000000000000000101000000000000000000000000000000000000000000000000;
		29720: Delta = 69'sb111111111111111111011000000000000000000000000000000000000000000000000;
		48226: Delta = 69'sb000000000000000001001000000000000000000000000000000000000000000000000;
		41608: Delta = 69'sb111111111111111111001000000000000000000000000000000000000000000000000;
		9253: Delta = 69'sb000000000000000000111000000000000000000000000000000000000000000000000;
		2635: Delta = 69'sb111111111111111110111000000000000000000000000000000000000000000000000;
		674: Delta = 69'sb000000000000000010001000000000000000000000000000000000000000000000000;
		38299: Delta = 69'sb111111111111111110001000000000000000000000000000000000000000000000000;
		12562: Delta = 69'sb000000000000000001111000000000000000000000000000000000000000000000000;
		50187: Delta = 69'sb111111111111111101111000000000000000000000000000000000000000000000000;
		7292: Delta = 69'sb000000000000000100001000000000000000000000000000000000000000000000000;
		31681: Delta = 69'sb111111111111111100001000000000000000000000000000000000000000000000000;
		19180: Delta = 69'sb000000000000000011111000000000000000000000000000000000000000000000000;
		43569: Delta = 69'sb111111111111111011111000000000000000000000000000000000000000000000000;
		20528: Delta = 69'sb000000000000001000001000000000000000000000000000000000000000000000000;
		18445: Delta = 69'sb111111111111111000001000000000000000000000000000000000000000000000000;
		32416: Delta = 69'sb000000000000000111111000000000000000000000000000000000000000000000000;
		30333: Delta = 69'sb111111111111110111111000000000000000000000000000000000000000000000000;
		47000: Delta = 69'sb000000000000010000001000000000000000000000000000000000000000000000000;
		42834: Delta = 69'sb111111111111110000001000000000000000000000000000000000000000000000000;
		8027: Delta = 69'sb000000000000001111111000000000000000000000000000000000000000000000000;
		3861: Delta = 69'sb111111111111101111111000000000000000000000000000000000000000000000000;
		49083: Delta = 69'sb000000000000100000001000000000000000000000000000000000000000000000000;
		40751: Delta = 69'sb111111111111100000001000000000000000000000000000000000000000000000000;
		10110: Delta = 69'sb000000000000011111111000000000000000000000000000000000000000000000000;
		1778: Delta = 69'sb111111111111011111111000000000000000000000000000000000000000000000000;
		2388: Delta = 69'sb000000000001000000001000000000000000000000000000000000000000000000000;
		36585: Delta = 69'sb111111111111000000001000000000000000000000000000000000000000000000000;
		14276: Delta = 69'sb000000000000111111111000000000000000000000000000000000000000000000000;
		48473: Delta = 69'sb111111111110111111111000000000000000000000000000000000000000000000000;
		10720: Delta = 69'sb000000000010000000001000000000000000000000000000000000000000000000000;
		28253: Delta = 69'sb111111111110000000001000000000000000000000000000000000000000000000000;
		22608: Delta = 69'sb000000000001111111111000000000000000000000000000000000000000000000000;
		40141: Delta = 69'sb111111111101111111111000000000000000000000000000000000000000000000000;
		27384: Delta = 69'sb000000000100000000001000000000000000000000000000000000000000000000000;
		11589: Delta = 69'sb111111111100000000001000000000000000000000000000000000000000000000000;
		39272: Delta = 69'sb000000000011111111111000000000000000000000000000000000000000000000000;
		23477: Delta = 69'sb111111111011111111111000000000000000000000000000000000000000000000000;
		9851: Delta = 69'sb000000001000000000001000000000000000000000000000000000000000000000000;
		29122: Delta = 69'sb111111111000000000001000000000000000000000000000000000000000000000000;
		21739: Delta = 69'sb000000000111111111111000000000000000000000000000000000000000000000000;
		41010: Delta = 69'sb111111110111111111111000000000000000000000000000000000000000000000000;
		25646: Delta = 69'sb000000010000000000001000000000000000000000000000000000000000000000000;
		13327: Delta = 69'sb111111110000000000001000000000000000000000000000000000000000000000000;
		37534: Delta = 69'sb000000001111111111111000000000000000000000000000000000000000000000000;
		25215: Delta = 69'sb111111101111111111111000000000000000000000000000000000000000000000000;
		6375: Delta = 69'sb000000100000000000001000000000000000000000000000000000000000000000000;
		32598: Delta = 69'sb111111100000000000001000000000000000000000000000000000000000000000000;
		18263: Delta = 69'sb000000011111111111111000000000000000000000000000000000000000000000000;
		44486: Delta = 69'sb111111011111111111111000000000000000000000000000000000000000000000000;
		18694: Delta = 69'sb000001000000000000001000000000000000000000000000000000000000000000000;
		20279: Delta = 69'sb111111000000000000001000000000000000000000000000000000000000000000000;
		30582: Delta = 69'sb000000111111111111111000000000000000000000000000000000000000000000000;
		32167: Delta = 69'sb111110111111111111111000000000000000000000000000000000000000000000000;
		43332: Delta = 69'sb000010000000000000001000000000000000000000000000000000000000000000000;
		46502: Delta = 69'sb111110000000000000001000000000000000000000000000000000000000000000000;
		4359: Delta = 69'sb000001111111111111111000000000000000000000000000000000000000000000000;
		7529: Delta = 69'sb111101111111111111111000000000000000000000000000000000000000000000000;
		41747: Delta = 69'sb000100000000000000001000000000000000000000000000000000000000000000000;
		48087: Delta = 69'sb111100000000000000001000000000000000000000000000000000000000000000000;
		2774: Delta = 69'sb000011111111111111111000000000000000000000000000000000000000000000000;
		9114: Delta = 69'sb111011111111111111111000000000000000000000000000000000000000000000000;
		38577: Delta = 69'sb001000000000000000001000000000000000000000000000000000000000000000000;
		396: Delta = 69'sb111000000000000000001000000000000000000000000000000000000000000000000;
		50465: Delta = 69'sb000111111111111111111000000000000000000000000000000000000000000000000;
		12284: Delta = 69'sb110111111111111111111000000000000000000000000000000000000000000000000;
		32237: Delta = 69'sb010000000000000000001000000000000000000000000000000000000000000000000;
		6736: Delta = 69'sb110000000000000000001000000000000000000000000000000000000000000000000;
		44125: Delta = 69'sb001111111111111111111000000000000000000000000000000000000000000000000;
		18624: Delta = 69'sb101111111111111111111000000000000000000000000000000000000000000000000;
		15197: Delta = 69'sb000000000000000000110000000000000000000000000000000000000000000000000;
		35664: Delta = 69'sb111111111111111111010000000000000000000000000000000000000000000000000;
		42282: Delta = 69'sb000000000000000001010000000000000000000000000000000000000000000000000;
		8579: Delta = 69'sb111111111111111110110000000000000000000000000000000000000000000000000;
		45591: Delta = 69'sb000000000000000010010000000000000000000000000000000000000000000000000;
		32355: Delta = 69'sb111111111111111110010000000000000000000000000000000000000000000000000;
		18506: Delta = 69'sb000000000000000001110000000000000000000000000000000000000000000000000;
		5270: Delta = 69'sb111111111111111101110000000000000000000000000000000000000000000000000;
		1348: Delta = 69'sb000000000000000100010000000000000000000000000000000000000000000000000;
		25737: Delta = 69'sb111111111111111100010000000000000000000000000000000000000000000000000;
		25124: Delta = 69'sb000000000000000011110000000000000000000000000000000000000000000000000;
		49513: Delta = 69'sb111111111111111011110000000000000000000000000000000000000000000000000;
		14584: Delta = 69'sb000000000000001000010000000000000000000000000000000000000000000000000;
		12501: Delta = 69'sb111111111111111000010000000000000000000000000000000000000000000000000;
		38360: Delta = 69'sb000000000000000111110000000000000000000000000000000000000000000000000;
		36277: Delta = 69'sb111111111111110111110000000000000000000000000000000000000000000000000;
		41056: Delta = 69'sb000000000000010000010000000000000000000000000000000000000000000000000;
		36890: Delta = 69'sb111111111111110000010000000000000000000000000000000000000000000000000;
		13971: Delta = 69'sb000000000000001111110000000000000000000000000000000000000000000000000;
		9805: Delta = 69'sb111111111111101111110000000000000000000000000000000000000000000000000;
		43139: Delta = 69'sb000000000000100000010000000000000000000000000000000000000000000000000;
		34807: Delta = 69'sb111111111111100000010000000000000000000000000000000000000000000000000;
		16054: Delta = 69'sb000000000000011111110000000000000000000000000000000000000000000000000;
		7722: Delta = 69'sb111111111111011111110000000000000000000000000000000000000000000000000;
		47305: Delta = 69'sb000000000001000000010000000000000000000000000000000000000000000000000;
		30641: Delta = 69'sb111111111111000000010000000000000000000000000000000000000000000000000;
		20220: Delta = 69'sb000000000000111111110000000000000000000000000000000000000000000000000;
		3556: Delta = 69'sb111111111110111111110000000000000000000000000000000000000000000000000;
		4776: Delta = 69'sb000000000010000000010000000000000000000000000000000000000000000000000;
		22309: Delta = 69'sb111111111110000000010000000000000000000000000000000000000000000000000;
		28552: Delta = 69'sb000000000001111111110000000000000000000000000000000000000000000000000;
		46085: Delta = 69'sb111111111101111111110000000000000000000000000000000000000000000000000;
		21440: Delta = 69'sb000000000100000000010000000000000000000000000000000000000000000000000;
		5645: Delta = 69'sb111111111100000000010000000000000000000000000000000000000000000000000;
		45216: Delta = 69'sb000000000011111111110000000000000000000000000000000000000000000000000;
		29421: Delta = 69'sb111111111011111111110000000000000000000000000000000000000000000000000;
		3907: Delta = 69'sb000000001000000000010000000000000000000000000000000000000000000000000;
		23178: Delta = 69'sb111111111000000000010000000000000000000000000000000000000000000000000;
		27683: Delta = 69'sb000000000111111111110000000000000000000000000000000000000000000000000;
		46954: Delta = 69'sb111111110111111111110000000000000000000000000000000000000000000000000;
		19702: Delta = 69'sb000000010000000000010000000000000000000000000000000000000000000000000;
		7383: Delta = 69'sb111111110000000000010000000000000000000000000000000000000000000000000;
		43478: Delta = 69'sb000000001111111111110000000000000000000000000000000000000000000000000;
		31159: Delta = 69'sb111111101111111111110000000000000000000000000000000000000000000000000;
		431: Delta = 69'sb000000100000000000010000000000000000000000000000000000000000000000000;
		26654: Delta = 69'sb111111100000000000010000000000000000000000000000000000000000000000000;
		24207: Delta = 69'sb000000011111111111110000000000000000000000000000000000000000000000000;
		50430: Delta = 69'sb111111011111111111110000000000000000000000000000000000000000000000000;
		12750: Delta = 69'sb000001000000000000010000000000000000000000000000000000000000000000000;
		14335: Delta = 69'sb111111000000000000010000000000000000000000000000000000000000000000000;
		36526: Delta = 69'sb000000111111111111110000000000000000000000000000000000000000000000000;
		38111: Delta = 69'sb111110111111111111110000000000000000000000000000000000000000000000000;
		37388: Delta = 69'sb000010000000000000010000000000000000000000000000000000000000000000000;
		40558: Delta = 69'sb111110000000000000010000000000000000000000000000000000000000000000000;
		10303: Delta = 69'sb000001111111111111110000000000000000000000000000000000000000000000000;
		13473: Delta = 69'sb111101111111111111110000000000000000000000000000000000000000000000000;
		35803: Delta = 69'sb000100000000000000010000000000000000000000000000000000000000000000000;
		42143: Delta = 69'sb111100000000000000010000000000000000000000000000000000000000000000000;
		8718: Delta = 69'sb000011111111111111110000000000000000000000000000000000000000000000000;
		15058: Delta = 69'sb111011111111111111110000000000000000000000000000000000000000000000000;
		32633: Delta = 69'sb001000000000000000010000000000000000000000000000000000000000000000000;
		45313: Delta = 69'sb111000000000000000010000000000000000000000000000000000000000000000000;
		5548: Delta = 69'sb000111111111111111110000000000000000000000000000000000000000000000000;
		18228: Delta = 69'sb110111111111111111110000000000000000000000000000000000000000000000000;
		26293: Delta = 69'sb010000000000000000010000000000000000000000000000000000000000000000000;
		792: Delta = 69'sb110000000000000000010000000000000000000000000000000000000000000000000;
		50069: Delta = 69'sb001111111111111111110000000000000000000000000000000000000000000000000;
		24568: Delta = 69'sb101111111111111111110000000000000000000000000000000000000000000000000;
		30394: Delta = 69'sb000000000000000001100000000000000000000000000000000000000000000000000;
		20467: Delta = 69'sb111111111111111110100000000000000000000000000000000000000000000000000;
		33703: Delta = 69'sb000000000000000010100000000000000000000000000000000000000000000000000;
		17158: Delta = 69'sb111111111111111101100000000000000000000000000000000000000000000000000;
		40321: Delta = 69'sb000000000000000100100000000000000000000000000000000000000000000000000;
		13849: Delta = 69'sb111111111111111100100000000000000000000000000000000000000000000000000;
		37012: Delta = 69'sb000000000000000011100000000000000000000000000000000000000000000000000;
		10540: Delta = 69'sb111111111111111011100000000000000000000000000000000000000000000000000;
		2696: Delta = 69'sb000000000000001000100000000000000000000000000000000000000000000000000;
		613: Delta = 69'sb111111111111111000100000000000000000000000000000000000000000000000000;
		50248: Delta = 69'sb000000000000000111100000000000000000000000000000000000000000000000000;
		48165: Delta = 69'sb111111111111110111100000000000000000000000000000000000000000000000000;
		29168: Delta = 69'sb000000000000010000100000000000000000000000000000000000000000000000000;
		25002: Delta = 69'sb111111111111110000100000000000000000000000000000000000000000000000000;
		25859: Delta = 69'sb000000000000001111100000000000000000000000000000000000000000000000000;
		21693: Delta = 69'sb111111111111101111100000000000000000000000000000000000000000000000000;
		31251: Delta = 69'sb000000000000100000100000000000000000000000000000000000000000000000000;
		22919: Delta = 69'sb111111111111100000100000000000000000000000000000000000000000000000000;
		27942: Delta = 69'sb000000000000011111100000000000000000000000000000000000000000000000000;
		19610: Delta = 69'sb111111111111011111100000000000000000000000000000000000000000000000000;
		35417: Delta = 69'sb000000000001000000100000000000000000000000000000000000000000000000000;
		18753: Delta = 69'sb111111111111000000100000000000000000000000000000000000000000000000000;
		32108: Delta = 69'sb000000000000111111100000000000000000000000000000000000000000000000000;
		15444: Delta = 69'sb111111111110111111100000000000000000000000000000000000000000000000000;
		43749: Delta = 69'sb000000000010000000100000000000000000000000000000000000000000000000000;
		10421: Delta = 69'sb111111111110000000100000000000000000000000000000000000000000000000000;
		40440: Delta = 69'sb000000000001111111100000000000000000000000000000000000000000000000000;
		7112: Delta = 69'sb111111111101111111100000000000000000000000000000000000000000000000000;
		9552: Delta = 69'sb000000000100000000100000000000000000000000000000000000000000000000000;
		44618: Delta = 69'sb111111111100000000100000000000000000000000000000000000000000000000000;
		6243: Delta = 69'sb000000000011111111100000000000000000000000000000000000000000000000000;
		41309: Delta = 69'sb111111111011111111100000000000000000000000000000000000000000000000000;
		42880: Delta = 69'sb000000001000000000100000000000000000000000000000000000000000000000000;
		11290: Delta = 69'sb111111111000000000100000000000000000000000000000000000000000000000000;
		39571: Delta = 69'sb000000000111111111100000000000000000000000000000000000000000000000000;
		7981: Delta = 69'sb111111110111111111100000000000000000000000000000000000000000000000000;
		7814: Delta = 69'sb000000010000000000100000000000000000000000000000000000000000000000000;
		46356: Delta = 69'sb111111110000000000100000000000000000000000000000000000000000000000000;
		4505: Delta = 69'sb000000001111111111100000000000000000000000000000000000000000000000000;
		43047: Delta = 69'sb111111101111111111100000000000000000000000000000000000000000000000000;
		39404: Delta = 69'sb000000100000000000100000000000000000000000000000000000000000000000000;
		14766: Delta = 69'sb111111100000000000100000000000000000000000000000000000000000000000000;
		36095: Delta = 69'sb000000011111111111100000000000000000000000000000000000000000000000000;
		11457: Delta = 69'sb111111011111111111100000000000000000000000000000000000000000000000000;
		862: Delta = 69'sb000001000000000000100000000000000000000000000000000000000000000000000;
		2447: Delta = 69'sb111111000000000000100000000000000000000000000000000000000000000000000;
		48414: Delta = 69'sb000000111111111111100000000000000000000000000000000000000000000000000;
		49999: Delta = 69'sb111110111111111111100000000000000000000000000000000000000000000000000;
		25500: Delta = 69'sb000010000000000000100000000000000000000000000000000000000000000000000;
		28670: Delta = 69'sb111110000000000000100000000000000000000000000000000000000000000000000;
		22191: Delta = 69'sb000001111111111111100000000000000000000000000000000000000000000000000;
		25361: Delta = 69'sb111101111111111111100000000000000000000000000000000000000000000000000;
		23915: Delta = 69'sb000100000000000000100000000000000000000000000000000000000000000000000;
		30255: Delta = 69'sb111100000000000000100000000000000000000000000000000000000000000000000;
		20606: Delta = 69'sb000011111111111111100000000000000000000000000000000000000000000000000;
		26946: Delta = 69'sb111011111111111111100000000000000000000000000000000000000000000000000;
		20745: Delta = 69'sb001000000000000000100000000000000000000000000000000000000000000000000;
		33425: Delta = 69'sb111000000000000000100000000000000000000000000000000000000000000000000;
		17436: Delta = 69'sb000111111111111111100000000000000000000000000000000000000000000000000;
		30116: Delta = 69'sb110111111111111111100000000000000000000000000000000000000000000000000;
		14405: Delta = 69'sb010000000000000000100000000000000000000000000000000000000000000000000;
		39765: Delta = 69'sb110000000000000000100000000000000000000000000000000000000000000000000;
		11096: Delta = 69'sb001111111111111111100000000000000000000000000000000000000000000000000;
		36456: Delta = 69'sb101111111111111111100000000000000000000000000000000000000000000000000;
		9927: Delta = 69'sb000000000000000011000000000000000000000000000000000000000000000000000;
		40934: Delta = 69'sb111111111111111101000000000000000000000000000000000000000000000000000;
		16545: Delta = 69'sb000000000000000101000000000000000000000000000000000000000000000000000;
		34316: Delta = 69'sb111111111111111011000000000000000000000000000000000000000000000000000;
		29781: Delta = 69'sb000000000000001001000000000000000000000000000000000000000000000000000;
		27698: Delta = 69'sb111111111111111001000000000000000000000000000000000000000000000000000;
		23163: Delta = 69'sb000000000000000111000000000000000000000000000000000000000000000000000;
		21080: Delta = 69'sb111111111111110111000000000000000000000000000000000000000000000000000;
		5392: Delta = 69'sb000000000000010001000000000000000000000000000000000000000000000000000;
		1226: Delta = 69'sb111111111111110001000000000000000000000000000000000000000000000000000;
		49635: Delta = 69'sb000000000000001111000000000000000000000000000000000000000000000000000;
		45469: Delta = 69'sb111111111111101111000000000000000000000000000000000000000000000000000;
		7475: Delta = 69'sb000000000000100001000000000000000000000000000000000000000000000000000;
		50004: Delta = 69'sb111111111111100001000000000000000000000000000000000000000000000000000;
		857: Delta = 69'sb000000000000011111000000000000000000000000000000000000000000000000000;
		43386: Delta = 69'sb111111111111011111000000000000000000000000000000000000000000000000000;
		11641: Delta = 69'sb000000000001000001000000000000000000000000000000000000000000000000000;
		45838: Delta = 69'sb111111111111000001000000000000000000000000000000000000000000000000000;
		5023: Delta = 69'sb000000000000111111000000000000000000000000000000000000000000000000000;
		39220: Delta = 69'sb111111111110111111000000000000000000000000000000000000000000000000000;
		19973: Delta = 69'sb000000000010000001000000000000000000000000000000000000000000000000000;
		37506: Delta = 69'sb111111111110000001000000000000000000000000000000000000000000000000000;
		13355: Delta = 69'sb000000000001111111000000000000000000000000000000000000000000000000000;
		30888: Delta = 69'sb111111111101111111000000000000000000000000000000000000000000000000000;
		36637: Delta = 69'sb000000000100000001000000000000000000000000000000000000000000000000000;
		20842: Delta = 69'sb111111111100000001000000000000000000000000000000000000000000000000000;
		30019: Delta = 69'sb000000000011111111000000000000000000000000000000000000000000000000000;
		14224: Delta = 69'sb111111111011111111000000000000000000000000000000000000000000000000000;
		19104: Delta = 69'sb000000001000000001000000000000000000000000000000000000000000000000000;
		38375: Delta = 69'sb111111111000000001000000000000000000000000000000000000000000000000000;
		12486: Delta = 69'sb000000000111111111000000000000000000000000000000000000000000000000000;
		31757: Delta = 69'sb111111110111111111000000000000000000000000000000000000000000000000000;
		34899: Delta = 69'sb000000010000000001000000000000000000000000000000000000000000000000000;
		22580: Delta = 69'sb111111110000000001000000000000000000000000000000000000000000000000000;
		28281: Delta = 69'sb000000001111111111000000000000000000000000000000000000000000000000000;
		15962: Delta = 69'sb111111101111111111000000000000000000000000000000000000000000000000000;
		15628: Delta = 69'sb000000100000000001000000000000000000000000000000000000000000000000000;
		41851: Delta = 69'sb111111100000000001000000000000000000000000000000000000000000000000000;
		9010: Delta = 69'sb000000011111111111000000000000000000000000000000000000000000000000000;
		35233: Delta = 69'sb111111011111111111000000000000000000000000000000000000000000000000000;
		27947: Delta = 69'sb000001000000000001000000000000000000000000000000000000000000000000000;
		29532: Delta = 69'sb111111000000000001000000000000000000000000000000000000000000000000000;
		21329: Delta = 69'sb000000111111111111000000000000000000000000000000000000000000000000000;
		22914: Delta = 69'sb111110111111111111000000000000000000000000000000000000000000000000000;
		1724: Delta = 69'sb000010000000000001000000000000000000000000000000000000000000000000000;
		4894: Delta = 69'sb111110000000000001000000000000000000000000000000000000000000000000000;
		45967: Delta = 69'sb000001111111111111000000000000000000000000000000000000000000000000000;
		49137: Delta = 69'sb111101111111111111000000000000000000000000000000000000000000000000000;
		139: Delta = 69'sb000100000000000001000000000000000000000000000000000000000000000000000;
		6479: Delta = 69'sb111100000000000001000000000000000000000000000000000000000000000000000;
		44382: Delta = 69'sb000011111111111111000000000000000000000000000000000000000000000000000;
		50722: Delta = 69'sb111011111111111111000000000000000000000000000000000000000000000000000;
		47830: Delta = 69'sb001000000000000001000000000000000000000000000000000000000000000000000;
		9649: Delta = 69'sb111000000000000001000000000000000000000000000000000000000000000000000;
		41212: Delta = 69'sb000111111111111111000000000000000000000000000000000000000000000000000;
		3031: Delta = 69'sb110111111111111111000000000000000000000000000000000000000000000000000;
		41490: Delta = 69'sb010000000000000001000000000000000000000000000000000000000000000000000;
		15989: Delta = 69'sb110000000000000001000000000000000000000000000000000000000000000000000;
		34872: Delta = 69'sb001111111111111111000000000000000000000000000000000000000000000000000;
		9371: Delta = 69'sb101111111111111111000000000000000000000000000000000000000000000000000;
		19854: Delta = 69'sb000000000000000110000000000000000000000000000000000000000000000000000;
		31007: Delta = 69'sb111111111111111010000000000000000000000000000000000000000000000000000;
		33090: Delta = 69'sb000000000000001010000000000000000000000000000000000000000000000000000;
		17771: Delta = 69'sb111111111111110110000000000000000000000000000000000000000000000000000;
		8701: Delta = 69'sb000000000000010010000000000000000000000000000000000000000000000000000;
		4535: Delta = 69'sb111111111111110010000000000000000000000000000000000000000000000000000;
		46326: Delta = 69'sb000000000000001110000000000000000000000000000000000000000000000000000;
		42160: Delta = 69'sb111111111111101110000000000000000000000000000000000000000000000000000;
		10784: Delta = 69'sb000000000000100010000000000000000000000000000000000000000000000000000;
		2452: Delta = 69'sb111111111111100010000000000000000000000000000000000000000000000000000;
		48409: Delta = 69'sb000000000000011110000000000000000000000000000000000000000000000000000;
		40077: Delta = 69'sb111111111111011110000000000000000000000000000000000000000000000000000;
		14950: Delta = 69'sb000000000001000010000000000000000000000000000000000000000000000000000;
		49147: Delta = 69'sb111111111111000010000000000000000000000000000000000000000000000000000;
		1714: Delta = 69'sb000000000000111110000000000000000000000000000000000000000000000000000;
		35911: Delta = 69'sb111111111110111110000000000000000000000000000000000000000000000000000;
		23282: Delta = 69'sb000000000010000010000000000000000000000000000000000000000000000000000;
		40815: Delta = 69'sb111111111110000010000000000000000000000000000000000000000000000000000;
		10046: Delta = 69'sb000000000001111110000000000000000000000000000000000000000000000000000;
		27579: Delta = 69'sb111111111101111110000000000000000000000000000000000000000000000000000;
		39946: Delta = 69'sb000000000100000010000000000000000000000000000000000000000000000000000;
		24151: Delta = 69'sb111111111100000010000000000000000000000000000000000000000000000000000;
		26710: Delta = 69'sb000000000011111110000000000000000000000000000000000000000000000000000;
		10915: Delta = 69'sb111111111011111110000000000000000000000000000000000000000000000000000;
		22413: Delta = 69'sb000000001000000010000000000000000000000000000000000000000000000000000;
		41684: Delta = 69'sb111111111000000010000000000000000000000000000000000000000000000000000;
		9177: Delta = 69'sb000000000111111110000000000000000000000000000000000000000000000000000;
		28448: Delta = 69'sb111111110111111110000000000000000000000000000000000000000000000000000;
		38208: Delta = 69'sb000000010000000010000000000000000000000000000000000000000000000000000;
		25889: Delta = 69'sb111111110000000010000000000000000000000000000000000000000000000000000;
		24972: Delta = 69'sb000000001111111110000000000000000000000000000000000000000000000000000;
		12653: Delta = 69'sb111111101111111110000000000000000000000000000000000000000000000000000;
		18937: Delta = 69'sb000000100000000010000000000000000000000000000000000000000000000000000;
		45160: Delta = 69'sb111111100000000010000000000000000000000000000000000000000000000000000;
		5701: Delta = 69'sb000000011111111110000000000000000000000000000000000000000000000000000;
		31924: Delta = 69'sb111111011111111110000000000000000000000000000000000000000000000000000;
		31256: Delta = 69'sb000001000000000010000000000000000000000000000000000000000000000000000;
		32841: Delta = 69'sb111111000000000010000000000000000000000000000000000000000000000000000;
		18020: Delta = 69'sb000000111111111110000000000000000000000000000000000000000000000000000;
		19605: Delta = 69'sb111110111111111110000000000000000000000000000000000000000000000000000;
		5033: Delta = 69'sb000010000000000010000000000000000000000000000000000000000000000000000;
		8203: Delta = 69'sb111110000000000010000000000000000000000000000000000000000000000000000;
		42658: Delta = 69'sb000001111111111110000000000000000000000000000000000000000000000000000;
		45828: Delta = 69'sb111101111111111110000000000000000000000000000000000000000000000000000;
		3448: Delta = 69'sb000100000000000010000000000000000000000000000000000000000000000000000;
		9788: Delta = 69'sb111100000000000010000000000000000000000000000000000000000000000000000;
		41073: Delta = 69'sb000011111111111110000000000000000000000000000000000000000000000000000;
		47413: Delta = 69'sb111011111111111110000000000000000000000000000000000000000000000000000;
		278: Delta = 69'sb001000000000000010000000000000000000000000000000000000000000000000000;
		12958: Delta = 69'sb111000000000000010000000000000000000000000000000000000000000000000000;
		37903: Delta = 69'sb000111111111111110000000000000000000000000000000000000000000000000000;
		50583: Delta = 69'sb110111111111111110000000000000000000000000000000000000000000000000000;
		44799: Delta = 69'sb010000000000000010000000000000000000000000000000000000000000000000000;
		19298: Delta = 69'sb110000000000000010000000000000000000000000000000000000000000000000000;
		31563: Delta = 69'sb001111111111111110000000000000000000000000000000000000000000000000000;
		6062: Delta = 69'sb101111111111111110000000000000000000000000000000000000000000000000000;
		39708: Delta = 69'sb000000000000001100000000000000000000000000000000000000000000000000000;
		11153: Delta = 69'sb111111111111110100000000000000000000000000000000000000000000000000000;
		15319: Delta = 69'sb000000000000010100000000000000000000000000000000000000000000000000000;
		35542: Delta = 69'sb111111111111101100000000000000000000000000000000000000000000000000000;
		17402: Delta = 69'sb000000000000100100000000000000000000000000000000000000000000000000000;
		9070: Delta = 69'sb111111111111100100000000000000000000000000000000000000000000000000000;
		41791: Delta = 69'sb000000000000011100000000000000000000000000000000000000000000000000000;
		33459: Delta = 69'sb111111111111011100000000000000000000000000000000000000000000000000000;
		21568: Delta = 69'sb000000000001000100000000000000000000000000000000000000000000000000000;
		4904: Delta = 69'sb111111111111000100000000000000000000000000000000000000000000000000000;
		45957: Delta = 69'sb000000000000111100000000000000000000000000000000000000000000000000000;
		29293: Delta = 69'sb111111111110111100000000000000000000000000000000000000000000000000000;
		29900: Delta = 69'sb000000000010000100000000000000000000000000000000000000000000000000000;
		47433: Delta = 69'sb111111111110000100000000000000000000000000000000000000000000000000000;
		3428: Delta = 69'sb000000000001111100000000000000000000000000000000000000000000000000000;
		20961: Delta = 69'sb111111111101111100000000000000000000000000000000000000000000000000000;
		46564: Delta = 69'sb000000000100000100000000000000000000000000000000000000000000000000000;
		30769: Delta = 69'sb111111111100000100000000000000000000000000000000000000000000000000000;
		20092: Delta = 69'sb000000000011111100000000000000000000000000000000000000000000000000000;
		4297: Delta = 69'sb111111111011111100000000000000000000000000000000000000000000000000000;
		29031: Delta = 69'sb000000001000000100000000000000000000000000000000000000000000000000000;
		48302: Delta = 69'sb111111111000000100000000000000000000000000000000000000000000000000000;
		2559: Delta = 69'sb000000000111111100000000000000000000000000000000000000000000000000000;
		21830: Delta = 69'sb111111110111111100000000000000000000000000000000000000000000000000000;
		44826: Delta = 69'sb000000010000000100000000000000000000000000000000000000000000000000000;
		32507: Delta = 69'sb111111110000000100000000000000000000000000000000000000000000000000000;
		18354: Delta = 69'sb000000001111111100000000000000000000000000000000000000000000000000000;
		6035: Delta = 69'sb111111101111111100000000000000000000000000000000000000000000000000000;
		25555: Delta = 69'sb000000100000000100000000000000000000000000000000000000000000000000000;
		917: Delta = 69'sb111111100000000100000000000000000000000000000000000000000000000000000;
		49944: Delta = 69'sb000000011111111100000000000000000000000000000000000000000000000000000;
		25306: Delta = 69'sb111111011111111100000000000000000000000000000000000000000000000000000;
		37874: Delta = 69'sb000001000000000100000000000000000000000000000000000000000000000000000;
		39459: Delta = 69'sb111111000000000100000000000000000000000000000000000000000000000000000;
		11402: Delta = 69'sb000000111111111100000000000000000000000000000000000000000000000000000;
		12987: Delta = 69'sb111110111111111100000000000000000000000000000000000000000000000000000;
		11651: Delta = 69'sb000010000000000100000000000000000000000000000000000000000000000000000;
		14821: Delta = 69'sb111110000000000100000000000000000000000000000000000000000000000000000;
		36040: Delta = 69'sb000001111111111100000000000000000000000000000000000000000000000000000;
		39210: Delta = 69'sb111101111111111100000000000000000000000000000000000000000000000000000;
		10066: Delta = 69'sb000100000000000100000000000000000000000000000000000000000000000000000;
		16406: Delta = 69'sb111100000000000100000000000000000000000000000000000000000000000000000;
		34455: Delta = 69'sb000011111111111100000000000000000000000000000000000000000000000000000;
		40795: Delta = 69'sb111011111111111100000000000000000000000000000000000000000000000000000;
		6896: Delta = 69'sb001000000000000100000000000000000000000000000000000000000000000000000;
		19576: Delta = 69'sb111000000000000100000000000000000000000000000000000000000000000000000;
		31285: Delta = 69'sb000111111111111100000000000000000000000000000000000000000000000000000;
		43965: Delta = 69'sb110111111111111100000000000000000000000000000000000000000000000000000;
		556: Delta = 69'sb010000000000000100000000000000000000000000000000000000000000000000000;
		25916: Delta = 69'sb110000000000000100000000000000000000000000000000000000000000000000000;
		24945: Delta = 69'sb001111111111111100000000000000000000000000000000000000000000000000000;
		50305: Delta = 69'sb101111111111111100000000000000000000000000000000000000000000000000000;
		28555: Delta = 69'sb000000000000011000000000000000000000000000000000000000000000000000000;
		22306: Delta = 69'sb111111111111101000000000000000000000000000000000000000000000000000000;
		30638: Delta = 69'sb000000000000101000000000000000000000000000000000000000000000000000000;
		20223: Delta = 69'sb111111111111011000000000000000000000000000000000000000000000000000000;
		34804: Delta = 69'sb000000000001001000000000000000000000000000000000000000000000000000000;
		18140: Delta = 69'sb111111111111001000000000000000000000000000000000000000000000000000000;
		32721: Delta = 69'sb000000000000111000000000000000000000000000000000000000000000000000000;
		16057: Delta = 69'sb111111111110111000000000000000000000000000000000000000000000000000000;
		43136: Delta = 69'sb000000000010001000000000000000000000000000000000000000000000000000000;
		9808: Delta = 69'sb111111111110001000000000000000000000000000000000000000000000000000000;
		41053: Delta = 69'sb000000000001111000000000000000000000000000000000000000000000000000000;
		7725: Delta = 69'sb111111111101111000000000000000000000000000000000000000000000000000000;
		8939: Delta = 69'sb000000000100001000000000000000000000000000000000000000000000000000000;
		44005: Delta = 69'sb111111111100001000000000000000000000000000000000000000000000000000000;
		6856: Delta = 69'sb000000000011111000000000000000000000000000000000000000000000000000000;
		41922: Delta = 69'sb111111111011111000000000000000000000000000000000000000000000000000000;
		42267: Delta = 69'sb000000001000001000000000000000000000000000000000000000000000000000000;
		10677: Delta = 69'sb111111111000001000000000000000000000000000000000000000000000000000000;
		40184: Delta = 69'sb000000000111111000000000000000000000000000000000000000000000000000000;
		8594: Delta = 69'sb111111110111111000000000000000000000000000000000000000000000000000000;
		7201: Delta = 69'sb000000010000001000000000000000000000000000000000000000000000000000000;
		45743: Delta = 69'sb111111110000001000000000000000000000000000000000000000000000000000000;
		5118: Delta = 69'sb000000001111111000000000000000000000000000000000000000000000000000000;
		43660: Delta = 69'sb111111101111111000000000000000000000000000000000000000000000000000000;
		38791: Delta = 69'sb000000100000001000000000000000000000000000000000000000000000000000000;
		14153: Delta = 69'sb111111100000001000000000000000000000000000000000000000000000000000000;
		36708: Delta = 69'sb000000011111111000000000000000000000000000000000000000000000000000000;
		12070: Delta = 69'sb111111011111111000000000000000000000000000000000000000000000000000000;
		249: Delta = 69'sb000001000000001000000000000000000000000000000000000000000000000000000;
		1834: Delta = 69'sb111111000000001000000000000000000000000000000000000000000000000000000;
		49027: Delta = 69'sb000000111111111000000000000000000000000000000000000000000000000000000;
		50612: Delta = 69'sb111110111111111000000000000000000000000000000000000000000000000000000;
		24887: Delta = 69'sb000010000000001000000000000000000000000000000000000000000000000000000;
		28057: Delta = 69'sb111110000000001000000000000000000000000000000000000000000000000000000;
		22804: Delta = 69'sb000001111111111000000000000000000000000000000000000000000000000000000;
		25974: Delta = 69'sb111101111111111000000000000000000000000000000000000000000000000000000;
		23302: Delta = 69'sb000100000000001000000000000000000000000000000000000000000000000000000;
		29642: Delta = 69'sb111100000000001000000000000000000000000000000000000000000000000000000;
		21219: Delta = 69'sb000011111111111000000000000000000000000000000000000000000000000000000;
		27559: Delta = 69'sb111011111111111000000000000000000000000000000000000000000000000000000;
		20132: Delta = 69'sb001000000000001000000000000000000000000000000000000000000000000000000;
		32812: Delta = 69'sb111000000000001000000000000000000000000000000000000000000000000000000;
		18049: Delta = 69'sb000111111111111000000000000000000000000000000000000000000000000000000;
		30729: Delta = 69'sb110111111111111000000000000000000000000000000000000000000000000000000;
		13792: Delta = 69'sb010000000000001000000000000000000000000000000000000000000000000000000;
		39152: Delta = 69'sb110000000000001000000000000000000000000000000000000000000000000000000;
		11709: Delta = 69'sb001111111111111000000000000000000000000000000000000000000000000000000;
		37069: Delta = 69'sb101111111111111000000000000000000000000000000000000000000000000000000;
		6249: Delta = 69'sb000000000000110000000000000000000000000000000000000000000000000000000;
		44612: Delta = 69'sb111111111111010000000000000000000000000000000000000000000000000000000;
		10415: Delta = 69'sb000000000001010000000000000000000000000000000000000000000000000000000;
		40446: Delta = 69'sb111111111110110000000000000000000000000000000000000000000000000000000;
		18747: Delta = 69'sb000000000010010000000000000000000000000000000000000000000000000000000;
		36280: Delta = 69'sb111111111110010000000000000000000000000000000000000000000000000000000;
		14581: Delta = 69'sb000000000001110000000000000000000000000000000000000000000000000000000;
		32114: Delta = 69'sb111111111101110000000000000000000000000000000000000000000000000000000;
		35411: Delta = 69'sb000000000100010000000000000000000000000000000000000000000000000000000;
		19616: Delta = 69'sb111111111100010000000000000000000000000000000000000000000000000000000;
		31245: Delta = 69'sb000000000011110000000000000000000000000000000000000000000000000000000;
		15450: Delta = 69'sb111111111011110000000000000000000000000000000000000000000000000000000;
		17878: Delta = 69'sb000000001000010000000000000000000000000000000000000000000000000000000;
		37149: Delta = 69'sb111111111000010000000000000000000000000000000000000000000000000000000;
		13712: Delta = 69'sb000000000111110000000000000000000000000000000000000000000000000000000;
		32983: Delta = 69'sb111111110111110000000000000000000000000000000000000000000000000000000;
		33673: Delta = 69'sb000000010000010000000000000000000000000000000000000000000000000000000;
		21354: Delta = 69'sb111111110000010000000000000000000000000000000000000000000000000000000;
		29507: Delta = 69'sb000000001111110000000000000000000000000000000000000000000000000000000;
		17188: Delta = 69'sb111111101111110000000000000000000000000000000000000000000000000000000;
		14402: Delta = 69'sb000000100000010000000000000000000000000000000000000000000000000000000;
		40625: Delta = 69'sb111111100000010000000000000000000000000000000000000000000000000000000;
		10236: Delta = 69'sb000000011111110000000000000000000000000000000000000000000000000000000;
		36459: Delta = 69'sb111111011111110000000000000000000000000000000000000000000000000000000;
		26721: Delta = 69'sb000001000000010000000000000000000000000000000000000000000000000000000;
		28306: Delta = 69'sb111111000000010000000000000000000000000000000000000000000000000000000;
		22555: Delta = 69'sb000000111111110000000000000000000000000000000000000000000000000000000;
		24140: Delta = 69'sb111110111111110000000000000000000000000000000000000000000000000000000;
		498: Delta = 69'sb000010000000010000000000000000000000000000000000000000000000000000000;
		3668: Delta = 69'sb111110000000010000000000000000000000000000000000000000000000000000000;
		47193: Delta = 69'sb000001111111110000000000000000000000000000000000000000000000000000000;
		50363: Delta = 69'sb111101111111110000000000000000000000000000000000000000000000000000000;
		49774: Delta = 69'sb000100000000010000000000000000000000000000000000000000000000000000000;
		5253: Delta = 69'sb111100000000010000000000000000000000000000000000000000000000000000000;
		45608: Delta = 69'sb000011111111110000000000000000000000000000000000000000000000000000000;
		1087: Delta = 69'sb111011111111110000000000000000000000000000000000000000000000000000000;
		46604: Delta = 69'sb001000000000010000000000000000000000000000000000000000000000000000000;
		8423: Delta = 69'sb111000000000010000000000000000000000000000000000000000000000000000000;
		42438: Delta = 69'sb000111111111110000000000000000000000000000000000000000000000000000000;
		4257: Delta = 69'sb110111111111110000000000000000000000000000000000000000000000000000000;
		40264: Delta = 69'sb010000000000010000000000000000000000000000000000000000000000000000000;
		14763: Delta = 69'sb110000000000010000000000000000000000000000000000000000000000000000000;
		36098: Delta = 69'sb001111111111110000000000000000000000000000000000000000000000000000000;
		10597: Delta = 69'sb101111111111110000000000000000000000000000000000000000000000000000000;
		12498: Delta = 69'sb000000000001100000000000000000000000000000000000000000000000000000000;
		38363: Delta = 69'sb111111111110100000000000000000000000000000000000000000000000000000000;
		20830: Delta = 69'sb000000000010100000000000000000000000000000000000000000000000000000000;
		30031: Delta = 69'sb111111111101100000000000000000000000000000000000000000000000000000000;
		37494: Delta = 69'sb000000000100100000000000000000000000000000000000000000000000000000000;
		21699: Delta = 69'sb111111111100100000000000000000000000000000000000000000000000000000000;
		29162: Delta = 69'sb000000000011100000000000000000000000000000000000000000000000000000000;
		13367: Delta = 69'sb111111111011100000000000000000000000000000000000000000000000000000000;
		19961: Delta = 69'sb000000001000100000000000000000000000000000000000000000000000000000000;
		39232: Delta = 69'sb111111111000100000000000000000000000000000000000000000000000000000000;
		11629: Delta = 69'sb000000000111100000000000000000000000000000000000000000000000000000000;
		30900: Delta = 69'sb111111110111100000000000000000000000000000000000000000000000000000000;
		35756: Delta = 69'sb000000010000100000000000000000000000000000000000000000000000000000000;
		23437: Delta = 69'sb111111110000100000000000000000000000000000000000000000000000000000000;
		27424: Delta = 69'sb000000001111100000000000000000000000000000000000000000000000000000000;
		15105: Delta = 69'sb111111101111100000000000000000000000000000000000000000000000000000000;
		16485: Delta = 69'sb000000100000100000000000000000000000000000000000000000000000000000000;
		42708: Delta = 69'sb111111100000100000000000000000000000000000000000000000000000000000000;
		8153: Delta = 69'sb000000011111100000000000000000000000000000000000000000000000000000000;
		34376: Delta = 69'sb111111011111100000000000000000000000000000000000000000000000000000000;
		28804: Delta = 69'sb000001000000100000000000000000000000000000000000000000000000000000000;
		30389: Delta = 69'sb111111000000100000000000000000000000000000000000000000000000000000000;
		20472: Delta = 69'sb000000111111100000000000000000000000000000000000000000000000000000000;
		22057: Delta = 69'sb111110111111100000000000000000000000000000000000000000000000000000000;
		2581: Delta = 69'sb000010000000100000000000000000000000000000000000000000000000000000000;
		5751: Delta = 69'sb111110000000100000000000000000000000000000000000000000000000000000000;
		45110: Delta = 69'sb000001111111100000000000000000000000000000000000000000000000000000000;
		48280: Delta = 69'sb111101111111100000000000000000000000000000000000000000000000000000000;
		996: Delta = 69'sb000100000000100000000000000000000000000000000000000000000000000000000;
		7336: Delta = 69'sb111100000000100000000000000000000000000000000000000000000000000000000;
		43525: Delta = 69'sb000011111111100000000000000000000000000000000000000000000000000000000;
		49865: Delta = 69'sb111011111111100000000000000000000000000000000000000000000000000000000;
		48687: Delta = 69'sb001000000000100000000000000000000000000000000000000000000000000000000;
		10506: Delta = 69'sb111000000000100000000000000000000000000000000000000000000000000000000;
		40355: Delta = 69'sb000111111111100000000000000000000000000000000000000000000000000000000;
		2174: Delta = 69'sb110111111111100000000000000000000000000000000000000000000000000000000;
		42347: Delta = 69'sb010000000000100000000000000000000000000000000000000000000000000000000;
		16846: Delta = 69'sb110000000000100000000000000000000000000000000000000000000000000000000;
		34015: Delta = 69'sb001111111111100000000000000000000000000000000000000000000000000000000;
		8514: Delta = 69'sb101111111111100000000000000000000000000000000000000000000000000000000;
		24996: Delta = 69'sb000000000011000000000000000000000000000000000000000000000000000000000;
		25865: Delta = 69'sb111111111101000000000000000000000000000000000000000000000000000000000;
		41660: Delta = 69'sb000000000101000000000000000000000000000000000000000000000000000000000;
		9201: Delta = 69'sb111111111011000000000000000000000000000000000000000000000000000000000;
		24127: Delta = 69'sb000000001001000000000000000000000000000000000000000000000000000000000;
		43398: Delta = 69'sb111111111001000000000000000000000000000000000000000000000000000000000;
		7463: Delta = 69'sb000000000111000000000000000000000000000000000000000000000000000000000;
		26734: Delta = 69'sb111111110111000000000000000000000000000000000000000000000000000000000;
		39922: Delta = 69'sb000000010001000000000000000000000000000000000000000000000000000000000;
		27603: Delta = 69'sb111111110001000000000000000000000000000000000000000000000000000000000;
		23258: Delta = 69'sb000000001111000000000000000000000000000000000000000000000000000000000;
		10939: Delta = 69'sb111111101111000000000000000000000000000000000000000000000000000000000;
		20651: Delta = 69'sb000000100001000000000000000000000000000000000000000000000000000000000;
		46874: Delta = 69'sb111111100001000000000000000000000000000000000000000000000000000000000;
		3987: Delta = 69'sb000000011111000000000000000000000000000000000000000000000000000000000;
		30210: Delta = 69'sb111111011111000000000000000000000000000000000000000000000000000000000;
		32970: Delta = 69'sb000001000001000000000000000000000000000000000000000000000000000000000;
		34555: Delta = 69'sb111111000001000000000000000000000000000000000000000000000000000000000;
		16306: Delta = 69'sb000000111111000000000000000000000000000000000000000000000000000000000;
		17891: Delta = 69'sb111110111111000000000000000000000000000000000000000000000000000000000;
		6747: Delta = 69'sb000010000001000000000000000000000000000000000000000000000000000000000;
		9917: Delta = 69'sb111110000001000000000000000000000000000000000000000000000000000000000;
		40944: Delta = 69'sb000001111111000000000000000000000000000000000000000000000000000000000;
		44114: Delta = 69'sb111101111111000000000000000000000000000000000000000000000000000000000;
		5162: Delta = 69'sb000100000001000000000000000000000000000000000000000000000000000000000;
		11502: Delta = 69'sb111100000001000000000000000000000000000000000000000000000000000000000;
		39359: Delta = 69'sb000011111111000000000000000000000000000000000000000000000000000000000;
		45699: Delta = 69'sb111011111111000000000000000000000000000000000000000000000000000000000;
		1992: Delta = 69'sb001000000001000000000000000000000000000000000000000000000000000000000;
		14672: Delta = 69'sb111000000001000000000000000000000000000000000000000000000000000000000;
		36189: Delta = 69'sb000111111111000000000000000000000000000000000000000000000000000000000;
		48869: Delta = 69'sb110111111111000000000000000000000000000000000000000000000000000000000;
		46513: Delta = 69'sb010000000001000000000000000000000000000000000000000000000000000000000;
		21012: Delta = 69'sb110000000001000000000000000000000000000000000000000000000000000000000;
		29849: Delta = 69'sb001111111111000000000000000000000000000000000000000000000000000000000;
		4348: Delta = 69'sb101111111111000000000000000000000000000000000000000000000000000000000;
		49992: Delta = 69'sb000000000110000000000000000000000000000000000000000000000000000000000;
		869: Delta = 69'sb111111111010000000000000000000000000000000000000000000000000000000000;
		32459: Delta = 69'sb000000001010000000000000000000000000000000000000000000000000000000000;
		18402: Delta = 69'sb111111110110000000000000000000000000000000000000000000000000000000000;
		48254: Delta = 69'sb000000010010000000000000000000000000000000000000000000000000000000000;
		35935: Delta = 69'sb111111110010000000000000000000000000000000000000000000000000000000000;
		14926: Delta = 69'sb000000001110000000000000000000000000000000000000000000000000000000000;
		2607: Delta = 69'sb111111101110000000000000000000000000000000000000000000000000000000000;
		28983: Delta = 69'sb000000100010000000000000000000000000000000000000000000000000000000000;
		4345: Delta = 69'sb111111100010000000000000000000000000000000000000000000000000000000000;
		46516: Delta = 69'sb000000011110000000000000000000000000000000000000000000000000000000000;
		21878: Delta = 69'sb111111011110000000000000000000000000000000000000000000000000000000000;
		41302: Delta = 69'sb000001000010000000000000000000000000000000000000000000000000000000000;
		42887: Delta = 69'sb111111000010000000000000000000000000000000000000000000000000000000000;
		7974: Delta = 69'sb000000111110000000000000000000000000000000000000000000000000000000000;
		9559: Delta = 69'sb111110111110000000000000000000000000000000000000000000000000000000000;
		15079: Delta = 69'sb000010000010000000000000000000000000000000000000000000000000000000000;
		18249: Delta = 69'sb111110000010000000000000000000000000000000000000000000000000000000000;
		32612: Delta = 69'sb000001111110000000000000000000000000000000000000000000000000000000000;
		35782: Delta = 69'sb111101111110000000000000000000000000000000000000000000000000000000000;
		13494: Delta = 69'sb000100000010000000000000000000000000000000000000000000000000000000000;
		19834: Delta = 69'sb111100000010000000000000000000000000000000000000000000000000000000000;
		31027: Delta = 69'sb000011111110000000000000000000000000000000000000000000000000000000000;
		37367: Delta = 69'sb111011111110000000000000000000000000000000000000000000000000000000000;
		10324: Delta = 69'sb001000000010000000000000000000000000000000000000000000000000000000000;
		23004: Delta = 69'sb111000000010000000000000000000000000000000000000000000000000000000000;
		27857: Delta = 69'sb000111111110000000000000000000000000000000000000000000000000000000000;
		40537: Delta = 69'sb110111111110000000000000000000000000000000000000000000000000000000000;
		3984: Delta = 69'sb010000000010000000000000000000000000000000000000000000000000000000000;
		29344: Delta = 69'sb110000000010000000000000000000000000000000000000000000000000000000000;
		21517: Delta = 69'sb001111111110000000000000000000000000000000000000000000000000000000000;
		46877: Delta = 69'sb101111111110000000000000000000000000000000000000000000000000000000000;
		49123: Delta = 69'sb000000001100000000000000000000000000000000000000000000000000000000000;
		1738: Delta = 69'sb111111110100000000000000000000000000000000000000000000000000000000000;
		14057: Delta = 69'sb000000010100000000000000000000000000000000000000000000000000000000000;
		36804: Delta = 69'sb111111101100000000000000000000000000000000000000000000000000000000000;
		45647: Delta = 69'sb000000100100000000000000000000000000000000000000000000000000000000000;
		21009: Delta = 69'sb111111100100000000000000000000000000000000000000000000000000000000000;
		29852: Delta = 69'sb000000011100000000000000000000000000000000000000000000000000000000000;
		5214: Delta = 69'sb111111011100000000000000000000000000000000000000000000000000000000000;
		7105: Delta = 69'sb000001000100000000000000000000000000000000000000000000000000000000000;
		8690: Delta = 69'sb111111000100000000000000000000000000000000000000000000000000000000000;
		42171: Delta = 69'sb000000111100000000000000000000000000000000000000000000000000000000000;
		43756: Delta = 69'sb111110111100000000000000000000000000000000000000000000000000000000000;
		31743: Delta = 69'sb000010000100000000000000000000000000000000000000000000000000000000000;
		34913: Delta = 69'sb111110000100000000000000000000000000000000000000000000000000000000000;
		15948: Delta = 69'sb000001111100000000000000000000000000000000000000000000000000000000000;
		19118: Delta = 69'sb111101111100000000000000000000000000000000000000000000000000000000000;
		30158: Delta = 69'sb000100000100000000000000000000000000000000000000000000000000000000000;
		36498: Delta = 69'sb111100000100000000000000000000000000000000000000000000000000000000000;
		14363: Delta = 69'sb000011111100000000000000000000000000000000000000000000000000000000000;
		20703: Delta = 69'sb111011111100000000000000000000000000000000000000000000000000000000000;
		26988: Delta = 69'sb001000000100000000000000000000000000000000000000000000000000000000000;
		39668: Delta = 69'sb111000000100000000000000000000000000000000000000000000000000000000000;
		11193: Delta = 69'sb000111111100000000000000000000000000000000000000000000000000000000000;
		23873: Delta = 69'sb110111111100000000000000000000000000000000000000000000000000000000000;
		20648: Delta = 69'sb010000000100000000000000000000000000000000000000000000000000000000000;
		46008: Delta = 69'sb110000000100000000000000000000000000000000000000000000000000000000000;
		4853: Delta = 69'sb001111111100000000000000000000000000000000000000000000000000000000000;
		30213: Delta = 69'sb101111111100000000000000000000000000000000000000000000000000000000000;
		47385: Delta = 69'sb000000011000000000000000000000000000000000000000000000000000000000000;
		3476: Delta = 69'sb111111101000000000000000000000000000000000000000000000000000000000000;
		28114: Delta = 69'sb000000101000000000000000000000000000000000000000000000000000000000000;
		22747: Delta = 69'sb111111011000000000000000000000000000000000000000000000000000000000000;
		40433: Delta = 69'sb000001001000000000000000000000000000000000000000000000000000000000000;
		42018: Delta = 69'sb111111001000000000000000000000000000000000000000000000000000000000000;
		8843: Delta = 69'sb000000111000000000000000000000000000000000000000000000000000000000000;
		10428: Delta = 69'sb111110111000000000000000000000000000000000000000000000000000000000000;
		14210: Delta = 69'sb000010001000000000000000000000000000000000000000000000000000000000000;
		17380: Delta = 69'sb111110001000000000000000000000000000000000000000000000000000000000000;
		33481: Delta = 69'sb000001111000000000000000000000000000000000000000000000000000000000000;
		36651: Delta = 69'sb111101111000000000000000000000000000000000000000000000000000000000000;
		12625: Delta = 69'sb000100001000000000000000000000000000000000000000000000000000000000000;
		18965: Delta = 69'sb111100001000000000000000000000000000000000000000000000000000000000000;
		31896: Delta = 69'sb000011111000000000000000000000000000000000000000000000000000000000000;
		38236: Delta = 69'sb111011111000000000000000000000000000000000000000000000000000000000000;
		9455: Delta = 69'sb001000001000000000000000000000000000000000000000000000000000000000000;
		22135: Delta = 69'sb111000001000000000000000000000000000000000000000000000000000000000000;
		28726: Delta = 69'sb000111111000000000000000000000000000000000000000000000000000000000000;
		41406: Delta = 69'sb110111111000000000000000000000000000000000000000000000000000000000000;
		3115: Delta = 69'sb010000001000000000000000000000000000000000000000000000000000000000000;
		28475: Delta = 69'sb110000001000000000000000000000000000000000000000000000000000000000000;
		22386: Delta = 69'sb001111111000000000000000000000000000000000000000000000000000000000000;
		47746: Delta = 69'sb101111111000000000000000000000000000000000000000000000000000000000000;
		43909: Delta = 69'sb000000110000000000000000000000000000000000000000000000000000000000000;
		6952: Delta = 69'sb111111010000000000000000000000000000000000000000000000000000000000000;
		5367: Delta = 69'sb000001010000000000000000000000000000000000000000000000000000000000000;
		45494: Delta = 69'sb111110110000000000000000000000000000000000000000000000000000000000000;
		30005: Delta = 69'sb000010010000000000000000000000000000000000000000000000000000000000000;
		33175: Delta = 69'sb111110010000000000000000000000000000000000000000000000000000000000000;
		17686: Delta = 69'sb000001110000000000000000000000000000000000000000000000000000000000000;
		20856: Delta = 69'sb111101110000000000000000000000000000000000000000000000000000000000000;
		28420: Delta = 69'sb000100010000000000000000000000000000000000000000000000000000000000000;
		34760: Delta = 69'sb111100010000000000000000000000000000000000000000000000000000000000000;
		16101: Delta = 69'sb000011110000000000000000000000000000000000000000000000000000000000000;
		22441: Delta = 69'sb111011110000000000000000000000000000000000000000000000000000000000000;
		25250: Delta = 69'sb001000010000000000000000000000000000000000000000000000000000000000000;
		37930: Delta = 69'sb111000010000000000000000000000000000000000000000000000000000000000000;
		12931: Delta = 69'sb000111110000000000000000000000000000000000000000000000000000000000000;
		25611: Delta = 69'sb110111110000000000000000000000000000000000000000000000000000000000000;
		18910: Delta = 69'sb010000010000000000000000000000000000000000000000000000000000000000000;
		44270: Delta = 69'sb110000010000000000000000000000000000000000000000000000000000000000000;
		6591: Delta = 69'sb001111110000000000000000000000000000000000000000000000000000000000000;
		31951: Delta = 69'sb101111110000000000000000000000000000000000000000000000000000000000000;
		36957: Delta = 69'sb000001100000000000000000000000000000000000000000000000000000000000000;
		13904: Delta = 69'sb111110100000000000000000000000000000000000000000000000000000000000000;
		10734: Delta = 69'sb000010100000000000000000000000000000000000000000000000000000000000000;
		40127: Delta = 69'sb111101100000000000000000000000000000000000000000000000000000000000000;
		9149: Delta = 69'sb000100100000000000000000000000000000000000000000000000000000000000000;
		15489: Delta = 69'sb111100100000000000000000000000000000000000000000000000000000000000000;
		35372: Delta = 69'sb000011100000000000000000000000000000000000000000000000000000000000000;
		41712: Delta = 69'sb111011100000000000000000000000000000000000000000000000000000000000000;
		5979: Delta = 69'sb001000100000000000000000000000000000000000000000000000000000000000000;
		18659: Delta = 69'sb111000100000000000000000000000000000000000000000000000000000000000000;
		32202: Delta = 69'sb000111100000000000000000000000000000000000000000000000000000000000000;
		44882: Delta = 69'sb110111100000000000000000000000000000000000000000000000000000000000000;
		50500: Delta = 69'sb010000100000000000000000000000000000000000000000000000000000000000000;
		24999: Delta = 69'sb110000100000000000000000000000000000000000000000000000000000000000000;
		25862: Delta = 69'sb001111100000000000000000000000000000000000000000000000000000000000000;
		361: Delta = 69'sb101111100000000000000000000000000000000000000000000000000000000000000;
		23053: Delta = 69'sb000011000000000000000000000000000000000000000000000000000000000000000;
		27808: Delta = 69'sb111101000000000000000000000000000000000000000000000000000000000000000;
		21468: Delta = 69'sb000101000000000000000000000000000000000000000000000000000000000000000;
		29393: Delta = 69'sb111011000000000000000000000000000000000000000000000000000000000000000;
		18298: Delta = 69'sb001001000000000000000000000000000000000000000000000000000000000000000;
		30978: Delta = 69'sb111001000000000000000000000000000000000000000000000000000000000000000;
		19883: Delta = 69'sb000111000000000000000000000000000000000000000000000000000000000000000;
		32563: Delta = 69'sb110111000000000000000000000000000000000000000000000000000000000000000;
		11958: Delta = 69'sb010001000000000000000000000000000000000000000000000000000000000000000;
		37318: Delta = 69'sb110001000000000000000000000000000000000000000000000000000000000000000;
		13543: Delta = 69'sb001111000000000000000000000000000000000000000000000000000000000000000;
		38903: Delta = 69'sb101111000000000000000000000000000000000000000000000000000000000000000;
		46106: Delta = 69'sb000110000000000000000000000000000000000000000000000000000000000000000;
		4755: Delta = 69'sb111010000000000000000000000000000000000000000000000000000000000000000;
		42936: Delta = 69'sb001010000000000000000000000000000000000000000000000000000000000000000;
		7925: Delta = 69'sb110110000000000000000000000000000000000000000000000000000000000000000;
		36596: Delta = 69'sb010010000000000000000000000000000000000000000000000000000000000000000;
		11095: Delta = 69'sb110010000000000000000000000000000000000000000000000000000000000000000;
		39766: Delta = 69'sb001110000000000000000000000000000000000000000000000000000000000000000;
		14265: Delta = 69'sb101110000000000000000000000000000000000000000000000000000000000000000;
		41351: Delta = 69'sb001100000000000000000000000000000000000000000000000000000000000000000;
		9510: Delta = 69'sb110100000000000000000000000000000000000000000000000000000000000000000;
		35011: Delta = 69'sb010100000000000000000000000000000000000000000000000000000000000000000;
		15850: Delta = 69'sb101100000000000000000000000000000000000000000000000000000000000000000;
		31841: Delta = 69'sb011000000000000000000000000000000000000000000000000000000000000000000;
		19020: Delta = 69'sb101000000000000000000000000000000000000000000000000000000000000000000;
		default: Delta =69'sb0;
	endcase
end

wire signed [W_BITS-1:0] W_signed;
assign W_signed = (W - Delta);

always@(posedge clk or negedge rst_n) begin
   if(!rst_n) begin
     	ps <= idle;
    end
   else begin
        case(ps)
            idle: begin
                found <= 0;
                R <= 0;
        	Q <= 0;
                ps <= pre;
                end
	    pre: begin
		 Q <= W / A;
		 ps <= load;
		end
            load: begin
                 R <= W - (A * Q);
		 ps <= LUT;
		end
	    LUT: begin
		  if(Delta != 0)begin
		      N <= W_signed / A ;	
		      found <= 1;
                      ps <= idle;
		  end
		  else begin
		      N <= Q;
		      found <= 1;
                      ps <= idle;
		  end
		end
	endcase
    end
end

endmodule

// Product (AN) Code DEC_LUT_Decoder
// DEC_LUT_Decoder16bits.v
// Received codeword W = AN + E, E is double AWE (E = e1 + e2), +2^i or -2^i.
module DEC_LUT_Decoder16bits_clk(clk, rst_n, W, found, N);

//=========================================================================
//   PARAMETER AND LOCALPARAM FOR FSM
//   W_BITS 要考慮 OVERFLOW 問題
//   N_BITS 也要考慮 OVERFLOW 問題
//=========================================================================
parameter A = 4547 , W_BITS = 30, A_BITS = 13 , N_BITS = 17;

localparam [1:0] idle=2'b00, pre=2'b01,load=2'b10, LUT=2'b11;

reg [1:0] ps;
//==========================================
//   INPUT AND OUTPUT DECLARATION
//==========================================
input   clk, rst_n;
input 	[W_BITS-1:0]	W;
output	reg  [N_BITS-1:0] N;
output  reg  found;

reg 	[N_BITS-1:0]	Q;
reg 	[A_BITS-1:0]	R;


reg	signed	[29:0]	Delta;
always@(*) begin
	case(R)
		1: Delta = 30'sb000000000000000000000000000001;
		4546: Delta = 30'sb111111111111111111111111111111;
		2: Delta = 30'sb000000000000000000000000000010;
		4545: Delta = 30'sb111111111111111111111111111110;
		4: Delta = 30'sb000000000000000000000000000100;
		4543: Delta = 30'sb111111111111111111111111111100;
		8: Delta = 30'sb000000000000000000000000001000;
		4539: Delta = 30'sb111111111111111111111111111000;
		16: Delta = 30'sb000000000000000000000000010000;
		4531: Delta = 30'sb111111111111111111111111110000;
		32: Delta = 30'sb000000000000000000000000100000;
		4515: Delta = 30'sb111111111111111111111111100000;
		64: Delta = 30'sb000000000000000000000001000000;
		4483: Delta = 30'sb111111111111111111111111000000;
		128: Delta = 30'sb000000000000000000000010000000;
		4419: Delta = 30'sb111111111111111111111110000000;
		256: Delta = 30'sb000000000000000000000100000000;
		4291: Delta = 30'sb111111111111111111111100000000;
		512: Delta = 30'sb000000000000000000001000000000;
		4035: Delta = 30'sb111111111111111111111000000000;
		1024: Delta = 30'sb000000000000000000010000000000;
		3523: Delta = 30'sb111111111111111111110000000000;
		2048: Delta = 30'sb000000000000000000100000000000;
		2499: Delta = 30'sb111111111111111111100000000000;
		4096: Delta = 30'sb000000000000000001000000000000;
		451: Delta = 30'sb111111111111111111000000000000;
		3645: Delta = 30'sb000000000000000010000000000000;
		902: Delta = 30'sb111111111111111110000000000000;
		2743: Delta = 30'sb000000000000000100000000000000;
		1804: Delta = 30'sb111111111111111100000000000000;
		939: Delta = 30'sb000000000000001000000000000000;
		3608: Delta = 30'sb111111111111111000000000000000;
		1878: Delta = 30'sb000000000000010000000000000000;
		2669: Delta = 30'sb111111111111110000000000000000;
		3756: Delta = 30'sb000000000000100000000000000000;
		791: Delta = 30'sb111111111111100000000000000000;
		2965: Delta = 30'sb000000000001000000000000000000;
		1582: Delta = 30'sb111111111111000000000000000000;
		1383: Delta = 30'sb000000000010000000000000000000;
		3164: Delta = 30'sb111111111110000000000000000000;
		2766: Delta = 30'sb000000000100000000000000000000;
		1781: Delta = 30'sb111111111100000000000000000000;
		985: Delta = 30'sb000000001000000000000000000000;
		3562: Delta = 30'sb111111111000000000000000000000;
		1970: Delta = 30'sb000000010000000000000000000000;
		2577: Delta = 30'sb111111110000000000000000000000;
		3940: Delta = 30'sb000000100000000000000000000000;
		607: Delta = 30'sb111111100000000000000000000000;
		3333: Delta = 30'sb000001000000000000000000000000;
		1214: Delta = 30'sb111111000000000000000000000000;
		2119: Delta = 30'sb000010000000000000000000000000;
		2428: Delta = 30'sb111110000000000000000000000000;
		4238: Delta = 30'sb000100000000000000000000000000;
		309: Delta = 30'sb111100000000000000000000000000;
		3929: Delta = 30'sb001000000000000000000000000000;
		618: Delta = 30'sb111000000000000000000000000000;
		3311: Delta = 30'sb010000000000000000000000000000;
		1236: Delta = 30'sb110000000000000000000000000000;
		3: Delta = 30'sb000000000000000000000000000011;
		4544: Delta = 30'sb111111111111111111111111111101;
		5: Delta = 30'sb000000000000000000000000000101;
		4542: Delta = 30'sb111111111111111111111111111011;
		9: Delta = 30'sb000000000000000000000000001001;
		4540: Delta = 30'sb111111111111111111111111111001;
		7: Delta = 30'sb000000000000000000000000000111;
		4538: Delta = 30'sb111111111111111111111111110111;
		17: Delta = 30'sb000000000000000000000000010001;
		4532: Delta = 30'sb111111111111111111111111110001;
		15: Delta = 30'sb000000000000000000000000001111;
		4530: Delta = 30'sb111111111111111111111111101111;
		33: Delta = 30'sb000000000000000000000000100001;
		4516: Delta = 30'sb111111111111111111111111100001;
		31: Delta = 30'sb000000000000000000000000011111;
		4514: Delta = 30'sb111111111111111111111111011111;
		65: Delta = 30'sb000000000000000000000001000001;
		4484: Delta = 30'sb111111111111111111111111000001;
		63: Delta = 30'sb000000000000000000000000111111;
		4482: Delta = 30'sb111111111111111111111110111111;
		129: Delta = 30'sb000000000000000000000010000001;
		4420: Delta = 30'sb111111111111111111111110000001;
		127: Delta = 30'sb000000000000000000000001111111;
		4418: Delta = 30'sb111111111111111111111101111111;
		257: Delta = 30'sb000000000000000000000100000001;
		4292: Delta = 30'sb111111111111111111111100000001;
		255: Delta = 30'sb000000000000000000000011111111;
		4290: Delta = 30'sb111111111111111111111011111111;
		513: Delta = 30'sb000000000000000000001000000001;
		4036: Delta = 30'sb111111111111111111111000000001;
		511: Delta = 30'sb000000000000000000000111111111;
		4034: Delta = 30'sb111111111111111111110111111111;
		1025: Delta = 30'sb000000000000000000010000000001;
		3524: Delta = 30'sb111111111111111111110000000001;
		1023: Delta = 30'sb000000000000000000001111111111;
		3522: Delta = 30'sb111111111111111111101111111111;
		2049: Delta = 30'sb000000000000000000100000000001;
		2500: Delta = 30'sb111111111111111111100000000001;
		2047: Delta = 30'sb000000000000000000011111111111;
		2498: Delta = 30'sb111111111111111111011111111111;
		4097: Delta = 30'sb000000000000000001000000000001;
		452: Delta = 30'sb111111111111111111000000000001;
		4095: Delta = 30'sb000000000000000000111111111111;
		450: Delta = 30'sb111111111111111110111111111111;
		3646: Delta = 30'sb000000000000000010000000000001;
		903: Delta = 30'sb111111111111111110000000000001;
		3644: Delta = 30'sb000000000000000001111111111111;
		901: Delta = 30'sb111111111111111101111111111111;
		2744: Delta = 30'sb000000000000000100000000000001;
		1805: Delta = 30'sb111111111111111100000000000001;
		2742: Delta = 30'sb000000000000000011111111111111;
		1803: Delta = 30'sb111111111111111011111111111111;
		940: Delta = 30'sb000000000000001000000000000001;
		3609: Delta = 30'sb111111111111111000000000000001;
		938: Delta = 30'sb000000000000000111111111111111;
		3607: Delta = 30'sb111111111111110111111111111111;
		1879: Delta = 30'sb000000000000010000000000000001;
		2670: Delta = 30'sb111111111111110000000000000001;
		1877: Delta = 30'sb000000000000001111111111111111;
		2668: Delta = 30'sb111111111111101111111111111111;
		3757: Delta = 30'sb000000000000100000000000000001;
		792: Delta = 30'sb111111111111100000000000000001;
		3755: Delta = 30'sb000000000000011111111111111111;
		790: Delta = 30'sb111111111111011111111111111111;
		2966: Delta = 30'sb000000000001000000000000000001;
		1583: Delta = 30'sb111111111111000000000000000001;
		2964: Delta = 30'sb000000000000111111111111111111;
		1581: Delta = 30'sb111111111110111111111111111111;
		1384: Delta = 30'sb000000000010000000000000000001;
		3165: Delta = 30'sb111111111110000000000000000001;
		1382: Delta = 30'sb000000000001111111111111111111;
		3163: Delta = 30'sb111111111101111111111111111111;
		2767: Delta = 30'sb000000000100000000000000000001;
		1782: Delta = 30'sb111111111100000000000000000001;
		2765: Delta = 30'sb000000000011111111111111111111;
		1780: Delta = 30'sb111111111011111111111111111111;
		986: Delta = 30'sb000000001000000000000000000001;
		3563: Delta = 30'sb111111111000000000000000000001;
		984: Delta = 30'sb000000000111111111111111111111;
		3561: Delta = 30'sb111111110111111111111111111111;
		1971: Delta = 30'sb000000010000000000000000000001;
		2578: Delta = 30'sb111111110000000000000000000001;
		1969: Delta = 30'sb000000001111111111111111111111;
		2576: Delta = 30'sb111111101111111111111111111111;
		3941: Delta = 30'sb000000100000000000000000000001;
		608: Delta = 30'sb111111100000000000000000000001;
		3939: Delta = 30'sb000000011111111111111111111111;
		606: Delta = 30'sb111111011111111111111111111111;
		3334: Delta = 30'sb000001000000000000000000000001;
		1215: Delta = 30'sb111111000000000000000000000001;
		3332: Delta = 30'sb000000111111111111111111111111;
		1213: Delta = 30'sb111110111111111111111111111111;
		2120: Delta = 30'sb000010000000000000000000000001;
		2429: Delta = 30'sb111110000000000000000000000001;
		2118: Delta = 30'sb000001111111111111111111111111;
		2427: Delta = 30'sb111101111111111111111111111111;
		4239: Delta = 30'sb000100000000000000000000000001;
		310: Delta = 30'sb111100000000000000000000000001;
		4237: Delta = 30'sb000011111111111111111111111111;
		308: Delta = 30'sb111011111111111111111111111111;
		3930: Delta = 30'sb001000000000000000000000000001;
		619: Delta = 30'sb111000000000000000000000000001;
		3928: Delta = 30'sb000111111111111111111111111111;
		617: Delta = 30'sb110111111111111111111111111111;
		3312: Delta = 30'sb010000000000000000000000000001;
		1237: Delta = 30'sb110000000000000000000000000001;
		3310: Delta = 30'sb001111111111111111111111111111;
		1235: Delta = 30'sb101111111111111111111111111111;
		6: Delta = 30'sb000000000000000000000000000110;
		4541: Delta = 30'sb111111111111111111111111111010;
		10: Delta = 30'sb000000000000000000000000001010;
		4537: Delta = 30'sb111111111111111111111111110110;
		18: Delta = 30'sb000000000000000000000000010010;
		4533: Delta = 30'sb111111111111111111111111110010;
		14: Delta = 30'sb000000000000000000000000001110;
		4529: Delta = 30'sb111111111111111111111111101110;
		34: Delta = 30'sb000000000000000000000000100010;
		4517: Delta = 30'sb111111111111111111111111100010;
		30: Delta = 30'sb000000000000000000000000011110;
		4513: Delta = 30'sb111111111111111111111111011110;
		66: Delta = 30'sb000000000000000000000001000010;
		4485: Delta = 30'sb111111111111111111111111000010;
		62: Delta = 30'sb000000000000000000000000111110;
		4481: Delta = 30'sb111111111111111111111110111110;
		130: Delta = 30'sb000000000000000000000010000010;
		4421: Delta = 30'sb111111111111111111111110000010;
		126: Delta = 30'sb000000000000000000000001111110;
		4417: Delta = 30'sb111111111111111111111101111110;
		258: Delta = 30'sb000000000000000000000100000010;
		4293: Delta = 30'sb111111111111111111111100000010;
		254: Delta = 30'sb000000000000000000000011111110;
		4289: Delta = 30'sb111111111111111111111011111110;
		514: Delta = 30'sb000000000000000000001000000010;
		4037: Delta = 30'sb111111111111111111111000000010;
		510: Delta = 30'sb000000000000000000000111111110;
		4033: Delta = 30'sb111111111111111111110111111110;
		1026: Delta = 30'sb000000000000000000010000000010;
		3525: Delta = 30'sb111111111111111111110000000010;
		1022: Delta = 30'sb000000000000000000001111111110;
		3521: Delta = 30'sb111111111111111111101111111110;
		2050: Delta = 30'sb000000000000000000100000000010;
		2501: Delta = 30'sb111111111111111111100000000010;
		2046: Delta = 30'sb000000000000000000011111111110;
		2497: Delta = 30'sb111111111111111111011111111110;
		4098: Delta = 30'sb000000000000000001000000000010;
		453: Delta = 30'sb111111111111111111000000000010;
		4094: Delta = 30'sb000000000000000000111111111110;
		449: Delta = 30'sb111111111111111110111111111110;
		3647: Delta = 30'sb000000000000000010000000000010;
		904: Delta = 30'sb111111111111111110000000000010;
		3643: Delta = 30'sb000000000000000001111111111110;
		900: Delta = 30'sb111111111111111101111111111110;
		2745: Delta = 30'sb000000000000000100000000000010;
		1806: Delta = 30'sb111111111111111100000000000010;
		2741: Delta = 30'sb000000000000000011111111111110;
		1802: Delta = 30'sb111111111111111011111111111110;
		941: Delta = 30'sb000000000000001000000000000010;
		3610: Delta = 30'sb111111111111111000000000000010;
		937: Delta = 30'sb000000000000000111111111111110;
		3606: Delta = 30'sb111111111111110111111111111110;
		1880: Delta = 30'sb000000000000010000000000000010;
		2671: Delta = 30'sb111111111111110000000000000010;
		1876: Delta = 30'sb000000000000001111111111111110;
		2667: Delta = 30'sb111111111111101111111111111110;
		3758: Delta = 30'sb000000000000100000000000000010;
		793: Delta = 30'sb111111111111100000000000000010;
		3754: Delta = 30'sb000000000000011111111111111110;
		789: Delta = 30'sb111111111111011111111111111110;
		2967: Delta = 30'sb000000000001000000000000000010;
		1584: Delta = 30'sb111111111111000000000000000010;
		2963: Delta = 30'sb000000000000111111111111111110;
		1580: Delta = 30'sb111111111110111111111111111110;
		1385: Delta = 30'sb000000000010000000000000000010;
		3166: Delta = 30'sb111111111110000000000000000010;
		1381: Delta = 30'sb000000000001111111111111111110;
		3162: Delta = 30'sb111111111101111111111111111110;
		2768: Delta = 30'sb000000000100000000000000000010;
		1783: Delta = 30'sb111111111100000000000000000010;
		2764: Delta = 30'sb000000000011111111111111111110;
		1779: Delta = 30'sb111111111011111111111111111110;
		987: Delta = 30'sb000000001000000000000000000010;
		3564: Delta = 30'sb111111111000000000000000000010;
		983: Delta = 30'sb000000000111111111111111111110;
		3560: Delta = 30'sb111111110111111111111111111110;
		1972: Delta = 30'sb000000010000000000000000000010;
		2579: Delta = 30'sb111111110000000000000000000010;
		1968: Delta = 30'sb000000001111111111111111111110;
		2575: Delta = 30'sb111111101111111111111111111110;
		3942: Delta = 30'sb000000100000000000000000000010;
		609: Delta = 30'sb111111100000000000000000000010;
		3938: Delta = 30'sb000000011111111111111111111110;
		605: Delta = 30'sb111111011111111111111111111110;
		3335: Delta = 30'sb000001000000000000000000000010;
		1216: Delta = 30'sb111111000000000000000000000010;
		3331: Delta = 30'sb000000111111111111111111111110;
		1212: Delta = 30'sb111110111111111111111111111110;
		2121: Delta = 30'sb000010000000000000000000000010;
		2430: Delta = 30'sb111110000000000000000000000010;
		2117: Delta = 30'sb000001111111111111111111111110;
		2426: Delta = 30'sb111101111111111111111111111110;
		4240: Delta = 30'sb000100000000000000000000000010;
		311: Delta = 30'sb111100000000000000000000000010;
		4236: Delta = 30'sb000011111111111111111111111110;
		307: Delta = 30'sb111011111111111111111111111110;
		3931: Delta = 30'sb001000000000000000000000000010;
		620: Delta = 30'sb111000000000000000000000000010;
		3927: Delta = 30'sb000111111111111111111111111110;
		616: Delta = 30'sb110111111111111111111111111110;
		3313: Delta = 30'sb010000000000000000000000000010;
		1238: Delta = 30'sb110000000000000000000000000010;
		3309: Delta = 30'sb001111111111111111111111111110;
		1234: Delta = 30'sb101111111111111111111111111110;
		12: Delta = 30'sb000000000000000000000000001100;
		4535: Delta = 30'sb111111111111111111111111110100;
		20: Delta = 30'sb000000000000000000000000010100;
		4527: Delta = 30'sb111111111111111111111111101100;
		36: Delta = 30'sb000000000000000000000000100100;
		4519: Delta = 30'sb111111111111111111111111100100;
		28: Delta = 30'sb000000000000000000000000011100;
		4511: Delta = 30'sb111111111111111111111111011100;
		68: Delta = 30'sb000000000000000000000001000100;
		4487: Delta = 30'sb111111111111111111111111000100;
		60: Delta = 30'sb000000000000000000000000111100;
		4479: Delta = 30'sb111111111111111111111110111100;
		132: Delta = 30'sb000000000000000000000010000100;
		4423: Delta = 30'sb111111111111111111111110000100;
		124: Delta = 30'sb000000000000000000000001111100;
		4415: Delta = 30'sb111111111111111111111101111100;
		260: Delta = 30'sb000000000000000000000100000100;
		4295: Delta = 30'sb111111111111111111111100000100;
		252: Delta = 30'sb000000000000000000000011111100;
		4287: Delta = 30'sb111111111111111111111011111100;
		516: Delta = 30'sb000000000000000000001000000100;
		4039: Delta = 30'sb111111111111111111111000000100;
		508: Delta = 30'sb000000000000000000000111111100;
		4031: Delta = 30'sb111111111111111111110111111100;
		1028: Delta = 30'sb000000000000000000010000000100;
		3527: Delta = 30'sb111111111111111111110000000100;
		1020: Delta = 30'sb000000000000000000001111111100;
		3519: Delta = 30'sb111111111111111111101111111100;
		2052: Delta = 30'sb000000000000000000100000000100;
		2503: Delta = 30'sb111111111111111111100000000100;
		2044: Delta = 30'sb000000000000000000011111111100;
		2495: Delta = 30'sb111111111111111111011111111100;
		4100: Delta = 30'sb000000000000000001000000000100;
		455: Delta = 30'sb111111111111111111000000000100;
		4092: Delta = 30'sb000000000000000000111111111100;
		447: Delta = 30'sb111111111111111110111111111100;
		3649: Delta = 30'sb000000000000000010000000000100;
		906: Delta = 30'sb111111111111111110000000000100;
		3641: Delta = 30'sb000000000000000001111111111100;
		898: Delta = 30'sb111111111111111101111111111100;
		2747: Delta = 30'sb000000000000000100000000000100;
		1808: Delta = 30'sb111111111111111100000000000100;
		2739: Delta = 30'sb000000000000000011111111111100;
		1800: Delta = 30'sb111111111111111011111111111100;
		943: Delta = 30'sb000000000000001000000000000100;
		3612: Delta = 30'sb111111111111111000000000000100;
		935: Delta = 30'sb000000000000000111111111111100;
		3604: Delta = 30'sb111111111111110111111111111100;
		1882: Delta = 30'sb000000000000010000000000000100;
		2673: Delta = 30'sb111111111111110000000000000100;
		1874: Delta = 30'sb000000000000001111111111111100;
		2665: Delta = 30'sb111111111111101111111111111100;
		3760: Delta = 30'sb000000000000100000000000000100;
		795: Delta = 30'sb111111111111100000000000000100;
		3752: Delta = 30'sb000000000000011111111111111100;
		787: Delta = 30'sb111111111111011111111111111100;
		2969: Delta = 30'sb000000000001000000000000000100;
		1586: Delta = 30'sb111111111111000000000000000100;
		2961: Delta = 30'sb000000000000111111111111111100;
		1578: Delta = 30'sb111111111110111111111111111100;
		1387: Delta = 30'sb000000000010000000000000000100;
		3168: Delta = 30'sb111111111110000000000000000100;
		1379: Delta = 30'sb000000000001111111111111111100;
		3160: Delta = 30'sb111111111101111111111111111100;
		2770: Delta = 30'sb000000000100000000000000000100;
		1785: Delta = 30'sb111111111100000000000000000100;
		2762: Delta = 30'sb000000000011111111111111111100;
		1777: Delta = 30'sb111111111011111111111111111100;
		989: Delta = 30'sb000000001000000000000000000100;
		3566: Delta = 30'sb111111111000000000000000000100;
		981: Delta = 30'sb000000000111111111111111111100;
		3558: Delta = 30'sb111111110111111111111111111100;
		1974: Delta = 30'sb000000010000000000000000000100;
		2581: Delta = 30'sb111111110000000000000000000100;
		1966: Delta = 30'sb000000001111111111111111111100;
		2573: Delta = 30'sb111111101111111111111111111100;
		3944: Delta = 30'sb000000100000000000000000000100;
		611: Delta = 30'sb111111100000000000000000000100;
		3936: Delta = 30'sb000000011111111111111111111100;
		603: Delta = 30'sb111111011111111111111111111100;
		3337: Delta = 30'sb000001000000000000000000000100;
		1218: Delta = 30'sb111111000000000000000000000100;
		3329: Delta = 30'sb000000111111111111111111111100;
		1210: Delta = 30'sb111110111111111111111111111100;
		2123: Delta = 30'sb000010000000000000000000000100;
		2432: Delta = 30'sb111110000000000000000000000100;
		2115: Delta = 30'sb000001111111111111111111111100;
		2424: Delta = 30'sb111101111111111111111111111100;
		4242: Delta = 30'sb000100000000000000000000000100;
		313: Delta = 30'sb111100000000000000000000000100;
		4234: Delta = 30'sb000011111111111111111111111100;
		305: Delta = 30'sb111011111111111111111111111100;
		3933: Delta = 30'sb001000000000000000000000000100;
		622: Delta = 30'sb111000000000000000000000000100;
		3925: Delta = 30'sb000111111111111111111111111100;
		614: Delta = 30'sb110111111111111111111111111100;
		3315: Delta = 30'sb010000000000000000000000000100;
		1240: Delta = 30'sb110000000000000000000000000100;
		3307: Delta = 30'sb001111111111111111111111111100;
		1232: Delta = 30'sb101111111111111111111111111100;
		24: Delta = 30'sb000000000000000000000000011000;
		4523: Delta = 30'sb111111111111111111111111101000;
		40: Delta = 30'sb000000000000000000000000101000;
		4507: Delta = 30'sb111111111111111111111111011000;
		72: Delta = 30'sb000000000000000000000001001000;
		4491: Delta = 30'sb111111111111111111111111001000;
		56: Delta = 30'sb000000000000000000000000111000;
		4475: Delta = 30'sb111111111111111111111110111000;
		136: Delta = 30'sb000000000000000000000010001000;
		4427: Delta = 30'sb111111111111111111111110001000;
		120: Delta = 30'sb000000000000000000000001111000;
		4411: Delta = 30'sb111111111111111111111101111000;
		264: Delta = 30'sb000000000000000000000100001000;
		4299: Delta = 30'sb111111111111111111111100001000;
		248: Delta = 30'sb000000000000000000000011111000;
		4283: Delta = 30'sb111111111111111111111011111000;
		520: Delta = 30'sb000000000000000000001000001000;
		4043: Delta = 30'sb111111111111111111111000001000;
		504: Delta = 30'sb000000000000000000000111111000;
		4027: Delta = 30'sb111111111111111111110111111000;
		1032: Delta = 30'sb000000000000000000010000001000;
		3531: Delta = 30'sb111111111111111111110000001000;
		1016: Delta = 30'sb000000000000000000001111111000;
		3515: Delta = 30'sb111111111111111111101111111000;
		2056: Delta = 30'sb000000000000000000100000001000;
		2507: Delta = 30'sb111111111111111111100000001000;
		2040: Delta = 30'sb000000000000000000011111111000;
		2491: Delta = 30'sb111111111111111111011111111000;
		4104: Delta = 30'sb000000000000000001000000001000;
		459: Delta = 30'sb111111111111111111000000001000;
		4088: Delta = 30'sb000000000000000000111111111000;
		443: Delta = 30'sb111111111111111110111111111000;
		3653: Delta = 30'sb000000000000000010000000001000;
		910: Delta = 30'sb111111111111111110000000001000;
		3637: Delta = 30'sb000000000000000001111111111000;
		894: Delta = 30'sb111111111111111101111111111000;
		2751: Delta = 30'sb000000000000000100000000001000;
		1812: Delta = 30'sb111111111111111100000000001000;
		2735: Delta = 30'sb000000000000000011111111111000;
		1796: Delta = 30'sb111111111111111011111111111000;
		947: Delta = 30'sb000000000000001000000000001000;
		3616: Delta = 30'sb111111111111111000000000001000;
		931: Delta = 30'sb000000000000000111111111111000;
		3600: Delta = 30'sb111111111111110111111111111000;
		1886: Delta = 30'sb000000000000010000000000001000;
		2677: Delta = 30'sb111111111111110000000000001000;
		1870: Delta = 30'sb000000000000001111111111111000;
		2661: Delta = 30'sb111111111111101111111111111000;
		3764: Delta = 30'sb000000000000100000000000001000;
		799: Delta = 30'sb111111111111100000000000001000;
		3748: Delta = 30'sb000000000000011111111111111000;
		783: Delta = 30'sb111111111111011111111111111000;
		2973: Delta = 30'sb000000000001000000000000001000;
		1590: Delta = 30'sb111111111111000000000000001000;
		2957: Delta = 30'sb000000000000111111111111111000;
		1574: Delta = 30'sb111111111110111111111111111000;
		1391: Delta = 30'sb000000000010000000000000001000;
		3172: Delta = 30'sb111111111110000000000000001000;
		1375: Delta = 30'sb000000000001111111111111111000;
		3156: Delta = 30'sb111111111101111111111111111000;
		2774: Delta = 30'sb000000000100000000000000001000;
		1789: Delta = 30'sb111111111100000000000000001000;
		2758: Delta = 30'sb000000000011111111111111111000;
		1773: Delta = 30'sb111111111011111111111111111000;
		993: Delta = 30'sb000000001000000000000000001000;
		3570: Delta = 30'sb111111111000000000000000001000;
		977: Delta = 30'sb000000000111111111111111111000;
		3554: Delta = 30'sb111111110111111111111111111000;
		1978: Delta = 30'sb000000010000000000000000001000;
		2585: Delta = 30'sb111111110000000000000000001000;
		1962: Delta = 30'sb000000001111111111111111111000;
		2569: Delta = 30'sb111111101111111111111111111000;
		3948: Delta = 30'sb000000100000000000000000001000;
		615: Delta = 30'sb111111100000000000000000001000;
		3932: Delta = 30'sb000000011111111111111111111000;
		599: Delta = 30'sb111111011111111111111111111000;
		3341: Delta = 30'sb000001000000000000000000001000;
		1222: Delta = 30'sb111111000000000000000000001000;
		3325: Delta = 30'sb000000111111111111111111111000;
		1206: Delta = 30'sb111110111111111111111111111000;
		2127: Delta = 30'sb000010000000000000000000001000;
		2436: Delta = 30'sb111110000000000000000000001000;
		2111: Delta = 30'sb000001111111111111111111111000;
		2420: Delta = 30'sb111101111111111111111111111000;
		4246: Delta = 30'sb000100000000000000000000001000;
		317: Delta = 30'sb111100000000000000000000001000;
		4230: Delta = 30'sb000011111111111111111111111000;
		301: Delta = 30'sb111011111111111111111111111000;
		3937: Delta = 30'sb001000000000000000000000001000;
		626: Delta = 30'sb111000000000000000000000001000;
		3921: Delta = 30'sb000111111111111111111111111000;
		610: Delta = 30'sb110111111111111111111111111000;
		3319: Delta = 30'sb010000000000000000000000001000;
		1244: Delta = 30'sb110000000000000000000000001000;
		3303: Delta = 30'sb001111111111111111111111111000;
		1228: Delta = 30'sb101111111111111111111111111000;
		48: Delta = 30'sb000000000000000000000000110000;
		4499: Delta = 30'sb111111111111111111111111010000;
		80: Delta = 30'sb000000000000000000000001010000;
		4467: Delta = 30'sb111111111111111111111110110000;
		144: Delta = 30'sb000000000000000000000010010000;
		4435: Delta = 30'sb111111111111111111111110010000;
		112: Delta = 30'sb000000000000000000000001110000;
		4403: Delta = 30'sb111111111111111111111101110000;
		272: Delta = 30'sb000000000000000000000100010000;
		4307: Delta = 30'sb111111111111111111111100010000;
		240: Delta = 30'sb000000000000000000000011110000;
		4275: Delta = 30'sb111111111111111111111011110000;
		528: Delta = 30'sb000000000000000000001000010000;
		4051: Delta = 30'sb111111111111111111111000010000;
		496: Delta = 30'sb000000000000000000000111110000;
		4019: Delta = 30'sb111111111111111111110111110000;
		1040: Delta = 30'sb000000000000000000010000010000;
		3539: Delta = 30'sb111111111111111111110000010000;
		1008: Delta = 30'sb000000000000000000001111110000;
		3507: Delta = 30'sb111111111111111111101111110000;
		2064: Delta = 30'sb000000000000000000100000010000;
		2515: Delta = 30'sb111111111111111111100000010000;
		2032: Delta = 30'sb000000000000000000011111110000;
		2483: Delta = 30'sb111111111111111111011111110000;
		4112: Delta = 30'sb000000000000000001000000010000;
		467: Delta = 30'sb111111111111111111000000010000;
		4080: Delta = 30'sb000000000000000000111111110000;
		435: Delta = 30'sb111111111111111110111111110000;
		3661: Delta = 30'sb000000000000000010000000010000;
		918: Delta = 30'sb111111111111111110000000010000;
		3629: Delta = 30'sb000000000000000001111111110000;
		886: Delta = 30'sb111111111111111101111111110000;
		2759: Delta = 30'sb000000000000000100000000010000;
		1820: Delta = 30'sb111111111111111100000000010000;
		2727: Delta = 30'sb000000000000000011111111110000;
		1788: Delta = 30'sb111111111111111011111111110000;
		955: Delta = 30'sb000000000000001000000000010000;
		3624: Delta = 30'sb111111111111111000000000010000;
		923: Delta = 30'sb000000000000000111111111110000;
		3592: Delta = 30'sb111111111111110111111111110000;
		1894: Delta = 30'sb000000000000010000000000010000;
		2685: Delta = 30'sb111111111111110000000000010000;
		1862: Delta = 30'sb000000000000001111111111110000;
		2653: Delta = 30'sb111111111111101111111111110000;
		3772: Delta = 30'sb000000000000100000000000010000;
		807: Delta = 30'sb111111111111100000000000010000;
		3740: Delta = 30'sb000000000000011111111111110000;
		775: Delta = 30'sb111111111111011111111111110000;
		2981: Delta = 30'sb000000000001000000000000010000;
		1598: Delta = 30'sb111111111111000000000000010000;
		2949: Delta = 30'sb000000000000111111111111110000;
		1566: Delta = 30'sb111111111110111111111111110000;
		1399: Delta = 30'sb000000000010000000000000010000;
		3180: Delta = 30'sb111111111110000000000000010000;
		1367: Delta = 30'sb000000000001111111111111110000;
		3148: Delta = 30'sb111111111101111111111111110000;
		2782: Delta = 30'sb000000000100000000000000010000;
		1797: Delta = 30'sb111111111100000000000000010000;
		2750: Delta = 30'sb000000000011111111111111110000;
		1765: Delta = 30'sb111111111011111111111111110000;
		1001: Delta = 30'sb000000001000000000000000010000;
		3578: Delta = 30'sb111111111000000000000000010000;
		969: Delta = 30'sb000000000111111111111111110000;
		3546: Delta = 30'sb111111110111111111111111110000;
		1986: Delta = 30'sb000000010000000000000000010000;
		2593: Delta = 30'sb111111110000000000000000010000;
		1954: Delta = 30'sb000000001111111111111111110000;
		2561: Delta = 30'sb111111101111111111111111110000;
		3956: Delta = 30'sb000000100000000000000000010000;
		623: Delta = 30'sb111111100000000000000000010000;
		3924: Delta = 30'sb000000011111111111111111110000;
		591: Delta = 30'sb111111011111111111111111110000;
		3349: Delta = 30'sb000001000000000000000000010000;
		1230: Delta = 30'sb111111000000000000000000010000;
		3317: Delta = 30'sb000000111111111111111111110000;
		1198: Delta = 30'sb111110111111111111111111110000;
		2135: Delta = 30'sb000010000000000000000000010000;
		2444: Delta = 30'sb111110000000000000000000010000;
		2103: Delta = 30'sb000001111111111111111111110000;
		2412: Delta = 30'sb111101111111111111111111110000;
		4254: Delta = 30'sb000100000000000000000000010000;
		325: Delta = 30'sb111100000000000000000000010000;
		4222: Delta = 30'sb000011111111111111111111110000;
		293: Delta = 30'sb111011111111111111111111110000;
		3945: Delta = 30'sb001000000000000000000000010000;
		634: Delta = 30'sb111000000000000000000000010000;
		3913: Delta = 30'sb000111111111111111111111110000;
		602: Delta = 30'sb110111111111111111111111110000;
		3327: Delta = 30'sb010000000000000000000000010000;
		1252: Delta = 30'sb110000000000000000000000010000;
		3295: Delta = 30'sb001111111111111111111111110000;
		1220: Delta = 30'sb101111111111111111111111110000;
		96: Delta = 30'sb000000000000000000000001100000;
		4451: Delta = 30'sb111111111111111111111110100000;
		160: Delta = 30'sb000000000000000000000010100000;
		4387: Delta = 30'sb111111111111111111111101100000;
		288: Delta = 30'sb000000000000000000000100100000;
		4323: Delta = 30'sb111111111111111111111100100000;
		224: Delta = 30'sb000000000000000000000011100000;
		4259: Delta = 30'sb111111111111111111111011100000;
		544: Delta = 30'sb000000000000000000001000100000;
		4067: Delta = 30'sb111111111111111111111000100000;
		480: Delta = 30'sb000000000000000000000111100000;
		4003: Delta = 30'sb111111111111111111110111100000;
		1056: Delta = 30'sb000000000000000000010000100000;
		3555: Delta = 30'sb111111111111111111110000100000;
		992: Delta = 30'sb000000000000000000001111100000;
		3491: Delta = 30'sb111111111111111111101111100000;
		2080: Delta = 30'sb000000000000000000100000100000;
		2531: Delta = 30'sb111111111111111111100000100000;
		2016: Delta = 30'sb000000000000000000011111100000;
		2467: Delta = 30'sb111111111111111111011111100000;
		4128: Delta = 30'sb000000000000000001000000100000;
		483: Delta = 30'sb111111111111111111000000100000;
		4064: Delta = 30'sb000000000000000000111111100000;
		419: Delta = 30'sb111111111111111110111111100000;
		3677: Delta = 30'sb000000000000000010000000100000;
		934: Delta = 30'sb111111111111111110000000100000;
		3613: Delta = 30'sb000000000000000001111111100000;
		870: Delta = 30'sb111111111111111101111111100000;
		2775: Delta = 30'sb000000000000000100000000100000;
		1836: Delta = 30'sb111111111111111100000000100000;
		2711: Delta = 30'sb000000000000000011111111100000;
		1772: Delta = 30'sb111111111111111011111111100000;
		971: Delta = 30'sb000000000000001000000000100000;
		3640: Delta = 30'sb111111111111111000000000100000;
		907: Delta = 30'sb000000000000000111111111100000;
		3576: Delta = 30'sb111111111111110111111111100000;
		1910: Delta = 30'sb000000000000010000000000100000;
		2701: Delta = 30'sb111111111111110000000000100000;
		1846: Delta = 30'sb000000000000001111111111100000;
		2637: Delta = 30'sb111111111111101111111111100000;
		3788: Delta = 30'sb000000000000100000000000100000;
		823: Delta = 30'sb111111111111100000000000100000;
		3724: Delta = 30'sb000000000000011111111111100000;
		759: Delta = 30'sb111111111111011111111111100000;
		2997: Delta = 30'sb000000000001000000000000100000;
		1614: Delta = 30'sb111111111111000000000000100000;
		2933: Delta = 30'sb000000000000111111111111100000;
		1550: Delta = 30'sb111111111110111111111111100000;
		1415: Delta = 30'sb000000000010000000000000100000;
		3196: Delta = 30'sb111111111110000000000000100000;
		1351: Delta = 30'sb000000000001111111111111100000;
		3132: Delta = 30'sb111111111101111111111111100000;
		2798: Delta = 30'sb000000000100000000000000100000;
		1813: Delta = 30'sb111111111100000000000000100000;
		2734: Delta = 30'sb000000000011111111111111100000;
		1749: Delta = 30'sb111111111011111111111111100000;
		1017: Delta = 30'sb000000001000000000000000100000;
		3594: Delta = 30'sb111111111000000000000000100000;
		953: Delta = 30'sb000000000111111111111111100000;
		3530: Delta = 30'sb111111110111111111111111100000;
		2002: Delta = 30'sb000000010000000000000000100000;
		2609: Delta = 30'sb111111110000000000000000100000;
		1938: Delta = 30'sb000000001111111111111111100000;
		2545: Delta = 30'sb111111101111111111111111100000;
		3972: Delta = 30'sb000000100000000000000000100000;
		639: Delta = 30'sb111111100000000000000000100000;
		3908: Delta = 30'sb000000011111111111111111100000;
		575: Delta = 30'sb111111011111111111111111100000;
		3365: Delta = 30'sb000001000000000000000000100000;
		1246: Delta = 30'sb111111000000000000000000100000;
		3301: Delta = 30'sb000000111111111111111111100000;
		1182: Delta = 30'sb111110111111111111111111100000;
		2151: Delta = 30'sb000010000000000000000000100000;
		2460: Delta = 30'sb111110000000000000000000100000;
		2087: Delta = 30'sb000001111111111111111111100000;
		2396: Delta = 30'sb111101111111111111111111100000;
		4270: Delta = 30'sb000100000000000000000000100000;
		341: Delta = 30'sb111100000000000000000000100000;
		4206: Delta = 30'sb000011111111111111111111100000;
		277: Delta = 30'sb111011111111111111111111100000;
		3961: Delta = 30'sb001000000000000000000000100000;
		650: Delta = 30'sb111000000000000000000000100000;
		3897: Delta = 30'sb000111111111111111111111100000;
		586: Delta = 30'sb110111111111111111111111100000;
		3343: Delta = 30'sb010000000000000000000000100000;
		1268: Delta = 30'sb110000000000000000000000100000;
		3279: Delta = 30'sb001111111111111111111111100000;
		1204: Delta = 30'sb101111111111111111111111100000;
		192: Delta = 30'sb000000000000000000000011000000;
		4355: Delta = 30'sb111111111111111111111101000000;
		320: Delta = 30'sb000000000000000000000101000000;
		4227: Delta = 30'sb111111111111111111111011000000;
		576: Delta = 30'sb000000000000000000001001000000;
		4099: Delta = 30'sb111111111111111111111001000000;
		448: Delta = 30'sb000000000000000000000111000000;
		3971: Delta = 30'sb111111111111111111110111000000;
		1088: Delta = 30'sb000000000000000000010001000000;
		3587: Delta = 30'sb111111111111111111110001000000;
		960: Delta = 30'sb000000000000000000001111000000;
		3459: Delta = 30'sb111111111111111111101111000000;
		2112: Delta = 30'sb000000000000000000100001000000;
		2563: Delta = 30'sb111111111111111111100001000000;
		1984: Delta = 30'sb000000000000000000011111000000;
		2435: Delta = 30'sb111111111111111111011111000000;
		4160: Delta = 30'sb000000000000000001000001000000;
		515: Delta = 30'sb111111111111111111000001000000;
		4032: Delta = 30'sb000000000000000000111111000000;
		387: Delta = 30'sb111111111111111110111111000000;
		3709: Delta = 30'sb000000000000000010000001000000;
		966: Delta = 30'sb111111111111111110000001000000;
		3581: Delta = 30'sb000000000000000001111111000000;
		838: Delta = 30'sb111111111111111101111111000000;
		2807: Delta = 30'sb000000000000000100000001000000;
		1868: Delta = 30'sb111111111111111100000001000000;
		2679: Delta = 30'sb000000000000000011111111000000;
		1740: Delta = 30'sb111111111111111011111111000000;
		1003: Delta = 30'sb000000000000001000000001000000;
		3672: Delta = 30'sb111111111111111000000001000000;
		875: Delta = 30'sb000000000000000111111111000000;
		3544: Delta = 30'sb111111111111110111111111000000;
		1942: Delta = 30'sb000000000000010000000001000000;
		2733: Delta = 30'sb111111111111110000000001000000;
		1814: Delta = 30'sb000000000000001111111111000000;
		2605: Delta = 30'sb111111111111101111111111000000;
		3820: Delta = 30'sb000000000000100000000001000000;
		855: Delta = 30'sb111111111111100000000001000000;
		3692: Delta = 30'sb000000000000011111111111000000;
		727: Delta = 30'sb111111111111011111111111000000;
		3029: Delta = 30'sb000000000001000000000001000000;
		1646: Delta = 30'sb111111111111000000000001000000;
		2901: Delta = 30'sb000000000000111111111111000000;
		1518: Delta = 30'sb111111111110111111111111000000;
		1447: Delta = 30'sb000000000010000000000001000000;
		3228: Delta = 30'sb111111111110000000000001000000;
		1319: Delta = 30'sb000000000001111111111111000000;
		3100: Delta = 30'sb111111111101111111111111000000;
		2830: Delta = 30'sb000000000100000000000001000000;
		1845: Delta = 30'sb111111111100000000000001000000;
		2702: Delta = 30'sb000000000011111111111111000000;
		1717: Delta = 30'sb111111111011111111111111000000;
		1049: Delta = 30'sb000000001000000000000001000000;
		3626: Delta = 30'sb111111111000000000000001000000;
		921: Delta = 30'sb000000000111111111111111000000;
		3498: Delta = 30'sb111111110111111111111111000000;
		2034: Delta = 30'sb000000010000000000000001000000;
		2641: Delta = 30'sb111111110000000000000001000000;
		1906: Delta = 30'sb000000001111111111111111000000;
		2513: Delta = 30'sb111111101111111111111111000000;
		4004: Delta = 30'sb000000100000000000000001000000;
		671: Delta = 30'sb111111100000000000000001000000;
		3876: Delta = 30'sb000000011111111111111111000000;
		543: Delta = 30'sb111111011111111111111111000000;
		3397: Delta = 30'sb000001000000000000000001000000;
		1278: Delta = 30'sb111111000000000000000001000000;
		3269: Delta = 30'sb000000111111111111111111000000;
		1150: Delta = 30'sb111110111111111111111111000000;
		2183: Delta = 30'sb000010000000000000000001000000;
		2492: Delta = 30'sb111110000000000000000001000000;
		2055: Delta = 30'sb000001111111111111111111000000;
		2364: Delta = 30'sb111101111111111111111111000000;
		4302: Delta = 30'sb000100000000000000000001000000;
		373: Delta = 30'sb111100000000000000000001000000;
		4174: Delta = 30'sb000011111111111111111111000000;
		245: Delta = 30'sb111011111111111111111111000000;
		3993: Delta = 30'sb001000000000000000000001000000;
		682: Delta = 30'sb111000000000000000000001000000;
		3865: Delta = 30'sb000111111111111111111111000000;
		554: Delta = 30'sb110111111111111111111111000000;
		3375: Delta = 30'sb010000000000000000000001000000;
		1300: Delta = 30'sb110000000000000000000001000000;
		3247: Delta = 30'sb001111111111111111111111000000;
		1172: Delta = 30'sb101111111111111111111111000000;
		384: Delta = 30'sb000000000000000000000110000000;
		4163: Delta = 30'sb111111111111111111111010000000;
		640: Delta = 30'sb000000000000000000001010000000;
		3907: Delta = 30'sb111111111111111111110110000000;
		1152: Delta = 30'sb000000000000000000010010000000;
		3651: Delta = 30'sb111111111111111111110010000000;
		896: Delta = 30'sb000000000000000000001110000000;
		3395: Delta = 30'sb111111111111111111101110000000;
		2176: Delta = 30'sb000000000000000000100010000000;
		2627: Delta = 30'sb111111111111111111100010000000;
		1920: Delta = 30'sb000000000000000000011110000000;
		2371: Delta = 30'sb111111111111111111011110000000;
		4224: Delta = 30'sb000000000000000001000010000000;
		579: Delta = 30'sb111111111111111111000010000000;
		3968: Delta = 30'sb000000000000000000111110000000;
		323: Delta = 30'sb111111111111111110111110000000;
		3773: Delta = 30'sb000000000000000010000010000000;
		1030: Delta = 30'sb111111111111111110000010000000;
		3517: Delta = 30'sb000000000000000001111110000000;
		774: Delta = 30'sb111111111111111101111110000000;
		2871: Delta = 30'sb000000000000000100000010000000;
		1932: Delta = 30'sb111111111111111100000010000000;
		2615: Delta = 30'sb000000000000000011111110000000;
		1676: Delta = 30'sb111111111111111011111110000000;
		1067: Delta = 30'sb000000000000001000000010000000;
		3736: Delta = 30'sb111111111111111000000010000000;
		811: Delta = 30'sb000000000000000111111110000000;
		3480: Delta = 30'sb111111111111110111111110000000;
		2006: Delta = 30'sb000000000000010000000010000000;
		2797: Delta = 30'sb111111111111110000000010000000;
		1750: Delta = 30'sb000000000000001111111110000000;
		2541: Delta = 30'sb111111111111101111111110000000;
		3884: Delta = 30'sb000000000000100000000010000000;
		919: Delta = 30'sb111111111111100000000010000000;
		3628: Delta = 30'sb000000000000011111111110000000;
		663: Delta = 30'sb111111111111011111111110000000;
		3093: Delta = 30'sb000000000001000000000010000000;
		1710: Delta = 30'sb111111111111000000000010000000;
		2837: Delta = 30'sb000000000000111111111110000000;
		1454: Delta = 30'sb111111111110111111111110000000;
		1511: Delta = 30'sb000000000010000000000010000000;
		3292: Delta = 30'sb111111111110000000000010000000;
		1255: Delta = 30'sb000000000001111111111110000000;
		3036: Delta = 30'sb111111111101111111111110000000;
		2894: Delta = 30'sb000000000100000000000010000000;
		1909: Delta = 30'sb111111111100000000000010000000;
		2638: Delta = 30'sb000000000011111111111110000000;
		1653: Delta = 30'sb111111111011111111111110000000;
		1113: Delta = 30'sb000000001000000000000010000000;
		3690: Delta = 30'sb111111111000000000000010000000;
		857: Delta = 30'sb000000000111111111111110000000;
		3434: Delta = 30'sb111111110111111111111110000000;
		2098: Delta = 30'sb000000010000000000000010000000;
		2705: Delta = 30'sb111111110000000000000010000000;
		1842: Delta = 30'sb000000001111111111111110000000;
		2449: Delta = 30'sb111111101111111111111110000000;
		4068: Delta = 30'sb000000100000000000000010000000;
		735: Delta = 30'sb111111100000000000000010000000;
		3812: Delta = 30'sb000000011111111111111110000000;
		479: Delta = 30'sb111111011111111111111110000000;
		3461: Delta = 30'sb000001000000000000000010000000;
		1342: Delta = 30'sb111111000000000000000010000000;
		3205: Delta = 30'sb000000111111111111111110000000;
		1086: Delta = 30'sb111110111111111111111110000000;
		2247: Delta = 30'sb000010000000000000000010000000;
		2556: Delta = 30'sb111110000000000000000010000000;
		1991: Delta = 30'sb000001111111111111111110000000;
		2300: Delta = 30'sb111101111111111111111110000000;
		4366: Delta = 30'sb000100000000000000000010000000;
		437: Delta = 30'sb111100000000000000000010000000;
		4110: Delta = 30'sb000011111111111111111110000000;
		181: Delta = 30'sb111011111111111111111110000000;
		4057: Delta = 30'sb001000000000000000000010000000;
		746: Delta = 30'sb111000000000000000000010000000;
		3801: Delta = 30'sb000111111111111111111110000000;
		490: Delta = 30'sb110111111111111111111110000000;
		3439: Delta = 30'sb010000000000000000000010000000;
		1364: Delta = 30'sb110000000000000000000010000000;
		3183: Delta = 30'sb001111111111111111111110000000;
		1108: Delta = 30'sb101111111111111111111110000000;
		768: Delta = 30'sb000000000000000000001100000000;
		3779: Delta = 30'sb111111111111111111110100000000;
		1280: Delta = 30'sb000000000000000000010100000000;
		3267: Delta = 30'sb111111111111111111101100000000;
		2304: Delta = 30'sb000000000000000000100100000000;
		2755: Delta = 30'sb111111111111111111100100000000;
		1792: Delta = 30'sb000000000000000000011100000000;
		2243: Delta = 30'sb111111111111111111011100000000;
		4352: Delta = 30'sb000000000000000001000100000000;
		707: Delta = 30'sb111111111111111111000100000000;
		3840: Delta = 30'sb000000000000000000111100000000;
		195: Delta = 30'sb111111111111111110111100000000;
		3901: Delta = 30'sb000000000000000010000100000000;
		1158: Delta = 30'sb111111111111111110000100000000;
		3389: Delta = 30'sb000000000000000001111100000000;
		646: Delta = 30'sb111111111111111101111100000000;
		2999: Delta = 30'sb000000000000000100000100000000;
		2060: Delta = 30'sb111111111111111100000100000000;
		2487: Delta = 30'sb000000000000000011111100000000;
		1548: Delta = 30'sb111111111111111011111100000000;
		1195: Delta = 30'sb000000000000001000000100000000;
		3864: Delta = 30'sb111111111111111000000100000000;
		683: Delta = 30'sb000000000000000111111100000000;
		3352: Delta = 30'sb111111111111110111111100000000;
		2134: Delta = 30'sb000000000000010000000100000000;
		2925: Delta = 30'sb111111111111110000000100000000;
		1622: Delta = 30'sb000000000000001111111100000000;
		2413: Delta = 30'sb111111111111101111111100000000;
		4012: Delta = 30'sb000000000000100000000100000000;
		1047: Delta = 30'sb111111111111100000000100000000;
		3500: Delta = 30'sb000000000000011111111100000000;
		535: Delta = 30'sb111111111111011111111100000000;
		3221: Delta = 30'sb000000000001000000000100000000;
		1838: Delta = 30'sb111111111111000000000100000000;
		2709: Delta = 30'sb000000000000111111111100000000;
		1326: Delta = 30'sb111111111110111111111100000000;
		1639: Delta = 30'sb000000000010000000000100000000;
		3420: Delta = 30'sb111111111110000000000100000000;
		1127: Delta = 30'sb000000000001111111111100000000;
		2908: Delta = 30'sb111111111101111111111100000000;
		3022: Delta = 30'sb000000000100000000000100000000;
		2037: Delta = 30'sb111111111100000000000100000000;
		2510: Delta = 30'sb000000000011111111111100000000;
		1525: Delta = 30'sb111111111011111111111100000000;
		1241: Delta = 30'sb000000001000000000000100000000;
		3818: Delta = 30'sb111111111000000000000100000000;
		729: Delta = 30'sb000000000111111111111100000000;
		3306: Delta = 30'sb111111110111111111111100000000;
		2226: Delta = 30'sb000000010000000000000100000000;
		2833: Delta = 30'sb111111110000000000000100000000;
		1714: Delta = 30'sb000000001111111111111100000000;
		2321: Delta = 30'sb111111101111111111111100000000;
		4196: Delta = 30'sb000000100000000000000100000000;
		863: Delta = 30'sb111111100000000000000100000000;
		3684: Delta = 30'sb000000011111111111111100000000;
		351: Delta = 30'sb111111011111111111111100000000;
		3589: Delta = 30'sb000001000000000000000100000000;
		1470: Delta = 30'sb111111000000000000000100000000;
		3077: Delta = 30'sb000000111111111111111100000000;
		958: Delta = 30'sb111110111111111111111100000000;
		2375: Delta = 30'sb000010000000000000000100000000;
		2684: Delta = 30'sb111110000000000000000100000000;
		1863: Delta = 30'sb000001111111111111111100000000;
		2172: Delta = 30'sb111101111111111111111100000000;
		4494: Delta = 30'sb000100000000000000000100000000;
		565: Delta = 30'sb111100000000000000000100000000;
		3982: Delta = 30'sb000011111111111111111100000000;
		53: Delta = 30'sb111011111111111111111100000000;
		4185: Delta = 30'sb001000000000000000000100000000;
		874: Delta = 30'sb111000000000000000000100000000;
		3673: Delta = 30'sb000111111111111111111100000000;
		362: Delta = 30'sb110111111111111111111100000000;
		3567: Delta = 30'sb010000000000000000000100000000;
		1492: Delta = 30'sb110000000000000000000100000000;
		3055: Delta = 30'sb001111111111111111111100000000;
		980: Delta = 30'sb101111111111111111111100000000;
		1536: Delta = 30'sb000000000000000000011000000000;
		3011: Delta = 30'sb111111111111111111101000000000;
		2560: Delta = 30'sb000000000000000000101000000000;
		1987: Delta = 30'sb111111111111111111011000000000;
		61: Delta = 30'sb000000000000000001001000000000;
		963: Delta = 30'sb111111111111111111001000000000;
		3584: Delta = 30'sb000000000000000000111000000000;
		4486: Delta = 30'sb111111111111111110111000000000;
		4157: Delta = 30'sb000000000000000010001000000000;
		1414: Delta = 30'sb111111111111111110001000000000;
		3133: Delta = 30'sb000000000000000001111000000000;
		390: Delta = 30'sb111111111111111101111000000000;
		3255: Delta = 30'sb000000000000000100001000000000;
		2316: Delta = 30'sb111111111111111100001000000000;
		2231: Delta = 30'sb000000000000000011111000000000;
		1292: Delta = 30'sb111111111111111011111000000000;
		1451: Delta = 30'sb000000000000001000001000000000;
		4120: Delta = 30'sb111111111111111000001000000000;
		427: Delta = 30'sb000000000000000111111000000000;
		3096: Delta = 30'sb111111111111110111111000000000;
		2390: Delta = 30'sb000000000000010000001000000000;
		3181: Delta = 30'sb111111111111110000001000000000;
		1366: Delta = 30'sb000000000000001111111000000000;
		2157: Delta = 30'sb111111111111101111111000000000;
		4268: Delta = 30'sb000000000000100000001000000000;
		1303: Delta = 30'sb111111111111100000001000000000;
		3244: Delta = 30'sb000000000000011111111000000000;
		279: Delta = 30'sb111111111111011111111000000000;
		3477: Delta = 30'sb000000000001000000001000000000;
		2094: Delta = 30'sb111111111111000000001000000000;
		2453: Delta = 30'sb000000000000111111111000000000;
		1070: Delta = 30'sb111111111110111111111000000000;
		1895: Delta = 30'sb000000000010000000001000000000;
		3676: Delta = 30'sb111111111110000000001000000000;
		871: Delta = 30'sb000000000001111111111000000000;
		2652: Delta = 30'sb111111111101111111111000000000;
		3278: Delta = 30'sb000000000100000000001000000000;
		2293: Delta = 30'sb111111111100000000001000000000;
		2254: Delta = 30'sb000000000011111111111000000000;
		1269: Delta = 30'sb111111111011111111111000000000;
		1497: Delta = 30'sb000000001000000000001000000000;
		4074: Delta = 30'sb111111111000000000001000000000;
		473: Delta = 30'sb000000000111111111111000000000;
		3050: Delta = 30'sb111111110111111111111000000000;
		2482: Delta = 30'sb000000010000000000001000000000;
		3089: Delta = 30'sb111111110000000000001000000000;
		1458: Delta = 30'sb000000001111111111111000000000;
		2065: Delta = 30'sb111111101111111111111000000000;
		4452: Delta = 30'sb000000100000000000001000000000;
		1119: Delta = 30'sb111111100000000000001000000000;
		3428: Delta = 30'sb000000011111111111111000000000;
		95: Delta = 30'sb111111011111111111111000000000;
		3845: Delta = 30'sb000001000000000000001000000000;
		1726: Delta = 30'sb111111000000000000001000000000;
		2821: Delta = 30'sb000000111111111111111000000000;
		702: Delta = 30'sb111110111111111111111000000000;
		2631: Delta = 30'sb000010000000000000001000000000;
		2940: Delta = 30'sb111110000000000000001000000000;
		1607: Delta = 30'sb000001111111111111111000000000;
		1916: Delta = 30'sb111101111111111111111000000000;
		203: Delta = 30'sb000100000000000000001000000000;
		821: Delta = 30'sb111100000000000000001000000000;
		3726: Delta = 30'sb000011111111111111111000000000;
		4344: Delta = 30'sb111011111111111111111000000000;
		4441: Delta = 30'sb001000000000000000001000000000;
		1130: Delta = 30'sb111000000000000000001000000000;
		3417: Delta = 30'sb000111111111111111111000000000;
		106: Delta = 30'sb110111111111111111111000000000;
		3823: Delta = 30'sb010000000000000000001000000000;
		1748: Delta = 30'sb110000000000000000001000000000;
		2799: Delta = 30'sb001111111111111111111000000000;
		724: Delta = 30'sb101111111111111111111000000000;
		3072: Delta = 30'sb000000000000000000110000000000;
		1475: Delta = 30'sb111111111111111111010000000000;
		573: Delta = 30'sb000000000000000001010000000000;
		3974: Delta = 30'sb111111111111111110110000000000;
		122: Delta = 30'sb000000000000000010010000000000;
		1926: Delta = 30'sb111111111111111110010000000000;
		2621: Delta = 30'sb000000000000000001110000000000;
		4425: Delta = 30'sb111111111111111101110000000000;
		3767: Delta = 30'sb000000000000000100010000000000;
		2828: Delta = 30'sb111111111111111100010000000000;
		1719: Delta = 30'sb000000000000000011110000000000;
		780: Delta = 30'sb111111111111111011110000000000;
		1963: Delta = 30'sb000000000000001000010000000000;
		85: Delta = 30'sb111111111111111000010000000000;
		4462: Delta = 30'sb000000000000000111110000000000;
		2584: Delta = 30'sb111111111111110111110000000000;
		2902: Delta = 30'sb000000000000010000010000000000;
		3693: Delta = 30'sb111111111111110000010000000000;
		854: Delta = 30'sb000000000000001111110000000000;
		1645: Delta = 30'sb111111111111101111110000000000;
		233: Delta = 30'sb000000000000100000010000000000;
		1815: Delta = 30'sb111111111111100000010000000000;
		2732: Delta = 30'sb000000000000011111110000000000;
		4314: Delta = 30'sb111111111111011111110000000000;
		3989: Delta = 30'sb000000000001000000010000000000;
		2606: Delta = 30'sb111111111111000000010000000000;
		1941: Delta = 30'sb000000000000111111110000000000;
		558: Delta = 30'sb111111111110111111110000000000;
		2407: Delta = 30'sb000000000010000000010000000000;
		4188: Delta = 30'sb111111111110000000010000000000;
		359: Delta = 30'sb000000000001111111110000000000;
		2140: Delta = 30'sb111111111101111111110000000000;
		3790: Delta = 30'sb000000000100000000010000000000;
		2805: Delta = 30'sb111111111100000000010000000000;
		1742: Delta = 30'sb000000000011111111110000000000;
		757: Delta = 30'sb111111111011111111110000000000;
		2009: Delta = 30'sb000000001000000000010000000000;
		39: Delta = 30'sb111111111000000000010000000000;
		4508: Delta = 30'sb000000000111111111110000000000;
		2538: Delta = 30'sb111111110111111111110000000000;
		2994: Delta = 30'sb000000010000000000010000000000;
		3601: Delta = 30'sb111111110000000000010000000000;
		946: Delta = 30'sb000000001111111111110000000000;
		1553: Delta = 30'sb111111101111111111110000000000;
		417: Delta = 30'sb000000100000000000010000000000;
		1631: Delta = 30'sb111111100000000000010000000000;
		2916: Delta = 30'sb000000011111111111110000000000;
		4130: Delta = 30'sb111111011111111111110000000000;
		4357: Delta = 30'sb000001000000000000010000000000;
		2238: Delta = 30'sb111111000000000000010000000000;
		2309: Delta = 30'sb000000111111111111110000000000;
		190: Delta = 30'sb111110111111111111110000000000;
		3143: Delta = 30'sb000010000000000000010000000000;
		3452: Delta = 30'sb111110000000000000010000000000;
		1095: Delta = 30'sb000001111111111111110000000000;
		1404: Delta = 30'sb111101111111111111110000000000;
		715: Delta = 30'sb000100000000000000010000000000;
		1333: Delta = 30'sb111100000000000000010000000000;
		3214: Delta = 30'sb000011111111111111110000000000;
		3832: Delta = 30'sb111011111111111111110000000000;
		406: Delta = 30'sb001000000000000000010000000000;
		1642: Delta = 30'sb111000000000000000010000000000;
		2905: Delta = 30'sb000111111111111111110000000000;
		4141: Delta = 30'sb110111111111111111110000000000;
		4335: Delta = 30'sb010000000000000000010000000000;
		2260: Delta = 30'sb110000000000000000010000000000;
		2287: Delta = 30'sb001111111111111111110000000000;
		212: Delta = 30'sb101111111111111111110000000000;
		1597: Delta = 30'sb000000000000000001100000000000;
		2950: Delta = 30'sb111111111111111110100000000000;
		1146: Delta = 30'sb000000000000000010100000000000;
		3401: Delta = 30'sb111111111111111101100000000000;
		244: Delta = 30'sb000000000000000100100000000000;
		3852: Delta = 30'sb111111111111111100100000000000;
		695: Delta = 30'sb000000000000000011100000000000;
		4303: Delta = 30'sb111111111111111011100000000000;
		2987: Delta = 30'sb000000000000001000100000000000;
		1109: Delta = 30'sb111111111111111000100000000000;
		3438: Delta = 30'sb000000000000000111100000000000;
		1560: Delta = 30'sb111111111111110111100000000000;
		3926: Delta = 30'sb000000000000010000100000000000;
		170: Delta = 30'sb111111111111110000100000000000;
		4377: Delta = 30'sb000000000000001111100000000000;
		621: Delta = 30'sb111111111111101111100000000000;
		1257: Delta = 30'sb000000000000100000100000000000;
		2839: Delta = 30'sb111111111111100000100000000000;
		1708: Delta = 30'sb000000000000011111100000000000;
		3290: Delta = 30'sb111111111111011111100000000000;
		466: Delta = 30'sb000000000001000000100000000000;
		3630: Delta = 30'sb111111111111000000100000000000;
		917: Delta = 30'sb000000000000111111100000000000;
		4081: Delta = 30'sb111111111110111111100000000000;
		3431: Delta = 30'sb000000000010000000100000000000;
		665: Delta = 30'sb111111111110000000100000000000;
		3882: Delta = 30'sb000000000001111111100000000000;
		1116: Delta = 30'sb111111111101111111100000000000;
		267: Delta = 30'sb000000000100000000100000000000;
		3829: Delta = 30'sb111111111100000000100000000000;
		718: Delta = 30'sb000000000011111111100000000000;
		4280: Delta = 30'sb111111111011111111100000000000;
		3033: Delta = 30'sb000000001000000000100000000000;
		1063: Delta = 30'sb111111111000000000100000000000;
		3484: Delta = 30'sb000000000111111111100000000000;
		1514: Delta = 30'sb111111110111111111100000000000;
		4018: Delta = 30'sb000000010000000000100000000000;
		78: Delta = 30'sb111111110000000000100000000000;
		4469: Delta = 30'sb000000001111111111100000000000;
		529: Delta = 30'sb111111101111111111100000000000;
		1441: Delta = 30'sb000000100000000000100000000000;
		2655: Delta = 30'sb111111100000000000100000000000;
		1892: Delta = 30'sb000000011111111111100000000000;
		3106: Delta = 30'sb111111011111111111100000000000;
		834: Delta = 30'sb000001000000000000100000000000;
		3262: Delta = 30'sb111111000000000000100000000000;
		1285: Delta = 30'sb000000111111111111100000000000;
		3713: Delta = 30'sb111110111111111111100000000000;
		4167: Delta = 30'sb000010000000000000100000000000;
		4476: Delta = 30'sb111110000000000000100000000000;
		71: Delta = 30'sb000001111111111111100000000000;
		380: Delta = 30'sb111101111111111111100000000000;
		1739: Delta = 30'sb000100000000000000100000000000;
		2357: Delta = 30'sb111100000000000000100000000000;
		2190: Delta = 30'sb000011111111111111100000000000;
		2808: Delta = 30'sb111011111111111111100000000000;
		1430: Delta = 30'sb001000000000000000100000000000;
		2666: Delta = 30'sb111000000000000000100000000000;
		1881: Delta = 30'sb000111111111111111100000000000;
		3117: Delta = 30'sb110111111111111111100000000000;
		812: Delta = 30'sb010000000000000000100000000000;
		3284: Delta = 30'sb110000000000000000100000000000;
		1263: Delta = 30'sb001111111111111111100000000000;
		3735: Delta = 30'sb101111111111111111100000000000;
		3194: Delta = 30'sb000000000000000011000000000000;
		1353: Delta = 30'sb111111111111111101000000000000;
		2292: Delta = 30'sb000000000000000101000000000000;
		2255: Delta = 30'sb111111111111111011000000000000;
		488: Delta = 30'sb000000000000001001000000000000;
		3157: Delta = 30'sb111111111111111001000000000000;
		1390: Delta = 30'sb000000000000000111000000000000;
		4059: Delta = 30'sb111111111111110111000000000000;
		1427: Delta = 30'sb000000000000010001000000000000;
		2218: Delta = 30'sb111111111111110001000000000000;
		2329: Delta = 30'sb000000000000001111000000000000;
		3120: Delta = 30'sb111111111111101111000000000000;
		3305: Delta = 30'sb000000000000100001000000000000;
		340: Delta = 30'sb111111111111100001000000000000;
		4207: Delta = 30'sb000000000000011111000000000000;
		1242: Delta = 30'sb111111111111011111000000000000;
		2514: Delta = 30'sb000000000001000001000000000000;
		1131: Delta = 30'sb111111111111000001000000000000;
		3416: Delta = 30'sb000000000000111111000000000000;
		2033: Delta = 30'sb111111111110111111000000000000;
		932: Delta = 30'sb000000000010000001000000000000;
		2713: Delta = 30'sb111111111110000001000000000000;
		1834: Delta = 30'sb000000000001111111000000000000;
		3615: Delta = 30'sb111111111101111111000000000000;
		2315: Delta = 30'sb000000000100000001000000000000;
		1330: Delta = 30'sb111111111100000001000000000000;
		3217: Delta = 30'sb000000000011111111000000000000;
		2232: Delta = 30'sb111111111011111111000000000000;
		534: Delta = 30'sb000000001000000001000000000000;
		3111: Delta = 30'sb111111111000000001000000000000;
		1436: Delta = 30'sb000000000111111111000000000000;
		4013: Delta = 30'sb111111110111111111000000000000;
		1519: Delta = 30'sb000000010000000001000000000000;
		2126: Delta = 30'sb111111110000000001000000000000;
		2421: Delta = 30'sb000000001111111111000000000000;
		3028: Delta = 30'sb111111101111111111000000000000;
		3489: Delta = 30'sb000000100000000001000000000000;
		156: Delta = 30'sb111111100000000001000000000000;
		4391: Delta = 30'sb000000011111111111000000000000;
		1058: Delta = 30'sb111111011111111111000000000000;
		2882: Delta = 30'sb000001000000000001000000000000;
		763: Delta = 30'sb111111000000000001000000000000;
		3784: Delta = 30'sb000000111111111111000000000000;
		1665: Delta = 30'sb111110111111111111000000000000;
		1668: Delta = 30'sb000010000000000001000000000000;
		1977: Delta = 30'sb111110000000000001000000000000;
		2570: Delta = 30'sb000001111111111111000000000000;
		2879: Delta = 30'sb111101111111111111000000000000;
		3787: Delta = 30'sb000100000000000001000000000000;
		4405: Delta = 30'sb111100000000000001000000000000;
		142: Delta = 30'sb000011111111111111000000000000;
		760: Delta = 30'sb111011111111111111000000000000;
		3478: Delta = 30'sb001000000000000001000000000000;
		167: Delta = 30'sb111000000000000001000000000000;
		4380: Delta = 30'sb000111111111111111000000000000;
		1069: Delta = 30'sb110111111111111111000000000000;
		2860: Delta = 30'sb010000000000000001000000000000;
		785: Delta = 30'sb110000000000000001000000000000;
		3762: Delta = 30'sb001111111111111111000000000000;
		1687: Delta = 30'sb101111111111111111000000000000;
		1841: Delta = 30'sb000000000000000110000000000000;
		2706: Delta = 30'sb111111111111111010000000000000;
		37: Delta = 30'sb000000000000001010000000000000;
		4510: Delta = 30'sb111111111111110110000000000000;
		976: Delta = 30'sb000000000000010010000000000000;
		1767: Delta = 30'sb111111111111110010000000000000;
		2780: Delta = 30'sb000000000000001110000000000000;
		3571: Delta = 30'sb111111111111101110000000000000;
		2854: Delta = 30'sb000000000000100010000000000000;
		4436: Delta = 30'sb111111111111100010000000000000;
		111: Delta = 30'sb000000000000011110000000000000;
		1693: Delta = 30'sb111111111111011110000000000000;
		2063: Delta = 30'sb000000000001000010000000000000;
		680: Delta = 30'sb111111111111000010000000000000;
		3867: Delta = 30'sb000000000000111110000000000000;
		2484: Delta = 30'sb111111111110111110000000000000;
		481: Delta = 30'sb000000000010000010000000000000;
		2262: Delta = 30'sb111111111110000010000000000000;
		2285: Delta = 30'sb000000000001111110000000000000;
		4066: Delta = 30'sb111111111101111110000000000000;
		1864: Delta = 30'sb000000000100000010000000000000;
		879: Delta = 30'sb111111111100000010000000000000;
		3668: Delta = 30'sb000000000011111110000000000000;
		2683: Delta = 30'sb111111111011111110000000000000;
		83: Delta = 30'sb000000001000000010000000000000;
		2660: Delta = 30'sb111111111000000010000000000000;
		1887: Delta = 30'sb000000000111111110000000000000;
		4464: Delta = 30'sb111111110111111110000000000000;
		1068: Delta = 30'sb000000010000000010000000000000;
		1675: Delta = 30'sb111111110000000010000000000000;
		2872: Delta = 30'sb000000001111111110000000000000;
		3479: Delta = 30'sb111111101111111110000000000000;
		3038: Delta = 30'sb000000100000000010000000000000;
		4252: Delta = 30'sb111111100000000010000000000000;
		295: Delta = 30'sb000000011111111110000000000000;
		1509: Delta = 30'sb111111011111111110000000000000;
		2431: Delta = 30'sb000001000000000010000000000000;
		312: Delta = 30'sb111111000000000010000000000000;
		4235: Delta = 30'sb000000111111111110000000000000;
		2116: Delta = 30'sb111110111111111110000000000000;
		1217: Delta = 30'sb000010000000000010000000000000;
		1526: Delta = 30'sb111110000000000010000000000000;
		3021: Delta = 30'sb000001111111111110000000000000;
		3330: Delta = 30'sb111101111111111110000000000000;
		3336: Delta = 30'sb000100000000000010000000000000;
		3954: Delta = 30'sb111100000000000010000000000000;
		593: Delta = 30'sb000011111111111110000000000000;
		1211: Delta = 30'sb111011111111111110000000000000;
		3027: Delta = 30'sb001000000000000010000000000000;
		4263: Delta = 30'sb111000000000000010000000000000;
		284: Delta = 30'sb000111111111111110000000000000;
		1520: Delta = 30'sb110111111111111110000000000000;
		2409: Delta = 30'sb010000000000000010000000000000;
		334: Delta = 30'sb110000000000000010000000000000;
		4213: Delta = 30'sb001111111111111110000000000000;
		2138: Delta = 30'sb101111111111111110000000000000;
		3682: Delta = 30'sb000000000000001100000000000000;
		865: Delta = 30'sb111111111111110100000000000000;
		74: Delta = 30'sb000000000000010100000000000000;
		4473: Delta = 30'sb111111111111101100000000000000;
		1952: Delta = 30'sb000000000000100100000000000000;
		3534: Delta = 30'sb111111111111100100000000000000;
		1013: Delta = 30'sb000000000000011100000000000000;
		2595: Delta = 30'sb111111111111011100000000000000;
		1161: Delta = 30'sb000000000001000100000000000000;
		4325: Delta = 30'sb111111111111000100000000000000;
		222: Delta = 30'sb000000000000111100000000000000;
		3386: Delta = 30'sb111111111110111100000000000000;
		4126: Delta = 30'sb000000000010000100000000000000;
		1360: Delta = 30'sb111111111110000100000000000000;
		3187: Delta = 30'sb000000000001111100000000000000;
		421: Delta = 30'sb111111111101111100000000000000;
		962: Delta = 30'sb000000000100000100000000000000;
		4524: Delta = 30'sb111111111100000100000000000000;
		23: Delta = 30'sb000000000011111100000000000000;
		3585: Delta = 30'sb111111111011111100000000000000;
		3728: Delta = 30'sb000000001000000100000000000000;
		1758: Delta = 30'sb111111111000000100000000000000;
		2789: Delta = 30'sb000000000111111100000000000000;
		819: Delta = 30'sb111111110111111100000000000000;
		166: Delta = 30'sb000000010000000100000000000000;
		773: Delta = 30'sb111111110000000100000000000000;
		3774: Delta = 30'sb000000001111111100000000000000;
		4381: Delta = 30'sb111111101111111100000000000000;
		2136: Delta = 30'sb000000100000000100000000000000;
		3350: Delta = 30'sb111111100000000100000000000000;
		1197: Delta = 30'sb000000011111111100000000000000;
		2411: Delta = 30'sb111111011111111100000000000000;
		1529: Delta = 30'sb000001000000000100000000000000;
		3957: Delta = 30'sb111111000000000100000000000000;
		590: Delta = 30'sb000000111111111100000000000000;
		3018: Delta = 30'sb111110111111111100000000000000;
		315: Delta = 30'sb000010000000000100000000000000;
		624: Delta = 30'sb111110000000000100000000000000;
		3923: Delta = 30'sb000001111111111100000000000000;
		4232: Delta = 30'sb111101111111111100000000000000;
		2434: Delta = 30'sb000100000000000100000000000000;
		3052: Delta = 30'sb111100000000000100000000000000;
		1495: Delta = 30'sb000011111111111100000000000000;
		2113: Delta = 30'sb111011111111111100000000000000;
		2125: Delta = 30'sb001000000000000100000000000000;
		3361: Delta = 30'sb111000000000000100000000000000;
		1186: Delta = 30'sb000111111111111100000000000000;
		2422: Delta = 30'sb110111111111111100000000000000;
		1507: Delta = 30'sb010000000000000100000000000000;
		3979: Delta = 30'sb110000000000000100000000000000;
		568: Delta = 30'sb001111111111111100000000000000;
		3040: Delta = 30'sb101111111111111100000000000000;
		2817: Delta = 30'sb000000000000011000000000000000;
		1730: Delta = 30'sb111111111111101000000000000000;
		148: Delta = 30'sb000000000000101000000000000000;
		4399: Delta = 30'sb111111111111011000000000000000;
		3904: Delta = 30'sb000000000001001000000000000000;
		2521: Delta = 30'sb111111111111001000000000000000;
		2026: Delta = 30'sb000000000000111000000000000000;
		643: Delta = 30'sb111111111110111000000000000000;
		2322: Delta = 30'sb000000000010001000000000000000;
		4103: Delta = 30'sb111111111110001000000000000000;
		444: Delta = 30'sb000000000001111000000000000000;
		2225: Delta = 30'sb111111111101111000000000000000;
		3705: Delta = 30'sb000000000100001000000000000000;
		2720: Delta = 30'sb111111111100001000000000000000;
		1827: Delta = 30'sb000000000011111000000000000000;
		842: Delta = 30'sb111111111011111000000000000000;
		1924: Delta = 30'sb000000001000001000000000000000;
		4501: Delta = 30'sb111111111000001000000000000000;
		46: Delta = 30'sb000000000111111000000000000000;
		2623: Delta = 30'sb111111110111111000000000000000;
		2909: Delta = 30'sb000000010000001000000000000000;
		3516: Delta = 30'sb111111110000001000000000000000;
		1031: Delta = 30'sb000000001111111000000000000000;
		1638: Delta = 30'sb111111101111111000000000000000;
		332: Delta = 30'sb000000100000001000000000000000;
		1546: Delta = 30'sb111111100000001000000000000000;
		3001: Delta = 30'sb000000011111111000000000000000;
		4215: Delta = 30'sb111111011111111000000000000000;
		4272: Delta = 30'sb000001000000001000000000000000;
		2153: Delta = 30'sb111111000000001000000000000000;
		2394: Delta = 30'sb000000111111111000000000000000;
		275: Delta = 30'sb111110111111111000000000000000;
		3058: Delta = 30'sb000010000000001000000000000000;
		3367: Delta = 30'sb111110000000001000000000000000;
		1180: Delta = 30'sb000001111111111000000000000000;
		1489: Delta = 30'sb111101111111111000000000000000;
		630: Delta = 30'sb000100000000001000000000000000;
		1248: Delta = 30'sb111100000000001000000000000000;
		3299: Delta = 30'sb000011111111111000000000000000;
		3917: Delta = 30'sb111011111111111000000000000000;
		321: Delta = 30'sb001000000000001000000000000000;
		1557: Delta = 30'sb111000000000001000000000000000;
		2990: Delta = 30'sb000111111111111000000000000000;
		4226: Delta = 30'sb110111111111111000000000000000;
		4250: Delta = 30'sb010000000000001000000000000000;
		2175: Delta = 30'sb110000000000001000000000000000;
		2372: Delta = 30'sb001111111111111000000000000000;
		297: Delta = 30'sb101111111111111000000000000000;
		1087: Delta = 30'sb000000000000110000000000000000;
		3460: Delta = 30'sb111111111111010000000000000000;
		296: Delta = 30'sb000000000001010000000000000000;
		4251: Delta = 30'sb111111111110110000000000000000;
		3261: Delta = 30'sb000000000010010000000000000000;
		495: Delta = 30'sb111111111110010000000000000000;
		4052: Delta = 30'sb000000000001110000000000000000;
		1286: Delta = 30'sb111111111101110000000000000000;
		97: Delta = 30'sb000000000100010000000000000000;
		3659: Delta = 30'sb111111111100010000000000000000;
		888: Delta = 30'sb000000000011110000000000000000;
		4450: Delta = 30'sb111111111011110000000000000000;
		2863: Delta = 30'sb000000001000010000000000000000;
		893: Delta = 30'sb111111111000010000000000000000;
		3654: Delta = 30'sb000000000111110000000000000000;
		1684: Delta = 30'sb111111110111110000000000000000;
		3848: Delta = 30'sb000000010000010000000000000000;
		4455: Delta = 30'sb111111110000010000000000000000;
		92: Delta = 30'sb000000001111110000000000000000;
		699: Delta = 30'sb111111101111110000000000000000;
		1271: Delta = 30'sb000000100000010000000000000000;
		2485: Delta = 30'sb111111100000010000000000000000;
		2062: Delta = 30'sb000000011111110000000000000000;
		3276: Delta = 30'sb111111011111110000000000000000;
		664: Delta = 30'sb000001000000010000000000000000;
		3092: Delta = 30'sb111111000000010000000000000000;
		1455: Delta = 30'sb000000111111110000000000000000;
		3883: Delta = 30'sb111110111111110000000000000000;
		3997: Delta = 30'sb000010000000010000000000000000;
		4306: Delta = 30'sb111110000000010000000000000000;
		241: Delta = 30'sb000001111111110000000000000000;
		550: Delta = 30'sb111101111111110000000000000000;
		1569: Delta = 30'sb000100000000010000000000000000;
		2187: Delta = 30'sb111100000000010000000000000000;
		2360: Delta = 30'sb000011111111110000000000000000;
		2978: Delta = 30'sb111011111111110000000000000000;
		1260: Delta = 30'sb001000000000010000000000000000;
		2496: Delta = 30'sb111000000000010000000000000000;
		2051: Delta = 30'sb000111111111110000000000000000;
		3287: Delta = 30'sb110111111111110000000000000000;
		642: Delta = 30'sb010000000000010000000000000000;
		3114: Delta = 30'sb110000000000010000000000000000;
		1433: Delta = 30'sb001111111111110000000000000000;
		3905: Delta = 30'sb101111111111110000000000000000;
		2174: Delta = 30'sb000000000001100000000000000000;
		2373: Delta = 30'sb111111111110100000000000000000;
		592: Delta = 30'sb000000000010100000000000000000;
		3955: Delta = 30'sb111111111101100000000000000000;
		1975: Delta = 30'sb000000000100100000000000000000;
		990: Delta = 30'sb111111111100100000000000000000;
		3557: Delta = 30'sb000000000011100000000000000000;
		2572: Delta = 30'sb111111111011100000000000000000;
		194: Delta = 30'sb000000001000100000000000000000;
		2771: Delta = 30'sb111111111000100000000000000000;
		1776: Delta = 30'sb000000000111100000000000000000;
		4353: Delta = 30'sb111111110111100000000000000000;
		1179: Delta = 30'sb000000010000100000000000000000;
		1786: Delta = 30'sb111111110000100000000000000000;
		2761: Delta = 30'sb000000001111100000000000000000;
		3368: Delta = 30'sb111111101111100000000000000000;
		3149: Delta = 30'sb000000100000100000000000000000;
		4363: Delta = 30'sb111111100000100000000000000000;
		184: Delta = 30'sb000000011111100000000000000000;
		1398: Delta = 30'sb111111011111100000000000000000;
		2542: Delta = 30'sb000001000000100000000000000000;
		423: Delta = 30'sb111111000000100000000000000000;
		4124: Delta = 30'sb000000111111100000000000000000;
		2005: Delta = 30'sb111110111111100000000000000000;
		1328: Delta = 30'sb000010000000100000000000000000;
		1637: Delta = 30'sb111110000000100000000000000000;
		2910: Delta = 30'sb000001111111100000000000000000;
		3219: Delta = 30'sb111101111111100000000000000000;
		3447: Delta = 30'sb000100000000100000000000000000;
		4065: Delta = 30'sb111100000000100000000000000000;
		482: Delta = 30'sb000011111111100000000000000000;
		1100: Delta = 30'sb111011111111100000000000000000;
		3138: Delta = 30'sb001000000000100000000000000000;
		4374: Delta = 30'sb111000000000100000000000000000;
		173: Delta = 30'sb000111111111100000000000000000;
		1409: Delta = 30'sb110111111111100000000000000000;
		2520: Delta = 30'sb010000000000100000000000000000;
		445: Delta = 30'sb110000000000100000000000000000;
		4102: Delta = 30'sb001111111111100000000000000000;
		2027: Delta = 30'sb101111111111100000000000000000;
		4348: Delta = 30'sb000000000011000000000000000000;
		199: Delta = 30'sb111111111101000000000000000000;
		1184: Delta = 30'sb000000000101000000000000000000;
		3363: Delta = 30'sb111111111011000000000000000000;
		3950: Delta = 30'sb000000001001000000000000000000;
		1980: Delta = 30'sb111111111001000000000000000000;
		2567: Delta = 30'sb000000000111000000000000000000;
		597: Delta = 30'sb111111110111000000000000000000;
		388: Delta = 30'sb000000010001000000000000000000;
		995: Delta = 30'sb111111110001000000000000000000;
		3552: Delta = 30'sb000000001111000000000000000000;
		4159: Delta = 30'sb111111101111000000000000000000;
		2358: Delta = 30'sb000000100001000000000000000000;
		3572: Delta = 30'sb111111100001000000000000000000;
		975: Delta = 30'sb000000011111000000000000000000;
		2189: Delta = 30'sb111111011111000000000000000000;
		1751: Delta = 30'sb000001000001000000000000000000;
		4179: Delta = 30'sb111111000001000000000000000000;
		368: Delta = 30'sb000000111111000000000000000000;
		2796: Delta = 30'sb111110111111000000000000000000;
		537: Delta = 30'sb000010000001000000000000000000;
		846: Delta = 30'sb111110000001000000000000000000;
		3701: Delta = 30'sb000001111111000000000000000000;
		4010: Delta = 30'sb111101111111000000000000000000;
		2656: Delta = 30'sb000100000001000000000000000000;
		3274: Delta = 30'sb111100000001000000000000000000;
		1273: Delta = 30'sb000011111111000000000000000000;
		1891: Delta = 30'sb111011111111000000000000000000;
		2347: Delta = 30'sb001000000001000000000000000000;
		3583: Delta = 30'sb111000000001000000000000000000;
		964: Delta = 30'sb000111111111000000000000000000;
		2200: Delta = 30'sb110111111111000000000000000000;
		1729: Delta = 30'sb010000000001000000000000000000;
		4201: Delta = 30'sb110000000001000000000000000000;
		346: Delta = 30'sb001111111111000000000000000000;
		2818: Delta = 30'sb101111111111000000000000000000;
		4149: Delta = 30'sb000000000110000000000000000000;
		398: Delta = 30'sb111111111010000000000000000000;
		2368: Delta = 30'sb000000001010000000000000000000;
		2179: Delta = 30'sb111111110110000000000000000000;
		3353: Delta = 30'sb000000010010000000000000000000;
		3960: Delta = 30'sb111111110010000000000000000000;
		587: Delta = 30'sb000000001110000000000000000000;
		1194: Delta = 30'sb111111101110000000000000000000;
		776: Delta = 30'sb000000100010000000000000000000;
		1990: Delta = 30'sb111111100010000000000000000000;
		2557: Delta = 30'sb000000011110000000000000000000;
		3771: Delta = 30'sb111111011110000000000000000000;
		169: Delta = 30'sb000001000010000000000000000000;
		2597: Delta = 30'sb111111000010000000000000000000;
		1950: Delta = 30'sb000000111110000000000000000000;
		4378: Delta = 30'sb111110111110000000000000000000;
		3502: Delta = 30'sb000010000010000000000000000000;
		3811: Delta = 30'sb111110000010000000000000000000;
		736: Delta = 30'sb000001111110000000000000000000;
		1045: Delta = 30'sb111101111110000000000000000000;
		1074: Delta = 30'sb000100000010000000000000000000;
		1692: Delta = 30'sb111100000010000000000000000000;
		2855: Delta = 30'sb000011111110000000000000000000;
		3473: Delta = 30'sb111011111110000000000000000000;
		765: Delta = 30'sb001000000010000000000000000000;
		2001: Delta = 30'sb111000000010000000000000000000;
		2546: Delta = 30'sb000111111110000000000000000000;
		3782: Delta = 30'sb110111111110000000000000000000;
		147: Delta = 30'sb010000000010000000000000000000;
		2619: Delta = 30'sb110000000010000000000000000000;
		1928: Delta = 30'sb001111111110000000000000000000;
		4400: Delta = 30'sb101111111110000000000000000000;
		3751: Delta = 30'sb000000001100000000000000000000;
		796: Delta = 30'sb111111110100000000000000000000;
		189: Delta = 30'sb000000010100000000000000000000;
		4358: Delta = 30'sb111111101100000000000000000000;
		2159: Delta = 30'sb000000100100000000000000000000;
		3373: Delta = 30'sb111111100100000000000000000000;
		1174: Delta = 30'sb000000011100000000000000000000;
		2388: Delta = 30'sb111111011100000000000000000000;
		1552: Delta = 30'sb000001000100000000000000000000;
		3980: Delta = 30'sb111111000100000000000000000000;
		567: Delta = 30'sb000000111100000000000000000000;
		2995: Delta = 30'sb111110111100000000000000000000;
		338: Delta = 30'sb000010000100000000000000000000;
		647: Delta = 30'sb111110000100000000000000000000;
		3900: Delta = 30'sb000001111100000000000000000000;
		4209: Delta = 30'sb111101111100000000000000000000;
		2457: Delta = 30'sb000100000100000000000000000000;
		3075: Delta = 30'sb111100000100000000000000000000;
		1472: Delta = 30'sb000011111100000000000000000000;
		2090: Delta = 30'sb111011111100000000000000000000;
		2148: Delta = 30'sb001000000100000000000000000000;
		3384: Delta = 30'sb111000000100000000000000000000;
		1163: Delta = 30'sb000111111100000000000000000000;
		2399: Delta = 30'sb110111111100000000000000000000;
		1530: Delta = 30'sb010000000100000000000000000000;
		4002: Delta = 30'sb110000000100000000000000000000;
		545: Delta = 30'sb001111111100000000000000000000;
		3017: Delta = 30'sb101111111100000000000000000000;
		2955: Delta = 30'sb000000011000000000000000000000;
		1592: Delta = 30'sb111111101000000000000000000000;
		378: Delta = 30'sb000000101000000000000000000000;
		4169: Delta = 30'sb111111011000000000000000000000;
		4318: Delta = 30'sb000001001000000000000000000000;
		2199: Delta = 30'sb111111001000000000000000000000;
		2348: Delta = 30'sb000000111000000000000000000000;
		229: Delta = 30'sb111110111000000000000000000000;
		3104: Delta = 30'sb000010001000000000000000000000;
		3413: Delta = 30'sb111110001000000000000000000000;
		1134: Delta = 30'sb000001111000000000000000000000;
		1443: Delta = 30'sb111101111000000000000000000000;
		676: Delta = 30'sb000100001000000000000000000000;
		1294: Delta = 30'sb111100001000000000000000000000;
		3253: Delta = 30'sb000011111000000000000000000000;
		3871: Delta = 30'sb111011111000000000000000000000;
		367: Delta = 30'sb001000001000000000000000000000;
		1603: Delta = 30'sb111000001000000000000000000000;
		2944: Delta = 30'sb000111111000000000000000000000;
		4180: Delta = 30'sb110111111000000000000000000000;
		4296: Delta = 30'sb010000001000000000000000000000;
		2221: Delta = 30'sb110000001000000000000000000000;
		2326: Delta = 30'sb001111111000000000000000000000;
		251: Delta = 30'sb101111111000000000000000000000;
		1363: Delta = 30'sb000000110000000000000000000000;
		3184: Delta = 30'sb111111010000000000000000000000;
		756: Delta = 30'sb000001010000000000000000000000;
		3791: Delta = 30'sb111110110000000000000000000000;
		4089: Delta = 30'sb000010010000000000000000000000;
		4398: Delta = 30'sb111110010000000000000000000000;
		149: Delta = 30'sb000001110000000000000000000000;
		458: Delta = 30'sb111101110000000000000000000000;
		1661: Delta = 30'sb000100010000000000000000000000;
		2279: Delta = 30'sb111100010000000000000000000000;
		2268: Delta = 30'sb000011110000000000000000000000;
		2886: Delta = 30'sb111011110000000000000000000000;
		1352: Delta = 30'sb001000010000000000000000000000;
		2588: Delta = 30'sb111000010000000000000000000000;
		1959: Delta = 30'sb000111110000000000000000000000;
		3195: Delta = 30'sb110111110000000000000000000000;
		734: Delta = 30'sb010000010000000000000000000000;
		3206: Delta = 30'sb110000010000000000000000000000;
		1341: Delta = 30'sb001111110000000000000000000000;
		3813: Delta = 30'sb101111110000000000000000000000;
		2726: Delta = 30'sb000001100000000000000000000000;
		1821: Delta = 30'sb111110100000000000000000000000;
		1512: Delta = 30'sb000010100000000000000000000000;
		3035: Delta = 30'sb111101100000000000000000000000;
		3631: Delta = 30'sb000100100000000000000000000000;
		4249: Delta = 30'sb111100100000000000000000000000;
		298: Delta = 30'sb000011100000000000000000000000;
		916: Delta = 30'sb111011100000000000000000000000;
		3322: Delta = 30'sb001000100000000000000000000000;
		11: Delta = 30'sb111000100000000000000000000000;
		4536: Delta = 30'sb000111100000000000000000000000;
		1225: Delta = 30'sb110111100000000000000000000000;
		2704: Delta = 30'sb010000100000000000000000000000;
		629: Delta = 30'sb110000100000000000000000000000;
		3918: Delta = 30'sb001111100000000000000000000000;
		1843: Delta = 30'sb101111100000000000000000000000;
		905: Delta = 30'sb000011000000000000000000000000;
		3642: Delta = 30'sb111101000000000000000000000000;
		3024: Delta = 30'sb000101000000000000000000000000;
		1523: Delta = 30'sb111011000000000000000000000000;
		2715: Delta = 30'sb001001000000000000000000000000;
		3951: Delta = 30'sb111001000000000000000000000000;
		596: Delta = 30'sb000111000000000000000000000000;
		1832: Delta = 30'sb110111000000000000000000000000;
		2097: Delta = 30'sb010001000000000000000000000000;
		22: Delta = 30'sb110001000000000000000000000000;
		4525: Delta = 30'sb001111000000000000000000000000;
		2450: Delta = 30'sb101111000000000000000000000000;
		1810: Delta = 30'sb000110000000000000000000000000;
		2737: Delta = 30'sb111010000000000000000000000000;
		1501: Delta = 30'sb001010000000000000000000000000;
		3046: Delta = 30'sb110110000000000000000000000000;
		883: Delta = 30'sb010010000000000000000000000000;
		3355: Delta = 30'sb110010000000000000000000000000;
		1192: Delta = 30'sb001110000000000000000000000000;
		3664: Delta = 30'sb101110000000000000000000000000;
		3620: Delta = 30'sb001100000000000000000000000000;
		927: Delta = 30'sb110100000000000000000000000000;
		3002: Delta = 30'sb010100000000000000000000000000;
		1545: Delta = 30'sb101100000000000000000000000000;
		2693: Delta = 30'sb011000000000000000000000000000;
		1854: Delta = 30'sb101000000000000000000000000000;
		default: Delta =30'sb0;
	endcase
end

wire signed [W_BITS-1:0] W_signed;
assign W_signed = (W - Delta);

always@(posedge clk or negedge rst_n) begin
   if(!rst_n) begin
     	ps <= idle;
    end
   else begin
        case(ps)
            idle: begin
                found <= 0;
                R <= 0;
        	Q <= 0;
                ps <= pre;
                end
	    pre: begin
		 Q <= W / A;
		 ps <= load;
		end
            load: begin
                 R <= W - (A * Q);
		 ps <= LUT;
		end
	    LUT: begin
		  if(Delta != 0)begin
		      N <= W_signed / A ;	
		      found <= 1;
                      ps <= idle;
		  end
		  else begin
		      N <= Q;
		      found <= 1;
                      ps <= idle;
		  end
		end
	endcase
    end
end

endmodule


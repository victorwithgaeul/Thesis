`timescale 1ns/1ps
module Tradeoff_52bits(clk, rst_n, W, found, N);

//=========================================================================
//   PARAMETER AND LOCALPARAM FOR FSM
//   W_BITS 要考慮 OVERFLOW 問題
//   N_BITS 也要考慮 OVERFLOW 問題
//=========================================================================
parameter A = 50861 , W_BITS = 69, A_BITS = 16 , N_BITS = 53 , L_BITS = 7;
localparam [2:0] idle=3'b000, pre=3'b001,load=3'b010, lLUT=3'b011, 
                 R2_stage=3'b100, rLUT=3'b101, out=3'b110, done=3'b111;
				 
//==========================================
//   INPUT AND OUTPUT DECLARATION
//==========================================
input clk, rst_n;
input   [W_BITS-1:0]   W;
output reg  [N_BITS-1:0]   N;
output reg  found;

reg [2:0] ps;

//==========================================
//    INSTANTIATE r-LUT l-LUT 
//==========================================
reg [A_BITS-1 :0] R2, R1;

wire signed [L_BITS:0] l_val;
SEC_rLUT52bits rLUT_inst (
    .r(R2),
    .l(l_val) 
);

reg signed [L_BITS:0] h1, h2;
wire  [A_BITS-1:0] r_val;
SEC_lLUT52bits lLUT_inst (
    .l(h1),
    .r(r_val) 
);

//==========================================
//    FUNCTION FOR |h1| |h2| value 
//==========================================
function [L_BITS:0] abs;
    input signed [L_BITS:0] val;
    abs = val[L_BITS] ? ~val + 1 : val;
endfunction

//==========================================
//    FSM for Trade-off Algorithm
//==========================================
reg     [L_BITS:0] H;
reg     s;              // 0 for -1, 1 for +1
reg 	[N_BITS-1:0]	Q;
reg 	[A_BITS-1:0]	R;


wire signed [A_BITS:0] decide;
assign decide = R - R1;

reg [W_BITS-1:0]  W_new;


always@(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        ps <= idle;
        R <= 0;
        Q <= 0;
        found <= 0;
        N <= 0;
        h1 <= 0;
        h2 <= 0;
        R1 <= 0;
        R2 <= 0;
    end
    else begin
        case(ps)
            idle: begin
                found <= 0;
                s <= 0;
                H <= 0;
                ps <= pre;
                end
		pre: begin
		     Q <= W / A;
		     ps <= load;
		   end
            load: begin
                R <= W - (A * Q);
                h1 <= (s == 0) ? -(H + 1) : (H + 1); 
                ps <= lLUT;
                end
            lLUT: begin
                if(R == 0) begin
                    N <= Q;
                    found <= 1;
                    ps <= idle;
                end
                else begin
                    R1 <= r_val;
                    ps <= R2_stage;
                    end
                end
            R2_stage: begin
                R2 <= (decide < 0) ? (decide + A) : (decide);
                ps <= rLUT;
            end
            rLUT: begin
                h2 <= l_val;
                ps <= out;
                end
	    	out: begin
		     W_new <= W - ((s ? 1 : -1) * (1 << (abs(h1) - 1))) - ((h2[L_BITS] ? -1 : 1) * (1 << (abs(h2) - 1)));
		     ps <= done;
		   end
            done: begin
                if(h2 != 0)begin
                   N <= W_new / A ;
                   found <= 1;
                   ps <= idle;
                end
                else begin
                    ps <= load; 
                    if (s == 0) 
                        s <= 1;
                    else begin 
                        s <= 0; 
                        H <= H + 1; 
                    end
                    if (H == (W_BITS - 1) && s == 1) begin
                        ps <= idle;     // not found
                        found <= 1;
                        N <= Q;
                    end
                end
            end
        endcase
    end
end
endmodule

// Product (AN) Code SEC l-LUT
// SEC_lLUT52bits.v
// Received single error location l, output remainder r.
module SEC_lLUT52bits(l, r);
input	signed	[7:0]	l;
output	reg	[15:0]	r;
always@(*) begin
	case(l)
		1: r = 1;
		-1: r = 50860;
		2: r = 2;
		-2: r = 50859;
		3: r = 4;
		-3: r = 50857;
		4: r = 8;
		-4: r = 50853;
		5: r = 16;
		-5: r = 50845;
		6: r = 32;
		-6: r = 50829;
		7: r = 64;
		-7: r = 50797;
		8: r = 128;
		-8: r = 50733;
		9: r = 256;
		-9: r = 50605;
		10: r = 512;
		-10: r = 50349;
		11: r = 1024;
		-11: r = 49837;
		12: r = 2048;
		-12: r = 48813;
		13: r = 4096;
		-13: r = 46765;
		14: r = 8192;
		-14: r = 42669;
		15: r = 16384;
		-15: r = 34477;
		16: r = 32768;
		-16: r = 18093;
		17: r = 14675;
		-17: r = 36186;
		18: r = 29350;
		-18: r = 21511;
		19: r = 7839;
		-19: r = 43022;
		20: r = 15678;
		-20: r = 35183;
		21: r = 31356;
		-21: r = 19505;
		22: r = 11851;
		-22: r = 39010;
		23: r = 23702;
		-23: r = 27159;
		24: r = 47404;
		-24: r = 3457;
		25: r = 43947;
		-25: r = 6914;
		26: r = 37033;
		-26: r = 13828;
		27: r = 23205;
		-27: r = 27656;
		28: r = 46410;
		-28: r = 4451;
		29: r = 41959;
		-29: r = 8902;
		30: r = 33057;
		-30: r = 17804;
		31: r = 15253;
		-31: r = 35608;
		32: r = 30506;
		-32: r = 20355;
		33: r = 10151;
		-33: r = 40710;
		34: r = 20302;
		-34: r = 30559;
		35: r = 40604;
		-35: r = 10257;
		36: r = 30347;
		-36: r = 20514;
		37: r = 9833;
		-37: r = 41028;
		38: r = 19666;
		-38: r = 31195;
		39: r = 39332;
		-39: r = 11529;
		40: r = 27803;
		-40: r = 23058;
		41: r = 4745;
		-41: r = 46116;
		42: r = 9490;
		-42: r = 41371;
		43: r = 18980;
		-43: r = 31881;
		44: r = 37960;
		-44: r = 12901;
		45: r = 25059;
		-45: r = 25802;
		46: r = 50118;
		-46: r = 743;
		47: r = 49375;
		-47: r = 1486;
		48: r = 47889;
		-48: r = 2972;
		49: r = 44917;
		-49: r = 5944;
		50: r = 38973;
		-50: r = 11888;
		51: r = 27085;
		-51: r = 23776;
		52: r = 3309;
		-52: r = 47552;
		53: r = 6618;
		-53: r = 44243;
		54: r = 13236;
		-54: r = 37625;
		55: r = 26472;
		-55: r = 24389;
		56: r = 2083;
		-56: r = 48778;
		57: r = 4166;
		-57: r = 46695;
		58: r = 8332;
		-58: r = 42529;
		59: r = 16664;
		-59: r = 34197;
		60: r = 33328;
		-60: r = 17533;
		61: r = 15795;
		-61: r = 35066;
		62: r = 31590;
		-62: r = 19271;
		63: r = 12319;
		-63: r = 38542;
		64: r = 24638;
		-64: r = 26223;
		65: r = 49276;
		-65: r = 1585;
		66: r = 47691;
		-66: r = 3170;
		67: r = 44521;
		-67: r = 6340;
		68: r = 38181;
		-68: r = 12680;
		default: r = 0;
	endcase
end

endmodule

// Product (AN) Code SEC r-LUT
// SEC_rLUT52bits.v
// Received remainder r, output single error location.
module SEC_rLUT52bits(r, l);
input 	[15:0]	r;
output	reg	signed	[7:0]	l;
always@(*) begin
	case(r)
		1: l = +1;
		50860: l = -1;
		2: l = +2;
		50859: l = -2;
		4: l = +3;
		50857: l = -3;
		8: l = +4;
		50853: l = -4;
		16: l = +5;
		50845: l = -5;
		32: l = +6;
		50829: l = -6;
		64: l = +7;
		50797: l = -7;
		128: l = +8;
		50733: l = -8;
		256: l = +9;
		50605: l = -9;
		512: l = +10;
		50349: l = -10;
		1024: l = +11;
		49837: l = -11;
		2048: l = +12;
		48813: l = -12;
		4096: l = +13;
		46765: l = -13;
		8192: l = +14;
		42669: l = -14;
		16384: l = +15;
		34477: l = -15;
		32768: l = +16;
		18093: l = -16;
		14675: l = +17;
		36186: l = -17;
		29350: l = +18;
		21511: l = -18;
		7839: l = +19;
		43022: l = -19;
		15678: l = +20;
		35183: l = -20;
		31356: l = +21;
		19505: l = -21;
		11851: l = +22;
		39010: l = -22;
		23702: l = +23;
		27159: l = -23;
		47404: l = +24;
		3457: l = -24;
		43947: l = +25;
		6914: l = -25;
		37033: l = +26;
		13828: l = -26;
		23205: l = +27;
		27656: l = -27;
		46410: l = +28;
		4451: l = -28;
		41959: l = +29;
		8902: l = -29;
		33057: l = +30;
		17804: l = -30;
		15253: l = +31;
		35608: l = -31;
		30506: l = +32;
		20355: l = -32;
		10151: l = +33;
		40710: l = -33;
		20302: l = +34;
		30559: l = -34;
		40604: l = +35;
		10257: l = -35;
		30347: l = +36;
		20514: l = -36;
		9833: l = +37;
		41028: l = -37;
		19666: l = +38;
		31195: l = -38;
		39332: l = +39;
		11529: l = -39;
		27803: l = +40;
		23058: l = -40;
		4745: l = +41;
		46116: l = -41;
		9490: l = +42;
		41371: l = -42;
		18980: l = +43;
		31881: l = -43;
		37960: l = +44;
		12901: l = -44;
		25059: l = +45;
		25802: l = -45;
		50118: l = +46;
		743: l = -46;
		49375: l = +47;
		1486: l = -47;
		47889: l = +48;
		2972: l = -48;
		44917: l = +49;
		5944: l = -49;
		38973: l = +50;
		11888: l = -50;
		27085: l = +51;
		23776: l = -51;
		3309: l = +52;
		47552: l = -52;
		6618: l = +53;
		44243: l = -53;
		13236: l = +54;
		37625: l = -54;
		26472: l = +55;
		24389: l = -55;
		2083: l = +56;
		48778: l = -56;
		4166: l = +57;
		46695: l = -57;
		8332: l = +58;
		42529: l = -58;
		16664: l = +59;
		34197: l = -59;
		33328: l = +60;
		17533: l = -60;
		15795: l = +61;
		35066: l = -61;
		31590: l = +62;
		19271: l = -62;
		12319: l = +63;
		38542: l = -63;
		24638: l = +64;
		26223: l = -64;
		49276: l = +65;
		1585: l = -65;
		47691: l = +66;
		3170: l = -66;
		44521: l = +67;
		6340: l = -67;
		38181: l = +68;
		12680: l = -68;
		default: l = 0;
	endcase
end

endmodule


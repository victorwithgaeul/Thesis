// Product (AN) Code DEC_LUT_Decoder
// DEC_LUT_Decoder8bits.v
// Received codeword W = AN + E, E is double AWE (E = e1 + e2), +2^i or -2^i.
module DEC_LUT_Decoder8bits_clk(clk, rst_n, W, found, N);

//=========================================================================
//   W_BITS 要考慮 OVERFLOW 問題 : 19-bits + 2^18 + 2^17
//   N_BITS 也要考慮 OVERFLOW 問題
//=========================================================================
parameter A = 1939 , W_BITS = 20, A_BITS = 11 , N_BITS = 9 , L_BITS = 5;
localparam [1:0] idle=2'b00, pre=2'b01,load=2'b10, LUT=2'b11;

reg [1:0] ps;
//==========================================
//   INPUT AND OUTPUT DECLARATION
//==========================================
input clk, rst_n;
input 	[W_BITS-1:0]	W;
output	reg  [N_BITS-1:0] N;
output  reg  found;

reg 	[N_BITS-1:0]	Q;
reg 	[A_BITS-1:0]	R;

reg   signed	[19:0]	Delta;
always@(*) begin
	case(R)
		1: Delta = 20'sb00000000000000000001;
		1938: Delta = 20'sb11111111111111111111;
		2: Delta = 20'sb00000000000000000010;
		1937: Delta = 20'sb11111111111111111110;
		4: Delta = 20'sb00000000000000000100;
		1935: Delta = 20'sb11111111111111111100;
		8: Delta = 20'sb00000000000000001000;
		1931: Delta = 20'sb11111111111111111000;
		16: Delta = 20'sb00000000000000010000;
		1923: Delta = 20'sb11111111111111110000;
		32: Delta = 20'sb00000000000000100000;
		1907: Delta = 20'sb11111111111111100000;
		64: Delta = 20'sb00000000000001000000;
		1875: Delta = 20'sb11111111111111000000;
		128: Delta = 20'sb00000000000010000000;
		1811: Delta = 20'sb11111111111110000000;
		256: Delta = 20'sb00000000000100000000;
		1683: Delta = 20'sb11111111111100000000;
		512: Delta = 20'sb00000000001000000000;
		1427: Delta = 20'sb11111111111000000000;
		1024: Delta = 20'sb00000000010000000000;
		915: Delta = 20'sb11111111110000000000;
		109: Delta = 20'sb00000000100000000000;
		1830: Delta = 20'sb11111111100000000000;
		218: Delta = 20'sb00000001000000000000;
		1721: Delta = 20'sb11111111000000000000;
		436: Delta = 20'sb00000010000000000000;
		1503: Delta = 20'sb11111110000000000000;
		872: Delta = 20'sb00000100000000000000;
		1067: Delta = 20'sb11111100000000000000;
		1744: Delta = 20'sb00001000000000000000;
		195: Delta = 20'sb11111000000000000000;
		1549: Delta = 20'sb00010000000000000000;
		390: Delta = 20'sb11110000000000000000;
		1159: Delta = 20'sb00100000000000000000;
		780: Delta = 20'sb11100000000000000000;
		379: Delta = 20'sb01000000000000000000;
		1560: Delta = 20'sb11000000000000000000;
		3: Delta = 20'sb00000000000000000011;
		1936: Delta = 20'sb11111111111111111101;
		5: Delta = 20'sb00000000000000000101;
		1934: Delta = 20'sb11111111111111111011;
		9: Delta = 20'sb00000000000000001001;
		1932: Delta = 20'sb11111111111111111001;
		7: Delta = 20'sb00000000000000000111;
		1930: Delta = 20'sb11111111111111110111;
		17: Delta = 20'sb00000000000000010001;
		1924: Delta = 20'sb11111111111111110001;
		15: Delta = 20'sb00000000000000001111;
		1922: Delta = 20'sb11111111111111101111;
		33: Delta = 20'sb00000000000000100001;
		1908: Delta = 20'sb11111111111111100001;
		31: Delta = 20'sb00000000000000011111;
		1906: Delta = 20'sb11111111111111011111;
		65: Delta = 20'sb00000000000001000001;
		1876: Delta = 20'sb11111111111111000001;
		63: Delta = 20'sb00000000000000111111;
		1874: Delta = 20'sb11111111111110111111;
		129: Delta = 20'sb00000000000010000001;
		1812: Delta = 20'sb11111111111110000001;
		127: Delta = 20'sb00000000000001111111;
		1810: Delta = 20'sb11111111111101111111;
		257: Delta = 20'sb00000000000100000001;
		1684: Delta = 20'sb11111111111100000001;
		255: Delta = 20'sb00000000000011111111;
		1682: Delta = 20'sb11111111111011111111;
		513: Delta = 20'sb00000000001000000001;
		1428: Delta = 20'sb11111111111000000001;
		511: Delta = 20'sb00000000000111111111;
		1426: Delta = 20'sb11111111110111111111;
		1025: Delta = 20'sb00000000010000000001;
		916: Delta = 20'sb11111111110000000001;
		1023: Delta = 20'sb00000000001111111111;
		914: Delta = 20'sb11111111101111111111;
		110: Delta = 20'sb00000000100000000001;
		1831: Delta = 20'sb11111111100000000001;
		108: Delta = 20'sb00000000011111111111;
		1829: Delta = 20'sb11111111011111111111;
		219: Delta = 20'sb00000001000000000001;
		1722: Delta = 20'sb11111111000000000001;
		217: Delta = 20'sb00000000111111111111;
		1720: Delta = 20'sb11111110111111111111;
		437: Delta = 20'sb00000010000000000001;
		1504: Delta = 20'sb11111110000000000001;
		435: Delta = 20'sb00000001111111111111;
		1502: Delta = 20'sb11111101111111111111;
		873: Delta = 20'sb00000100000000000001;
		1068: Delta = 20'sb11111100000000000001;
		871: Delta = 20'sb00000011111111111111;
		1066: Delta = 20'sb11111011111111111111;
		1745: Delta = 20'sb00001000000000000001;
		196: Delta = 20'sb11111000000000000001;
		1743: Delta = 20'sb00000111111111111111;
		194: Delta = 20'sb11110111111111111111;
		1550: Delta = 20'sb00010000000000000001;
		391: Delta = 20'sb11110000000000000001;
		1548: Delta = 20'sb00001111111111111111;
		389: Delta = 20'sb11101111111111111111;
		1160: Delta = 20'sb00100000000000000001;
		781: Delta = 20'sb11100000000000000001;
		1158: Delta = 20'sb00011111111111111111;
		779: Delta = 20'sb11011111111111111111;
		380: Delta = 20'sb01000000000000000001;
		1561: Delta = 20'sb11000000000000000001;
		378: Delta = 20'sb00111111111111111111;
		1559: Delta = 20'sb10111111111111111111;
		6: Delta = 20'sb00000000000000000110;
		1933: Delta = 20'sb11111111111111111010;
		10: Delta = 20'sb00000000000000001010;
		1929: Delta = 20'sb11111111111111110110;
		18: Delta = 20'sb00000000000000010010;
		1925: Delta = 20'sb11111111111111110010;
		14: Delta = 20'sb00000000000000001110;
		1921: Delta = 20'sb11111111111111101110;
		34: Delta = 20'sb00000000000000100010;
		1909: Delta = 20'sb11111111111111100010;
		30: Delta = 20'sb00000000000000011110;
		1905: Delta = 20'sb11111111111111011110;
		66: Delta = 20'sb00000000000001000010;
		1877: Delta = 20'sb11111111111111000010;
		62: Delta = 20'sb00000000000000111110;
		1873: Delta = 20'sb11111111111110111110;
		130: Delta = 20'sb00000000000010000010;
		1813: Delta = 20'sb11111111111110000010;
		126: Delta = 20'sb00000000000001111110;
		1809: Delta = 20'sb11111111111101111110;
		258: Delta = 20'sb00000000000100000010;
		1685: Delta = 20'sb11111111111100000010;
		254: Delta = 20'sb00000000000011111110;
		1681: Delta = 20'sb11111111111011111110;
		514: Delta = 20'sb00000000001000000010;
		1429: Delta = 20'sb11111111111000000010;
		510: Delta = 20'sb00000000000111111110;
		1425: Delta = 20'sb11111111110111111110;
		1026: Delta = 20'sb00000000010000000010;
		917: Delta = 20'sb11111111110000000010;
		1022: Delta = 20'sb00000000001111111110;
		913: Delta = 20'sb11111111101111111110;
		111: Delta = 20'sb00000000100000000010;
		1832: Delta = 20'sb11111111100000000010;
		107: Delta = 20'sb00000000011111111110;
		1828: Delta = 20'sb11111111011111111110;
		220: Delta = 20'sb00000001000000000010;
		1723: Delta = 20'sb11111111000000000010;
		216: Delta = 20'sb00000000111111111110;
		1719: Delta = 20'sb11111110111111111110;
		438: Delta = 20'sb00000010000000000010;
		1505: Delta = 20'sb11111110000000000010;
		434: Delta = 20'sb00000001111111111110;
		1501: Delta = 20'sb11111101111111111110;
		874: Delta = 20'sb00000100000000000010;
		1069: Delta = 20'sb11111100000000000010;
		870: Delta = 20'sb00000011111111111110;
		1065: Delta = 20'sb11111011111111111110;
		1746: Delta = 20'sb00001000000000000010;
		197: Delta = 20'sb11111000000000000010;
		1742: Delta = 20'sb00000111111111111110;
		193: Delta = 20'sb11110111111111111110;
		1551: Delta = 20'sb00010000000000000010;
		392: Delta = 20'sb11110000000000000010;
		1547: Delta = 20'sb00001111111111111110;
		388: Delta = 20'sb11101111111111111110;
		1161: Delta = 20'sb00100000000000000010;
		782: Delta = 20'sb11100000000000000010;
		1157: Delta = 20'sb00011111111111111110;
		778: Delta = 20'sb11011111111111111110;
		381: Delta = 20'sb01000000000000000010;
		1562: Delta = 20'sb11000000000000000010;
		377: Delta = 20'sb00111111111111111110;
		1558: Delta = 20'sb10111111111111111110;
		12: Delta = 20'sb00000000000000001100;
		1927: Delta = 20'sb11111111111111110100;
		20: Delta = 20'sb00000000000000010100;
		1919: Delta = 20'sb11111111111111101100;
		36: Delta = 20'sb00000000000000100100;
		1911: Delta = 20'sb11111111111111100100;
		28: Delta = 20'sb00000000000000011100;
		1903: Delta = 20'sb11111111111111011100;
		68: Delta = 20'sb00000000000001000100;
		1879: Delta = 20'sb11111111111111000100;
		60: Delta = 20'sb00000000000000111100;
		1871: Delta = 20'sb11111111111110111100;
		132: Delta = 20'sb00000000000010000100;
		1815: Delta = 20'sb11111111111110000100;
		124: Delta = 20'sb00000000000001111100;
		1807: Delta = 20'sb11111111111101111100;
		260: Delta = 20'sb00000000000100000100;
		1687: Delta = 20'sb11111111111100000100;
		252: Delta = 20'sb00000000000011111100;
		1679: Delta = 20'sb11111111111011111100;
		516: Delta = 20'sb00000000001000000100;
		1431: Delta = 20'sb11111111111000000100;
		508: Delta = 20'sb00000000000111111100;
		1423: Delta = 20'sb11111111110111111100;
		1028: Delta = 20'sb00000000010000000100;
		919: Delta = 20'sb11111111110000000100;
		1020: Delta = 20'sb00000000001111111100;
		911: Delta = 20'sb11111111101111111100;
		113: Delta = 20'sb00000000100000000100;
		1834: Delta = 20'sb11111111100000000100;
		105: Delta = 20'sb00000000011111111100;
		1826: Delta = 20'sb11111111011111111100;
		222: Delta = 20'sb00000001000000000100;
		1725: Delta = 20'sb11111111000000000100;
		214: Delta = 20'sb00000000111111111100;
		1717: Delta = 20'sb11111110111111111100;
		440: Delta = 20'sb00000010000000000100;
		1507: Delta = 20'sb11111110000000000100;
		432: Delta = 20'sb00000001111111111100;
		1499: Delta = 20'sb11111101111111111100;
		876: Delta = 20'sb00000100000000000100;
		1071: Delta = 20'sb11111100000000000100;
		868: Delta = 20'sb00000011111111111100;
		1063: Delta = 20'sb11111011111111111100;
		1748: Delta = 20'sb00001000000000000100;
		199: Delta = 20'sb11111000000000000100;
		1740: Delta = 20'sb00000111111111111100;
		191: Delta = 20'sb11110111111111111100;
		1553: Delta = 20'sb00010000000000000100;
		394: Delta = 20'sb11110000000000000100;
		1545: Delta = 20'sb00001111111111111100;
		386: Delta = 20'sb11101111111111111100;
		1163: Delta = 20'sb00100000000000000100;
		784: Delta = 20'sb11100000000000000100;
		1155: Delta = 20'sb00011111111111111100;
		776: Delta = 20'sb11011111111111111100;
		383: Delta = 20'sb01000000000000000100;
		1564: Delta = 20'sb11000000000000000100;
		375: Delta = 20'sb00111111111111111100;
		1556: Delta = 20'sb10111111111111111100;
		24: Delta = 20'sb00000000000000011000;
		1915: Delta = 20'sb11111111111111101000;
		40: Delta = 20'sb00000000000000101000;
		1899: Delta = 20'sb11111111111111011000;
		72: Delta = 20'sb00000000000001001000;
		1883: Delta = 20'sb11111111111111001000;
		56: Delta = 20'sb00000000000000111000;
		1867: Delta = 20'sb11111111111110111000;
		136: Delta = 20'sb00000000000010001000;
		1819: Delta = 20'sb11111111111110001000;
		120: Delta = 20'sb00000000000001111000;
		1803: Delta = 20'sb11111111111101111000;
		264: Delta = 20'sb00000000000100001000;
		1691: Delta = 20'sb11111111111100001000;
		248: Delta = 20'sb00000000000011111000;
		1675: Delta = 20'sb11111111111011111000;
		520: Delta = 20'sb00000000001000001000;
		1435: Delta = 20'sb11111111111000001000;
		504: Delta = 20'sb00000000000111111000;
		1419: Delta = 20'sb11111111110111111000;
		1032: Delta = 20'sb00000000010000001000;
		923: Delta = 20'sb11111111110000001000;
		1016: Delta = 20'sb00000000001111111000;
		907: Delta = 20'sb11111111101111111000;
		117: Delta = 20'sb00000000100000001000;
		1838: Delta = 20'sb11111111100000001000;
		101: Delta = 20'sb00000000011111111000;
		1822: Delta = 20'sb11111111011111111000;
		226: Delta = 20'sb00000001000000001000;
		1729: Delta = 20'sb11111111000000001000;
		210: Delta = 20'sb00000000111111111000;
		1713: Delta = 20'sb11111110111111111000;
		444: Delta = 20'sb00000010000000001000;
		1511: Delta = 20'sb11111110000000001000;
		428: Delta = 20'sb00000001111111111000;
		1495: Delta = 20'sb11111101111111111000;
		880: Delta = 20'sb00000100000000001000;
		1075: Delta = 20'sb11111100000000001000;
		864: Delta = 20'sb00000011111111111000;
		1059: Delta = 20'sb11111011111111111000;
		1752: Delta = 20'sb00001000000000001000;
		203: Delta = 20'sb11111000000000001000;
		1736: Delta = 20'sb00000111111111111000;
		187: Delta = 20'sb11110111111111111000;
		1557: Delta = 20'sb00010000000000001000;
		398: Delta = 20'sb11110000000000001000;
		1541: Delta = 20'sb00001111111111111000;
		382: Delta = 20'sb11101111111111111000;
		1167: Delta = 20'sb00100000000000001000;
		788: Delta = 20'sb11100000000000001000;
		1151: Delta = 20'sb00011111111111111000;
		772: Delta = 20'sb11011111111111111000;
		387: Delta = 20'sb01000000000000001000;
		1568: Delta = 20'sb11000000000000001000;
		371: Delta = 20'sb00111111111111111000;
		1552: Delta = 20'sb10111111111111111000;
		48: Delta = 20'sb00000000000000110000;
		1891: Delta = 20'sb11111111111111010000;
		80: Delta = 20'sb00000000000001010000;
		1859: Delta = 20'sb11111111111110110000;
		144: Delta = 20'sb00000000000010010000;
		1827: Delta = 20'sb11111111111110010000;
		112: Delta = 20'sb00000000000001110000;
		1795: Delta = 20'sb11111111111101110000;
		272: Delta = 20'sb00000000000100010000;
		1699: Delta = 20'sb11111111111100010000;
		240: Delta = 20'sb00000000000011110000;
		1667: Delta = 20'sb11111111111011110000;
		528: Delta = 20'sb00000000001000010000;
		1443: Delta = 20'sb11111111111000010000;
		496: Delta = 20'sb00000000000111110000;
		1411: Delta = 20'sb11111111110111110000;
		1040: Delta = 20'sb00000000010000010000;
		931: Delta = 20'sb11111111110000010000;
		1008: Delta = 20'sb00000000001111110000;
		899: Delta = 20'sb11111111101111110000;
		125: Delta = 20'sb00000000100000010000;
		1846: Delta = 20'sb11111111100000010000;
		93: Delta = 20'sb00000000011111110000;
		1814: Delta = 20'sb11111111011111110000;
		234: Delta = 20'sb00000001000000010000;
		1737: Delta = 20'sb11111111000000010000;
		202: Delta = 20'sb00000000111111110000;
		1705: Delta = 20'sb11111110111111110000;
		452: Delta = 20'sb00000010000000010000;
		1519: Delta = 20'sb11111110000000010000;
		420: Delta = 20'sb00000001111111110000;
		1487: Delta = 20'sb11111101111111110000;
		888: Delta = 20'sb00000100000000010000;
		1083: Delta = 20'sb11111100000000010000;
		856: Delta = 20'sb00000011111111110000;
		1051: Delta = 20'sb11111011111111110000;
		1760: Delta = 20'sb00001000000000010000;
		211: Delta = 20'sb11111000000000010000;
		1728: Delta = 20'sb00000111111111110000;
		179: Delta = 20'sb11110111111111110000;
		1565: Delta = 20'sb00010000000000010000;
		406: Delta = 20'sb11110000000000010000;
		1533: Delta = 20'sb00001111111111110000;
		374: Delta = 20'sb11101111111111110000;
		1175: Delta = 20'sb00100000000000010000;
		796: Delta = 20'sb11100000000000010000;
		1143: Delta = 20'sb00011111111111110000;
		764: Delta = 20'sb11011111111111110000;
		395: Delta = 20'sb01000000000000010000;
		1576: Delta = 20'sb11000000000000010000;
		363: Delta = 20'sb00111111111111110000;
		1544: Delta = 20'sb10111111111111110000;
		96: Delta = 20'sb00000000000001100000;
		1843: Delta = 20'sb11111111111110100000;
		160: Delta = 20'sb00000000000010100000;
		1779: Delta = 20'sb11111111111101100000;
		288: Delta = 20'sb00000000000100100000;
		1715: Delta = 20'sb11111111111100100000;
		224: Delta = 20'sb00000000000011100000;
		1651: Delta = 20'sb11111111111011100000;
		544: Delta = 20'sb00000000001000100000;
		1459: Delta = 20'sb11111111111000100000;
		480: Delta = 20'sb00000000000111100000;
		1395: Delta = 20'sb11111111110111100000;
		1056: Delta = 20'sb00000000010000100000;
		947: Delta = 20'sb11111111110000100000;
		992: Delta = 20'sb00000000001111100000;
		883: Delta = 20'sb11111111101111100000;
		141: Delta = 20'sb00000000100000100000;
		1862: Delta = 20'sb11111111100000100000;
		77: Delta = 20'sb00000000011111100000;
		1798: Delta = 20'sb11111111011111100000;
		250: Delta = 20'sb00000001000000100000;
		1753: Delta = 20'sb11111111000000100000;
		186: Delta = 20'sb00000000111111100000;
		1689: Delta = 20'sb11111110111111100000;
		468: Delta = 20'sb00000010000000100000;
		1535: Delta = 20'sb11111110000000100000;
		404: Delta = 20'sb00000001111111100000;
		1471: Delta = 20'sb11111101111111100000;
		904: Delta = 20'sb00000100000000100000;
		1099: Delta = 20'sb11111100000000100000;
		840: Delta = 20'sb00000011111111100000;
		1035: Delta = 20'sb11111011111111100000;
		1776: Delta = 20'sb00001000000000100000;
		227: Delta = 20'sb11111000000000100000;
		1712: Delta = 20'sb00000111111111100000;
		163: Delta = 20'sb11110111111111100000;
		1581: Delta = 20'sb00010000000000100000;
		422: Delta = 20'sb11110000000000100000;
		1517: Delta = 20'sb00001111111111100000;
		358: Delta = 20'sb11101111111111100000;
		1191: Delta = 20'sb00100000000000100000;
		812: Delta = 20'sb11100000000000100000;
		1127: Delta = 20'sb00011111111111100000;
		748: Delta = 20'sb11011111111111100000;
		411: Delta = 20'sb01000000000000100000;
		1592: Delta = 20'sb11000000000000100000;
		347: Delta = 20'sb00111111111111100000;
		1528: Delta = 20'sb10111111111111100000;
		192: Delta = 20'sb00000000000011000000;
		1747: Delta = 20'sb11111111111101000000;
		320: Delta = 20'sb00000000000101000000;
		1619: Delta = 20'sb11111111111011000000;
		576: Delta = 20'sb00000000001001000000;
		1491: Delta = 20'sb11111111111001000000;
		448: Delta = 20'sb00000000000111000000;
		1363: Delta = 20'sb11111111110111000000;
		1088: Delta = 20'sb00000000010001000000;
		979: Delta = 20'sb11111111110001000000;
		960: Delta = 20'sb00000000001111000000;
		851: Delta = 20'sb11111111101111000000;
		173: Delta = 20'sb00000000100001000000;
		1894: Delta = 20'sb11111111100001000000;
		45: Delta = 20'sb00000000011111000000;
		1766: Delta = 20'sb11111111011111000000;
		282: Delta = 20'sb00000001000001000000;
		1785: Delta = 20'sb11111111000001000000;
		154: Delta = 20'sb00000000111111000000;
		1657: Delta = 20'sb11111110111111000000;
		500: Delta = 20'sb00000010000001000000;
		1567: Delta = 20'sb11111110000001000000;
		372: Delta = 20'sb00000001111111000000;
		1439: Delta = 20'sb11111101111111000000;
		936: Delta = 20'sb00000100000001000000;
		1131: Delta = 20'sb11111100000001000000;
		808: Delta = 20'sb00000011111111000000;
		1003: Delta = 20'sb11111011111111000000;
		1808: Delta = 20'sb00001000000001000000;
		259: Delta = 20'sb11111000000001000000;
		1680: Delta = 20'sb00000111111111000000;
		131: Delta = 20'sb11110111111111000000;
		1613: Delta = 20'sb00010000000001000000;
		454: Delta = 20'sb11110000000001000000;
		1485: Delta = 20'sb00001111111111000000;
		326: Delta = 20'sb11101111111111000000;
		1223: Delta = 20'sb00100000000001000000;
		844: Delta = 20'sb11100000000001000000;
		1095: Delta = 20'sb00011111111111000000;
		716: Delta = 20'sb11011111111111000000;
		443: Delta = 20'sb01000000000001000000;
		1624: Delta = 20'sb11000000000001000000;
		315: Delta = 20'sb00111111111111000000;
		1496: Delta = 20'sb10111111111111000000;
		384: Delta = 20'sb00000000000110000000;
		1555: Delta = 20'sb11111111111010000000;
		640: Delta = 20'sb00000000001010000000;
		1299: Delta = 20'sb11111111110110000000;
		1152: Delta = 20'sb00000000010010000000;
		1043: Delta = 20'sb11111111110010000000;
		896: Delta = 20'sb00000000001110000000;
		787: Delta = 20'sb11111111101110000000;
		237: Delta = 20'sb00000000100010000000;
		19: Delta = 20'sb11111111100010000000;
		1920: Delta = 20'sb00000000011110000000;
		1702: Delta = 20'sb11111111011110000000;
		346: Delta = 20'sb00000001000010000000;
		1849: Delta = 20'sb11111111000010000000;
		90: Delta = 20'sb00000000111110000000;
		1593: Delta = 20'sb11111110111110000000;
		564: Delta = 20'sb00000010000010000000;
		1631: Delta = 20'sb11111110000010000000;
		308: Delta = 20'sb00000001111110000000;
		1375: Delta = 20'sb11111101111110000000;
		1000: Delta = 20'sb00000100000010000000;
		1195: Delta = 20'sb11111100000010000000;
		744: Delta = 20'sb00000011111110000000;
		939: Delta = 20'sb11111011111110000000;
		1872: Delta = 20'sb00001000000010000000;
		323: Delta = 20'sb11111000000010000000;
		1616: Delta = 20'sb00000111111110000000;
		67: Delta = 20'sb11110111111110000000;
		1677: Delta = 20'sb00010000000010000000;
		518: Delta = 20'sb11110000000010000000;
		1421: Delta = 20'sb00001111111110000000;
		262: Delta = 20'sb11101111111110000000;
		1287: Delta = 20'sb00100000000010000000;
		908: Delta = 20'sb11100000000010000000;
		1031: Delta = 20'sb00011111111110000000;
		652: Delta = 20'sb11011111111110000000;
		507: Delta = 20'sb01000000000010000000;
		1688: Delta = 20'sb11000000000010000000;
		251: Delta = 20'sb00111111111110000000;
		1432: Delta = 20'sb10111111111110000000;
		768: Delta = 20'sb00000000001100000000;
		1171: Delta = 20'sb11111111110100000000;
		1280: Delta = 20'sb00000000010100000000;
		659: Delta = 20'sb11111111101100000000;
		365: Delta = 20'sb00000000100100000000;
		147: Delta = 20'sb11111111100100000000;
		1792: Delta = 20'sb00000000011100000000;
		1574: Delta = 20'sb11111111011100000000;
		474: Delta = 20'sb00000001000100000000;
		38: Delta = 20'sb11111111000100000000;
		1901: Delta = 20'sb00000000111100000000;
		1465: Delta = 20'sb11111110111100000000;
		692: Delta = 20'sb00000010000100000000;
		1759: Delta = 20'sb11111110000100000000;
		180: Delta = 20'sb00000001111100000000;
		1247: Delta = 20'sb11111101111100000000;
		1128: Delta = 20'sb00000100000100000000;
		1323: Delta = 20'sb11111100000100000000;
		616: Delta = 20'sb00000011111100000000;
		811: Delta = 20'sb11111011111100000000;
		61: Delta = 20'sb00001000000100000000;
		451: Delta = 20'sb11111000000100000000;
		1488: Delta = 20'sb00000111111100000000;
		1878: Delta = 20'sb11110111111100000000;
		1805: Delta = 20'sb00010000000100000000;
		646: Delta = 20'sb11110000000100000000;
		1293: Delta = 20'sb00001111111100000000;
		134: Delta = 20'sb11101111111100000000;
		1415: Delta = 20'sb00100000000100000000;
		1036: Delta = 20'sb11100000000100000000;
		903: Delta = 20'sb00011111111100000000;
		524: Delta = 20'sb11011111111100000000;
		635: Delta = 20'sb01000000000100000000;
		1816: Delta = 20'sb11000000000100000000;
		123: Delta = 20'sb00111111111100000000;
		1304: Delta = 20'sb10111111111100000000;
		1536: Delta = 20'sb00000000011000000000;
		403: Delta = 20'sb11111111101000000000;
		621: Delta = 20'sb00000000101000000000;
		1318: Delta = 20'sb11111111011000000000;
		730: Delta = 20'sb00000001001000000000;
		294: Delta = 20'sb11111111001000000000;
		1645: Delta = 20'sb00000000111000000000;
		1209: Delta = 20'sb11111110111000000000;
		948: Delta = 20'sb00000010001000000000;
		76: Delta = 20'sb11111110001000000000;
		1863: Delta = 20'sb00000001111000000000;
		991: Delta = 20'sb11111101111000000000;
		1384: Delta = 20'sb00000100001000000000;
		1579: Delta = 20'sb11111100001000000000;
		360: Delta = 20'sb00000011111000000000;
		555: Delta = 20'sb11111011111000000000;
		317: Delta = 20'sb00001000001000000000;
		707: Delta = 20'sb11111000001000000000;
		1232: Delta = 20'sb00000111111000000000;
		1622: Delta = 20'sb11110111111000000000;
		122: Delta = 20'sb00010000001000000000;
		902: Delta = 20'sb11110000001000000000;
		1037: Delta = 20'sb00001111111000000000;
		1817: Delta = 20'sb11101111111000000000;
		1671: Delta = 20'sb00100000001000000000;
		1292: Delta = 20'sb11100000001000000000;
		647: Delta = 20'sb00011111111000000000;
		268: Delta = 20'sb11011111111000000000;
		891: Delta = 20'sb01000000001000000000;
		133: Delta = 20'sb11000000001000000000;
		1806: Delta = 20'sb00111111111000000000;
		1048: Delta = 20'sb10111111111000000000;
		1133: Delta = 20'sb00000000110000000000;
		806: Delta = 20'sb11111111010000000000;
		1242: Delta = 20'sb00000001010000000000;
		697: Delta = 20'sb11111110110000000000;
		1460: Delta = 20'sb00000010010000000000;
		588: Delta = 20'sb11111110010000000000;
		1351: Delta = 20'sb00000001110000000000;
		479: Delta = 20'sb11111101110000000000;
		1896: Delta = 20'sb00000100010000000000;
		152: Delta = 20'sb11111100010000000000;
		1787: Delta = 20'sb00000011110000000000;
		43: Delta = 20'sb11111011110000000000;
		829: Delta = 20'sb00001000010000000000;
		1219: Delta = 20'sb11111000010000000000;
		720: Delta = 20'sb00000111110000000000;
		1110: Delta = 20'sb11110111110000000000;
		634: Delta = 20'sb00010000010000000000;
		1414: Delta = 20'sb11110000010000000000;
		525: Delta = 20'sb00001111110000000000;
		1305: Delta = 20'sb11101111110000000000;
		244: Delta = 20'sb00100000010000000000;
		1804: Delta = 20'sb11100000010000000000;
		135: Delta = 20'sb00011111110000000000;
		1695: Delta = 20'sb11011111110000000000;
		1403: Delta = 20'sb01000000010000000000;
		645: Delta = 20'sb11000000010000000000;
		1294: Delta = 20'sb00111111110000000000;
		536: Delta = 20'sb10111111110000000000;
		327: Delta = 20'sb00000001100000000000;
		1612: Delta = 20'sb11111110100000000000;
		545: Delta = 20'sb00000010100000000000;
		1394: Delta = 20'sb11111101100000000000;
		981: Delta = 20'sb00000100100000000000;
		1176: Delta = 20'sb11111100100000000000;
		763: Delta = 20'sb00000011100000000000;
		958: Delta = 20'sb11111011100000000000;
		1853: Delta = 20'sb00001000100000000000;
		304: Delta = 20'sb11111000100000000000;
		1635: Delta = 20'sb00000111100000000000;
		86: Delta = 20'sb11110111100000000000;
		1658: Delta = 20'sb00010000100000000000;
		499: Delta = 20'sb11110000100000000000;
		1440: Delta = 20'sb00001111100000000000;
		281: Delta = 20'sb11101111100000000000;
		1268: Delta = 20'sb00100000100000000000;
		889: Delta = 20'sb11100000100000000000;
		1050: Delta = 20'sb00011111100000000000;
		671: Delta = 20'sb11011111100000000000;
		488: Delta = 20'sb01000000100000000000;
		1669: Delta = 20'sb11000000100000000000;
		270: Delta = 20'sb00111111100000000000;
		1451: Delta = 20'sb10111111100000000000;
		654: Delta = 20'sb00000011000000000000;
		1285: Delta = 20'sb11111101000000000000;
		1090: Delta = 20'sb00000101000000000000;
		849: Delta = 20'sb11111011000000000000;
		23: Delta = 20'sb00001001000000000000;
		413: Delta = 20'sb11111001000000000000;
		1526: Delta = 20'sb00000111000000000000;
		1916: Delta = 20'sb11110111000000000000;
		1767: Delta = 20'sb00010001000000000000;
		608: Delta = 20'sb11110001000000000000;
		1331: Delta = 20'sb00001111000000000000;
		172: Delta = 20'sb11101111000000000000;
		1377: Delta = 20'sb00100001000000000000;
		998: Delta = 20'sb11100001000000000000;
		941: Delta = 20'sb00011111000000000000;
		562: Delta = 20'sb11011111000000000000;
		597: Delta = 20'sb01000001000000000000;
		1778: Delta = 20'sb11000001000000000000;
		161: Delta = 20'sb00111111000000000000;
		1342: Delta = 20'sb10111111000000000000;
		1308: Delta = 20'sb00000110000000000000;
		631: Delta = 20'sb11111010000000000000;
		241: Delta = 20'sb00001010000000000000;
		1698: Delta = 20'sb11110110000000000000;
		46: Delta = 20'sb00010010000000000000;
		826: Delta = 20'sb11110010000000000000;
		1113: Delta = 20'sb00001110000000000000;
		1893: Delta = 20'sb11101110000000000000;
		1595: Delta = 20'sb00100010000000000000;
		1216: Delta = 20'sb11100010000000000000;
		723: Delta = 20'sb00011110000000000000;
		344: Delta = 20'sb11011110000000000000;
		815: Delta = 20'sb01000010000000000000;
		57: Delta = 20'sb11000010000000000000;
		1882: Delta = 20'sb00111110000000000000;
		1124: Delta = 20'sb10111110000000000000;
		677: Delta = 20'sb00001100000000000000;
		1262: Delta = 20'sb11110100000000000000;
		482: Delta = 20'sb00010100000000000000;
		1457: Delta = 20'sb11101100000000000000;
		92: Delta = 20'sb00100100000000000000;
		1652: Delta = 20'sb11100100000000000000;
		287: Delta = 20'sb00011100000000000000;
		1847: Delta = 20'sb11011100000000000000;
		1251: Delta = 20'sb01000100000000000000;
		493: Delta = 20'sb11000100000000000000;
		1446: Delta = 20'sb00111100000000000000;
		688: Delta = 20'sb10111100000000000000;
		1354: Delta = 20'sb00011000000000000000;
		585: Delta = 20'sb11101000000000000000;
		964: Delta = 20'sb00101000000000000000;
		975: Delta = 20'sb11011000000000000000;
		184: Delta = 20'sb01001000000000000000;
		1365: Delta = 20'sb11001000000000000000;
		574: Delta = 20'sb00111000000000000000;
		1755: Delta = 20'sb10111000000000000000;
		769: Delta = 20'sb00110000000000000000;
		1170: Delta = 20'sb11010000000000000000;
		1928: Delta = 20'sb01010000000000000000;
		11: Delta = 20'sb10110000000000000000;
		1538: Delta = 20'sb01100000000000000000;
		401: Delta = 20'sb10100000000000000000;
		default: Delta =20'sb0;
	endcase
end

wire signed [W_BITS-1:0] W_signed;
assign W_signed = (W - Delta);

always@(posedge clk or negedge rst_n) begin
   if(!rst_n) begin
     	ps <= idle;
    end
   else begin
        case(ps)
            idle: begin
                found <= 0;
                R <= 0;
        	Q <= 0;
                ps <= pre;
                end
	    pre: begin
		 Q <= W / A;
		 ps <= load;
		end
            load: begin
                 R <= W - (A * Q);
		 ps <= LUT;
		end
	    LUT: begin
		  if(Delta != 0)begin
		      N <= W_signed / A ;	
		      found <= 1;
                      ps <= idle;
		  end
		  else begin
		      N <= Q;
		      found <= 1;
                      ps <= idle;
		  end
		end
	endcase
    end
end

endmodule


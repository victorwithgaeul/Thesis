// Product (AN) Code DEC r-LUT
// DEC_rLUT20bits.v
// Used to do DEC, but corrected errors by locations, not AWE
// Received remainder r, output two error locations.
module DEC_rLUT20bits(r, l_1, l_2);
input 	[12:0]	r;
output	reg	signed	[6:0]	l_1;
output	reg	signed	[6:0]	l_2;
always@(*) begin
	case(r)
		1: begin l_1 = -1;
				 l_2 = +2; end
		6310: begin l_1 = +1;
				 l_2 = -2; end
		2: begin l_1 = +1;
				 l_2 = +1; end
		6309: begin l_1 = -1;
				 l_2 = -1; end
		4: begin l_1 = +2;
				 l_2 = +2; end
		6307: begin l_1 = -2;
				 l_2 = -2; end
		8: begin l_1 = +3;
				 l_2 = +3; end
		6303: begin l_1 = -3;
				 l_2 = -3; end
		16: begin l_1 = +4;
				 l_2 = +4; end
		6295: begin l_1 = -4;
				 l_2 = -4; end
		32: begin l_1 = +5;
				 l_2 = +5; end
		6279: begin l_1 = -5;
				 l_2 = -5; end
		64: begin l_1 = +6;
				 l_2 = +6; end
		6247: begin l_1 = -6;
				 l_2 = -6; end
		128: begin l_1 = +7;
				 l_2 = +7; end
		6183: begin l_1 = -7;
				 l_2 = -7; end
		256: begin l_1 = +8;
				 l_2 = +8; end
		6055: begin l_1 = -8;
				 l_2 = -8; end
		512: begin l_1 = +9;
				 l_2 = +9; end
		5799: begin l_1 = -9;
				 l_2 = -9; end
		1024: begin l_1 = +10;
				 l_2 = +10; end
		5287: begin l_1 = -10;
				 l_2 = -10; end
		2048: begin l_1 = +11;
				 l_2 = +11; end
		4263: begin l_1 = -11;
				 l_2 = -11; end
		4096: begin l_1 = +12;
				 l_2 = +12; end
		2215: begin l_1 = -12;
				 l_2 = -12; end
		1881: begin l_1 = +13;
				 l_2 = +13; end
		4430: begin l_1 = -13;
				 l_2 = -13; end
		3762: begin l_1 = +14;
				 l_2 = +14; end
		2549: begin l_1 = -14;
				 l_2 = -14; end
		1213: begin l_1 = +15;
				 l_2 = +15; end
		5098: begin l_1 = -15;
				 l_2 = -15; end
		2426: begin l_1 = +16;
				 l_2 = +16; end
		3885: begin l_1 = -16;
				 l_2 = -16; end
		4852: begin l_1 = +17;
				 l_2 = +17; end
		1459: begin l_1 = -17;
				 l_2 = -17; end
		3393: begin l_1 = +18;
				 l_2 = +18; end
		2918: begin l_1 = -18;
				 l_2 = -18; end
		475: begin l_1 = +19;
				 l_2 = +19; end
		5836: begin l_1 = -19;
				 l_2 = -19; end
		950: begin l_1 = +20;
				 l_2 = +20; end
		5361: begin l_1 = -20;
				 l_2 = -20; end
		1900: begin l_1 = +21;
				 l_2 = +21; end
		4411: begin l_1 = -21;
				 l_2 = -21; end
		3800: begin l_1 = +22;
				 l_2 = +22; end
		2511: begin l_1 = -22;
				 l_2 = -22; end
		1289: begin l_1 = +23;
				 l_2 = +23; end
		5022: begin l_1 = -23;
				 l_2 = -23; end
		2578: begin l_1 = +24;
				 l_2 = +24; end
		3733: begin l_1 = -24;
				 l_2 = -24; end
		5156: begin l_1 = +25;
				 l_2 = +25; end
		1155: begin l_1 = -25;
				 l_2 = -25; end
		4001: begin l_1 = +26;
				 l_2 = +26; end
		2310: begin l_1 = -26;
				 l_2 = -26; end
		1691: begin l_1 = +27;
				 l_2 = +27; end
		4620: begin l_1 = -27;
				 l_2 = -27; end
		3382: begin l_1 = +28;
				 l_2 = +28; end
		2929: begin l_1 = -28;
				 l_2 = -28; end
		453: begin l_1 = +29;
				 l_2 = +29; end
		5858: begin l_1 = -29;
				 l_2 = -29; end
		906: begin l_1 = +30;
				 l_2 = +30; end
		5405: begin l_1 = -30;
				 l_2 = -30; end
		1812: begin l_1 = +31;
				 l_2 = +31; end
		4499: begin l_1 = -31;
				 l_2 = -31; end
		3624: begin l_1 = +32;
				 l_2 = +32; end
		2687: begin l_1 = -32;
				 l_2 = -32; end
		3: begin l_1 = -1;
				 l_2 = +3; end
		6308: begin l_1 = -1;
				 l_2 = -2; end
		5: begin l_1 = +1;
				 l_2 = +3; end
		6306: begin l_1 = -1;
				 l_2 = -3; end
		9: begin l_1 = +1;
				 l_2 = +4; end
		6304: begin l_1 = +1;
				 l_2 = -4; end
		7: begin l_1 = -1;
				 l_2 = +4; end
		6302: begin l_1 = -1;
				 l_2 = -4; end
		17: begin l_1 = +1;
				 l_2 = +5; end
		6296: begin l_1 = +1;
				 l_2 = -5; end
		15: begin l_1 = -1;
				 l_2 = +5; end
		6294: begin l_1 = -1;
				 l_2 = -5; end
		33: begin l_1 = +1;
				 l_2 = +6; end
		6280: begin l_1 = +1;
				 l_2 = -6; end
		31: begin l_1 = -1;
				 l_2 = +6; end
		6278: begin l_1 = -1;
				 l_2 = -6; end
		65: begin l_1 = +1;
				 l_2 = +7; end
		6248: begin l_1 = +1;
				 l_2 = -7; end
		63: begin l_1 = -1;
				 l_2 = +7; end
		6246: begin l_1 = -1;
				 l_2 = -7; end
		129: begin l_1 = +1;
				 l_2 = +8; end
		6184: begin l_1 = +1;
				 l_2 = -8; end
		127: begin l_1 = -1;
				 l_2 = +8; end
		6182: begin l_1 = -1;
				 l_2 = -8; end
		257: begin l_1 = +1;
				 l_2 = +9; end
		6056: begin l_1 = +1;
				 l_2 = -9; end
		255: begin l_1 = -1;
				 l_2 = +9; end
		6054: begin l_1 = -1;
				 l_2 = -9; end
		513: begin l_1 = +1;
				 l_2 = +10; end
		5800: begin l_1 = +1;
				 l_2 = -10; end
		511: begin l_1 = -1;
				 l_2 = +10; end
		5798: begin l_1 = -1;
				 l_2 = -10; end
		1025: begin l_1 = +1;
				 l_2 = +11; end
		5288: begin l_1 = +1;
				 l_2 = -11; end
		1023: begin l_1 = -1;
				 l_2 = +11; end
		5286: begin l_1 = -1;
				 l_2 = -11; end
		2049: begin l_1 = +1;
				 l_2 = +12; end
		4264: begin l_1 = +1;
				 l_2 = -12; end
		2047: begin l_1 = -1;
				 l_2 = +12; end
		4262: begin l_1 = -1;
				 l_2 = -12; end
		4097: begin l_1 = +1;
				 l_2 = +13; end
		2216: begin l_1 = +1;
				 l_2 = -13; end
		4095: begin l_1 = -1;
				 l_2 = +13; end
		2214: begin l_1 = -1;
				 l_2 = -13; end
		1882: begin l_1 = +1;
				 l_2 = +14; end
		4431: begin l_1 = +1;
				 l_2 = -14; end
		1880: begin l_1 = -1;
				 l_2 = +14; end
		4429: begin l_1 = -1;
				 l_2 = -14; end
		3763: begin l_1 = +1;
				 l_2 = +15; end
		2550: begin l_1 = +1;
				 l_2 = -15; end
		3761: begin l_1 = -1;
				 l_2 = +15; end
		2548: begin l_1 = -1;
				 l_2 = -15; end
		1214: begin l_1 = +1;
				 l_2 = +16; end
		5099: begin l_1 = +1;
				 l_2 = -16; end
		1212: begin l_1 = -1;
				 l_2 = +16; end
		5097: begin l_1 = -1;
				 l_2 = -16; end
		2427: begin l_1 = +1;
				 l_2 = +17; end
		3886: begin l_1 = +1;
				 l_2 = -17; end
		2425: begin l_1 = -1;
				 l_2 = +17; end
		3884: begin l_1 = -1;
				 l_2 = -17; end
		4853: begin l_1 = +1;
				 l_2 = +18; end
		1460: begin l_1 = +1;
				 l_2 = -18; end
		4851: begin l_1 = -1;
				 l_2 = +18; end
		1458: begin l_1 = -1;
				 l_2 = -18; end
		3394: begin l_1 = +1;
				 l_2 = +19; end
		2919: begin l_1 = +1;
				 l_2 = -19; end
		3392: begin l_1 = -1;
				 l_2 = +19; end
		2917: begin l_1 = -1;
				 l_2 = -19; end
		476: begin l_1 = +1;
				 l_2 = +20; end
		5837: begin l_1 = +1;
				 l_2 = -20; end
		474: begin l_1 = -1;
				 l_2 = +20; end
		5835: begin l_1 = -1;
				 l_2 = -20; end
		951: begin l_1 = +1;
				 l_2 = +21; end
		5362: begin l_1 = +1;
				 l_2 = -21; end
		949: begin l_1 = -1;
				 l_2 = +21; end
		5360: begin l_1 = -1;
				 l_2 = -21; end
		1901: begin l_1 = +1;
				 l_2 = +22; end
		4412: begin l_1 = +1;
				 l_2 = -22; end
		1899: begin l_1 = -1;
				 l_2 = +22; end
		4410: begin l_1 = -1;
				 l_2 = -22; end
		3801: begin l_1 = +1;
				 l_2 = +23; end
		2512: begin l_1 = +1;
				 l_2 = -23; end
		3799: begin l_1 = -1;
				 l_2 = +23; end
		2510: begin l_1 = -1;
				 l_2 = -23; end
		1290: begin l_1 = +1;
				 l_2 = +24; end
		5023: begin l_1 = +1;
				 l_2 = -24; end
		1288: begin l_1 = -1;
				 l_2 = +24; end
		5021: begin l_1 = -1;
				 l_2 = -24; end
		2579: begin l_1 = +1;
				 l_2 = +25; end
		3734: begin l_1 = +1;
				 l_2 = -25; end
		2577: begin l_1 = -1;
				 l_2 = +25; end
		3732: begin l_1 = -1;
				 l_2 = -25; end
		5157: begin l_1 = +1;
				 l_2 = +26; end
		1156: begin l_1 = +1;
				 l_2 = -26; end
		5155: begin l_1 = -1;
				 l_2 = +26; end
		1154: begin l_1 = -1;
				 l_2 = -26; end
		4002: begin l_1 = +1;
				 l_2 = +27; end
		2311: begin l_1 = +1;
				 l_2 = -27; end
		4000: begin l_1 = -1;
				 l_2 = +27; end
		2309: begin l_1 = -1;
				 l_2 = -27; end
		1692: begin l_1 = +1;
				 l_2 = +28; end
		4621: begin l_1 = +1;
				 l_2 = -28; end
		1690: begin l_1 = -1;
				 l_2 = +28; end
		4619: begin l_1 = -1;
				 l_2 = -28; end
		3383: begin l_1 = +1;
				 l_2 = +29; end
		2930: begin l_1 = +1;
				 l_2 = -29; end
		3381: begin l_1 = -1;
				 l_2 = +29; end
		2928: begin l_1 = -1;
				 l_2 = -29; end
		454: begin l_1 = +1;
				 l_2 = +30; end
		5859: begin l_1 = +1;
				 l_2 = -30; end
		452: begin l_1 = -1;
				 l_2 = +30; end
		5857: begin l_1 = -1;
				 l_2 = -30; end
		907: begin l_1 = +1;
				 l_2 = +31; end
		5406: begin l_1 = +1;
				 l_2 = -31; end
		905: begin l_1 = -1;
				 l_2 = +31; end
		5404: begin l_1 = -1;
				 l_2 = -31; end
		1813: begin l_1 = +1;
				 l_2 = +32; end
		4500: begin l_1 = +1;
				 l_2 = -32; end
		1811: begin l_1 = -1;
				 l_2 = +32; end
		4498: begin l_1 = -1;
				 l_2 = -32; end
		3625: begin l_1 = +1;
				 l_2 = +33; end
		2688: begin l_1 = +1;
				 l_2 = -33; end
		3623: begin l_1 = -1;
				 l_2 = +33; end
		2686: begin l_1 = -1;
				 l_2 = -33; end
		6: begin l_1 = -2;
				 l_2 = +4; end
		6305: begin l_1 = -2;
				 l_2 = -3; end
		10: begin l_1 = +2;
				 l_2 = +4; end
		6301: begin l_1 = -2;
				 l_2 = -4; end
		18: begin l_1 = +2;
				 l_2 = +5; end
		6297: begin l_1 = +2;
				 l_2 = -5; end
		14: begin l_1 = -2;
				 l_2 = +5; end
		6293: begin l_1 = -2;
				 l_2 = -5; end
		34: begin l_1 = +2;
				 l_2 = +6; end
		6281: begin l_1 = +2;
				 l_2 = -6; end
		30: begin l_1 = -2;
				 l_2 = +6; end
		6277: begin l_1 = -2;
				 l_2 = -6; end
		66: begin l_1 = +2;
				 l_2 = +7; end
		6249: begin l_1 = +2;
				 l_2 = -7; end
		62: begin l_1 = -2;
				 l_2 = +7; end
		6245: begin l_1 = -2;
				 l_2 = -7; end
		130: begin l_1 = +2;
				 l_2 = +8; end
		6185: begin l_1 = +2;
				 l_2 = -8; end
		126: begin l_1 = -2;
				 l_2 = +8; end
		6181: begin l_1 = -2;
				 l_2 = -8; end
		258: begin l_1 = +2;
				 l_2 = +9; end
		6057: begin l_1 = +2;
				 l_2 = -9; end
		254: begin l_1 = -2;
				 l_2 = +9; end
		6053: begin l_1 = -2;
				 l_2 = -9; end
		514: begin l_1 = +2;
				 l_2 = +10; end
		5801: begin l_1 = +2;
				 l_2 = -10; end
		510: begin l_1 = -2;
				 l_2 = +10; end
		5797: begin l_1 = -2;
				 l_2 = -10; end
		1026: begin l_1 = +2;
				 l_2 = +11; end
		5289: begin l_1 = +2;
				 l_2 = -11; end
		1022: begin l_1 = -2;
				 l_2 = +11; end
		5285: begin l_1 = -2;
				 l_2 = -11; end
		2050: begin l_1 = +2;
				 l_2 = +12; end
		4265: begin l_1 = +2;
				 l_2 = -12; end
		2046: begin l_1 = -2;
				 l_2 = +12; end
		4261: begin l_1 = -2;
				 l_2 = -12; end
		4098: begin l_1 = +2;
				 l_2 = +13; end
		2217: begin l_1 = +2;
				 l_2 = -13; end
		4094: begin l_1 = -2;
				 l_2 = +13; end
		2213: begin l_1 = -2;
				 l_2 = -13; end
		1883: begin l_1 = +2;
				 l_2 = +14; end
		4432: begin l_1 = +2;
				 l_2 = -14; end
		1879: begin l_1 = -2;
				 l_2 = +14; end
		4428: begin l_1 = -2;
				 l_2 = -14; end
		3764: begin l_1 = +2;
				 l_2 = +15; end
		2551: begin l_1 = +2;
				 l_2 = -15; end
		3760: begin l_1 = -2;
				 l_2 = +15; end
		2547: begin l_1 = -2;
				 l_2 = -15; end
		1215: begin l_1 = +2;
				 l_2 = +16; end
		5100: begin l_1 = +2;
				 l_2 = -16; end
		1211: begin l_1 = -2;
				 l_2 = +16; end
		5096: begin l_1 = -2;
				 l_2 = -16; end
		2428: begin l_1 = +2;
				 l_2 = +17; end
		3887: begin l_1 = +2;
				 l_2 = -17; end
		2424: begin l_1 = -2;
				 l_2 = +17; end
		3883: begin l_1 = -2;
				 l_2 = -17; end
		4854: begin l_1 = +2;
				 l_2 = +18; end
		1461: begin l_1 = +2;
				 l_2 = -18; end
		4850: begin l_1 = -2;
				 l_2 = +18; end
		1457: begin l_1 = -2;
				 l_2 = -18; end
		3395: begin l_1 = +2;
				 l_2 = +19; end
		2920: begin l_1 = +2;
				 l_2 = -19; end
		3391: begin l_1 = -2;
				 l_2 = +19; end
		2916: begin l_1 = -2;
				 l_2 = -19; end
		477: begin l_1 = +2;
				 l_2 = +20; end
		5838: begin l_1 = +2;
				 l_2 = -20; end
		473: begin l_1 = -2;
				 l_2 = +20; end
		5834: begin l_1 = -2;
				 l_2 = -20; end
		952: begin l_1 = +2;
				 l_2 = +21; end
		5363: begin l_1 = +2;
				 l_2 = -21; end
		948: begin l_1 = -2;
				 l_2 = +21; end
		5359: begin l_1 = -2;
				 l_2 = -21; end
		1902: begin l_1 = +2;
				 l_2 = +22; end
		4413: begin l_1 = +2;
				 l_2 = -22; end
		1898: begin l_1 = -2;
				 l_2 = +22; end
		4409: begin l_1 = -2;
				 l_2 = -22; end
		3802: begin l_1 = +2;
				 l_2 = +23; end
		2513: begin l_1 = +2;
				 l_2 = -23; end
		3798: begin l_1 = -2;
				 l_2 = +23; end
		2509: begin l_1 = -2;
				 l_2 = -23; end
		1291: begin l_1 = +2;
				 l_2 = +24; end
		5024: begin l_1 = +2;
				 l_2 = -24; end
		1287: begin l_1 = -2;
				 l_2 = +24; end
		5020: begin l_1 = -2;
				 l_2 = -24; end
		2580: begin l_1 = +2;
				 l_2 = +25; end
		3735: begin l_1 = +2;
				 l_2 = -25; end
		2576: begin l_1 = -2;
				 l_2 = +25; end
		3731: begin l_1 = -2;
				 l_2 = -25; end
		5158: begin l_1 = +2;
				 l_2 = +26; end
		1157: begin l_1 = +2;
				 l_2 = -26; end
		5154: begin l_1 = -2;
				 l_2 = +26; end
		1153: begin l_1 = -2;
				 l_2 = -26; end
		4003: begin l_1 = +2;
				 l_2 = +27; end
		2312: begin l_1 = +2;
				 l_2 = -27; end
		3999: begin l_1 = -2;
				 l_2 = +27; end
		2308: begin l_1 = -2;
				 l_2 = -27; end
		1693: begin l_1 = +2;
				 l_2 = +28; end
		4622: begin l_1 = +2;
				 l_2 = -28; end
		1689: begin l_1 = -2;
				 l_2 = +28; end
		4618: begin l_1 = -2;
				 l_2 = -28; end
		3384: begin l_1 = +2;
				 l_2 = +29; end
		2931: begin l_1 = +2;
				 l_2 = -29; end
		3380: begin l_1 = -2;
				 l_2 = +29; end
		2927: begin l_1 = -2;
				 l_2 = -29; end
		455: begin l_1 = +2;
				 l_2 = +30; end
		5860: begin l_1 = +2;
				 l_2 = -30; end
		451: begin l_1 = -2;
				 l_2 = +30; end
		5856: begin l_1 = -2;
				 l_2 = -30; end
		908: begin l_1 = +2;
				 l_2 = +31; end
		5407: begin l_1 = +2;
				 l_2 = -31; end
		904: begin l_1 = -2;
				 l_2 = +31; end
		5403: begin l_1 = -2;
				 l_2 = -31; end
		1814: begin l_1 = +2;
				 l_2 = +32; end
		4501: begin l_1 = +2;
				 l_2 = -32; end
		1810: begin l_1 = -2;
				 l_2 = +32; end
		4497: begin l_1 = -2;
				 l_2 = -32; end
		3626: begin l_1 = +2;
				 l_2 = +33; end
		2689: begin l_1 = +2;
				 l_2 = -33; end
		3622: begin l_1 = -2;
				 l_2 = +33; end
		2685: begin l_1 = -2;
				 l_2 = -33; end
		12: begin l_1 = -3;
				 l_2 = +5; end
		6299: begin l_1 = -3;
				 l_2 = -4; end
		20: begin l_1 = +3;
				 l_2 = +5; end
		6291: begin l_1 = -3;
				 l_2 = -5; end
		36: begin l_1 = +3;
				 l_2 = +6; end
		6283: begin l_1 = +3;
				 l_2 = -6; end
		28: begin l_1 = -3;
				 l_2 = +6; end
		6275: begin l_1 = -3;
				 l_2 = -6; end
		68: begin l_1 = +3;
				 l_2 = +7; end
		6251: begin l_1 = +3;
				 l_2 = -7; end
		60: begin l_1 = -3;
				 l_2 = +7; end
		6243: begin l_1 = -3;
				 l_2 = -7; end
		132: begin l_1 = +3;
				 l_2 = +8; end
		6187: begin l_1 = +3;
				 l_2 = -8; end
		124: begin l_1 = -3;
				 l_2 = +8; end
		6179: begin l_1 = -3;
				 l_2 = -8; end
		260: begin l_1 = +3;
				 l_2 = +9; end
		6059: begin l_1 = +3;
				 l_2 = -9; end
		252: begin l_1 = -3;
				 l_2 = +9; end
		6051: begin l_1 = -3;
				 l_2 = -9; end
		516: begin l_1 = +3;
				 l_2 = +10; end
		5803: begin l_1 = +3;
				 l_2 = -10; end
		508: begin l_1 = -3;
				 l_2 = +10; end
		5795: begin l_1 = -3;
				 l_2 = -10; end
		1028: begin l_1 = +3;
				 l_2 = +11; end
		5291: begin l_1 = +3;
				 l_2 = -11; end
		1020: begin l_1 = -3;
				 l_2 = +11; end
		5283: begin l_1 = -3;
				 l_2 = -11; end
		2052: begin l_1 = +3;
				 l_2 = +12; end
		4267: begin l_1 = +3;
				 l_2 = -12; end
		2044: begin l_1 = -3;
				 l_2 = +12; end
		4259: begin l_1 = -3;
				 l_2 = -12; end
		4100: begin l_1 = +3;
				 l_2 = +13; end
		2219: begin l_1 = +3;
				 l_2 = -13; end
		4092: begin l_1 = -3;
				 l_2 = +13; end
		2211: begin l_1 = -3;
				 l_2 = -13; end
		1885: begin l_1 = +3;
				 l_2 = +14; end
		4434: begin l_1 = +3;
				 l_2 = -14; end
		1877: begin l_1 = -3;
				 l_2 = +14; end
		4426: begin l_1 = -3;
				 l_2 = -14; end
		3766: begin l_1 = +3;
				 l_2 = +15; end
		2553: begin l_1 = +3;
				 l_2 = -15; end
		3758: begin l_1 = -3;
				 l_2 = +15; end
		2545: begin l_1 = -3;
				 l_2 = -15; end
		1217: begin l_1 = +3;
				 l_2 = +16; end
		5102: begin l_1 = +3;
				 l_2 = -16; end
		1209: begin l_1 = -3;
				 l_2 = +16; end
		5094: begin l_1 = -3;
				 l_2 = -16; end
		2430: begin l_1 = +3;
				 l_2 = +17; end
		3889: begin l_1 = +3;
				 l_2 = -17; end
		2422: begin l_1 = -3;
				 l_2 = +17; end
		3881: begin l_1 = -3;
				 l_2 = -17; end
		4856: begin l_1 = +3;
				 l_2 = +18; end
		1463: begin l_1 = +3;
				 l_2 = -18; end
		4848: begin l_1 = -3;
				 l_2 = +18; end
		1455: begin l_1 = -3;
				 l_2 = -18; end
		3397: begin l_1 = +3;
				 l_2 = +19; end
		2922: begin l_1 = +3;
				 l_2 = -19; end
		3389: begin l_1 = -3;
				 l_2 = +19; end
		2914: begin l_1 = -3;
				 l_2 = -19; end
		479: begin l_1 = +3;
				 l_2 = +20; end
		5840: begin l_1 = +3;
				 l_2 = -20; end
		471: begin l_1 = -3;
				 l_2 = +20; end
		5832: begin l_1 = -3;
				 l_2 = -20; end
		954: begin l_1 = +3;
				 l_2 = +21; end
		5365: begin l_1 = +3;
				 l_2 = -21; end
		946: begin l_1 = -3;
				 l_2 = +21; end
		5357: begin l_1 = -3;
				 l_2 = -21; end
		1904: begin l_1 = +3;
				 l_2 = +22; end
		4415: begin l_1 = +3;
				 l_2 = -22; end
		1896: begin l_1 = -3;
				 l_2 = +22; end
		4407: begin l_1 = -3;
				 l_2 = -22; end
		3804: begin l_1 = +3;
				 l_2 = +23; end
		2515: begin l_1 = +3;
				 l_2 = -23; end
		3796: begin l_1 = -3;
				 l_2 = +23; end
		2507: begin l_1 = -3;
				 l_2 = -23; end
		1293: begin l_1 = +3;
				 l_2 = +24; end
		5026: begin l_1 = +3;
				 l_2 = -24; end
		1285: begin l_1 = -3;
				 l_2 = +24; end
		5018: begin l_1 = -3;
				 l_2 = -24; end
		2582: begin l_1 = +3;
				 l_2 = +25; end
		3737: begin l_1 = +3;
				 l_2 = -25; end
		2574: begin l_1 = -3;
				 l_2 = +25; end
		3729: begin l_1 = -3;
				 l_2 = -25; end
		5160: begin l_1 = +3;
				 l_2 = +26; end
		1159: begin l_1 = +3;
				 l_2 = -26; end
		5152: begin l_1 = -3;
				 l_2 = +26; end
		1151: begin l_1 = -3;
				 l_2 = -26; end
		4005: begin l_1 = +3;
				 l_2 = +27; end
		2314: begin l_1 = +3;
				 l_2 = -27; end
		3997: begin l_1 = -3;
				 l_2 = +27; end
		2306: begin l_1 = -3;
				 l_2 = -27; end
		1695: begin l_1 = +3;
				 l_2 = +28; end
		4624: begin l_1 = +3;
				 l_2 = -28; end
		1687: begin l_1 = -3;
				 l_2 = +28; end
		4616: begin l_1 = -3;
				 l_2 = -28; end
		3386: begin l_1 = +3;
				 l_2 = +29; end
		2933: begin l_1 = +3;
				 l_2 = -29; end
		3378: begin l_1 = -3;
				 l_2 = +29; end
		2925: begin l_1 = -3;
				 l_2 = -29; end
		457: begin l_1 = +3;
				 l_2 = +30; end
		5862: begin l_1 = +3;
				 l_2 = -30; end
		449: begin l_1 = -3;
				 l_2 = +30; end
		5854: begin l_1 = -3;
				 l_2 = -30; end
		910: begin l_1 = +3;
				 l_2 = +31; end
		5409: begin l_1 = +3;
				 l_2 = -31; end
		902: begin l_1 = -3;
				 l_2 = +31; end
		5401: begin l_1 = -3;
				 l_2 = -31; end
		1816: begin l_1 = +3;
				 l_2 = +32; end
		4503: begin l_1 = +3;
				 l_2 = -32; end
		1808: begin l_1 = -3;
				 l_2 = +32; end
		4495: begin l_1 = -3;
				 l_2 = -32; end
		3628: begin l_1 = +3;
				 l_2 = +33; end
		2691: begin l_1 = +3;
				 l_2 = -33; end
		3620: begin l_1 = -3;
				 l_2 = +33; end
		2683: begin l_1 = -3;
				 l_2 = -33; end
		24: begin l_1 = -4;
				 l_2 = +6; end
		6287: begin l_1 = -4;
				 l_2 = -5; end
		40: begin l_1 = +4;
				 l_2 = +6; end
		6271: begin l_1 = -4;
				 l_2 = -6; end
		72: begin l_1 = +4;
				 l_2 = +7; end
		6255: begin l_1 = +4;
				 l_2 = -7; end
		56: begin l_1 = -4;
				 l_2 = +7; end
		6239: begin l_1 = -4;
				 l_2 = -7; end
		136: begin l_1 = +4;
				 l_2 = +8; end
		6191: begin l_1 = +4;
				 l_2 = -8; end
		120: begin l_1 = -4;
				 l_2 = +8; end
		6175: begin l_1 = -4;
				 l_2 = -8; end
		264: begin l_1 = +4;
				 l_2 = +9; end
		6063: begin l_1 = +4;
				 l_2 = -9; end
		248: begin l_1 = -4;
				 l_2 = +9; end
		6047: begin l_1 = -4;
				 l_2 = -9; end
		520: begin l_1 = +4;
				 l_2 = +10; end
		5807: begin l_1 = +4;
				 l_2 = -10; end
		504: begin l_1 = -4;
				 l_2 = +10; end
		5791: begin l_1 = -4;
				 l_2 = -10; end
		1032: begin l_1 = +4;
				 l_2 = +11; end
		5295: begin l_1 = +4;
				 l_2 = -11; end
		1016: begin l_1 = -4;
				 l_2 = +11; end
		5279: begin l_1 = -4;
				 l_2 = -11; end
		2056: begin l_1 = +4;
				 l_2 = +12; end
		4271: begin l_1 = +4;
				 l_2 = -12; end
		2040: begin l_1 = -4;
				 l_2 = +12; end
		4255: begin l_1 = -4;
				 l_2 = -12; end
		4104: begin l_1 = +4;
				 l_2 = +13; end
		2223: begin l_1 = +4;
				 l_2 = -13; end
		4088: begin l_1 = -4;
				 l_2 = +13; end
		2207: begin l_1 = -4;
				 l_2 = -13; end
		1889: begin l_1 = +4;
				 l_2 = +14; end
		4438: begin l_1 = +4;
				 l_2 = -14; end
		1873: begin l_1 = -4;
				 l_2 = +14; end
		4422: begin l_1 = -4;
				 l_2 = -14; end
		3770: begin l_1 = +4;
				 l_2 = +15; end
		2557: begin l_1 = +4;
				 l_2 = -15; end
		3754: begin l_1 = -4;
				 l_2 = +15; end
		2541: begin l_1 = -4;
				 l_2 = -15; end
		1221: begin l_1 = +4;
				 l_2 = +16; end
		5106: begin l_1 = +4;
				 l_2 = -16; end
		1205: begin l_1 = -4;
				 l_2 = +16; end
		5090: begin l_1 = -4;
				 l_2 = -16; end
		2434: begin l_1 = +4;
				 l_2 = +17; end
		3893: begin l_1 = +4;
				 l_2 = -17; end
		2418: begin l_1 = -4;
				 l_2 = +17; end
		3877: begin l_1 = -4;
				 l_2 = -17; end
		4860: begin l_1 = +4;
				 l_2 = +18; end
		1467: begin l_1 = +4;
				 l_2 = -18; end
		4844: begin l_1 = -4;
				 l_2 = +18; end
		1451: begin l_1 = -4;
				 l_2 = -18; end
		3401: begin l_1 = +4;
				 l_2 = +19; end
		2926: begin l_1 = +4;
				 l_2 = -19; end
		3385: begin l_1 = -4;
				 l_2 = +19; end
		2910: begin l_1 = -4;
				 l_2 = -19; end
		483: begin l_1 = +4;
				 l_2 = +20; end
		5844: begin l_1 = +4;
				 l_2 = -20; end
		467: begin l_1 = -4;
				 l_2 = +20; end
		5828: begin l_1 = -4;
				 l_2 = -20; end
		958: begin l_1 = +4;
				 l_2 = +21; end
		5369: begin l_1 = +4;
				 l_2 = -21; end
		942: begin l_1 = -4;
				 l_2 = +21; end
		5353: begin l_1 = -4;
				 l_2 = -21; end
		1908: begin l_1 = +4;
				 l_2 = +22; end
		4419: begin l_1 = +4;
				 l_2 = -22; end
		1892: begin l_1 = -4;
				 l_2 = +22; end
		4403: begin l_1 = -4;
				 l_2 = -22; end
		3808: begin l_1 = +4;
				 l_2 = +23; end
		2519: begin l_1 = +4;
				 l_2 = -23; end
		3792: begin l_1 = -4;
				 l_2 = +23; end
		2503: begin l_1 = -4;
				 l_2 = -23; end
		1297: begin l_1 = +4;
				 l_2 = +24; end
		5030: begin l_1 = +4;
				 l_2 = -24; end
		1281: begin l_1 = -4;
				 l_2 = +24; end
		5014: begin l_1 = -4;
				 l_2 = -24; end
		2586: begin l_1 = +4;
				 l_2 = +25; end
		3741: begin l_1 = +4;
				 l_2 = -25; end
		2570: begin l_1 = -4;
				 l_2 = +25; end
		3725: begin l_1 = -4;
				 l_2 = -25; end
		5164: begin l_1 = +4;
				 l_2 = +26; end
		1163: begin l_1 = +4;
				 l_2 = -26; end
		5148: begin l_1 = -4;
				 l_2 = +26; end
		1147: begin l_1 = -4;
				 l_2 = -26; end
		4009: begin l_1 = +4;
				 l_2 = +27; end
		2318: begin l_1 = +4;
				 l_2 = -27; end
		3993: begin l_1 = -4;
				 l_2 = +27; end
		2302: begin l_1 = -4;
				 l_2 = -27; end
		1699: begin l_1 = +4;
				 l_2 = +28; end
		4628: begin l_1 = +4;
				 l_2 = -28; end
		1683: begin l_1 = -4;
				 l_2 = +28; end
		4612: begin l_1 = -4;
				 l_2 = -28; end
		3390: begin l_1 = +4;
				 l_2 = +29; end
		2937: begin l_1 = +4;
				 l_2 = -29; end
		3374: begin l_1 = -4;
				 l_2 = +29; end
		2921: begin l_1 = -4;
				 l_2 = -29; end
		461: begin l_1 = +4;
				 l_2 = +30; end
		5866: begin l_1 = +4;
				 l_2 = -30; end
		445: begin l_1 = -4;
				 l_2 = +30; end
		5850: begin l_1 = -4;
				 l_2 = -30; end
		914: begin l_1 = +4;
				 l_2 = +31; end
		5413: begin l_1 = +4;
				 l_2 = -31; end
		898: begin l_1 = -4;
				 l_2 = +31; end
		5397: begin l_1 = -4;
				 l_2 = -31; end
		1820: begin l_1 = +4;
				 l_2 = +32; end
		4507: begin l_1 = +4;
				 l_2 = -32; end
		1804: begin l_1 = -4;
				 l_2 = +32; end
		4491: begin l_1 = -4;
				 l_2 = -32; end
		3632: begin l_1 = +4;
				 l_2 = +33; end
		2695: begin l_1 = +4;
				 l_2 = -33; end
		3616: begin l_1 = -4;
				 l_2 = +33; end
		2679: begin l_1 = -4;
				 l_2 = -33; end
		48: begin l_1 = -5;
				 l_2 = +7; end
		6263: begin l_1 = -5;
				 l_2 = -6; end
		80: begin l_1 = +5;
				 l_2 = +7; end
		6231: begin l_1 = -5;
				 l_2 = -7; end
		144: begin l_1 = +5;
				 l_2 = +8; end
		6199: begin l_1 = +5;
				 l_2 = -8; end
		112: begin l_1 = -5;
				 l_2 = +8; end
		6167: begin l_1 = -5;
				 l_2 = -8; end
		272: begin l_1 = +5;
				 l_2 = +9; end
		6071: begin l_1 = +5;
				 l_2 = -9; end
		240: begin l_1 = -5;
				 l_2 = +9; end
		6039: begin l_1 = -5;
				 l_2 = -9; end
		528: begin l_1 = +5;
				 l_2 = +10; end
		5815: begin l_1 = +5;
				 l_2 = -10; end
		496: begin l_1 = -5;
				 l_2 = +10; end
		5783: begin l_1 = -5;
				 l_2 = -10; end
		1040: begin l_1 = +5;
				 l_2 = +11; end
		5303: begin l_1 = +5;
				 l_2 = -11; end
		1008: begin l_1 = -5;
				 l_2 = +11; end
		5271: begin l_1 = -5;
				 l_2 = -11; end
		2064: begin l_1 = +5;
				 l_2 = +12; end
		4279: begin l_1 = +5;
				 l_2 = -12; end
		2032: begin l_1 = -5;
				 l_2 = +12; end
		4247: begin l_1 = -5;
				 l_2 = -12; end
		4112: begin l_1 = +5;
				 l_2 = +13; end
		2231: begin l_1 = +5;
				 l_2 = -13; end
		4080: begin l_1 = -5;
				 l_2 = +13; end
		2199: begin l_1 = -5;
				 l_2 = -13; end
		1897: begin l_1 = +5;
				 l_2 = +14; end
		4446: begin l_1 = +5;
				 l_2 = -14; end
		1865: begin l_1 = -5;
				 l_2 = +14; end
		4414: begin l_1 = -5;
				 l_2 = -14; end
		3778: begin l_1 = +5;
				 l_2 = +15; end
		2565: begin l_1 = +5;
				 l_2 = -15; end
		3746: begin l_1 = -5;
				 l_2 = +15; end
		2533: begin l_1 = -5;
				 l_2 = -15; end
		1229: begin l_1 = +5;
				 l_2 = +16; end
		5114: begin l_1 = +5;
				 l_2 = -16; end
		1197: begin l_1 = -5;
				 l_2 = +16; end
		5082: begin l_1 = -5;
				 l_2 = -16; end
		2442: begin l_1 = +5;
				 l_2 = +17; end
		3901: begin l_1 = +5;
				 l_2 = -17; end
		2410: begin l_1 = -5;
				 l_2 = +17; end
		3869: begin l_1 = -5;
				 l_2 = -17; end
		4868: begin l_1 = +5;
				 l_2 = +18; end
		1475: begin l_1 = +5;
				 l_2 = -18; end
		4836: begin l_1 = -5;
				 l_2 = +18; end
		1443: begin l_1 = -5;
				 l_2 = -18; end
		3409: begin l_1 = +5;
				 l_2 = +19; end
		2934: begin l_1 = +5;
				 l_2 = -19; end
		3377: begin l_1 = -5;
				 l_2 = +19; end
		2902: begin l_1 = -5;
				 l_2 = -19; end
		491: begin l_1 = +5;
				 l_2 = +20; end
		5852: begin l_1 = +5;
				 l_2 = -20; end
		459: begin l_1 = -5;
				 l_2 = +20; end
		5820: begin l_1 = -5;
				 l_2 = -20; end
		966: begin l_1 = +5;
				 l_2 = +21; end
		5377: begin l_1 = +5;
				 l_2 = -21; end
		934: begin l_1 = -5;
				 l_2 = +21; end
		5345: begin l_1 = -5;
				 l_2 = -21; end
		1916: begin l_1 = +5;
				 l_2 = +22; end
		4427: begin l_1 = +5;
				 l_2 = -22; end
		1884: begin l_1 = -5;
				 l_2 = +22; end
		4395: begin l_1 = -5;
				 l_2 = -22; end
		3816: begin l_1 = +5;
				 l_2 = +23; end
		2527: begin l_1 = +5;
				 l_2 = -23; end
		3784: begin l_1 = -5;
				 l_2 = +23; end
		2495: begin l_1 = -5;
				 l_2 = -23; end
		1305: begin l_1 = +5;
				 l_2 = +24; end
		5038: begin l_1 = +5;
				 l_2 = -24; end
		1273: begin l_1 = -5;
				 l_2 = +24; end
		5006: begin l_1 = -5;
				 l_2 = -24; end
		2594: begin l_1 = +5;
				 l_2 = +25; end
		3749: begin l_1 = +5;
				 l_2 = -25; end
		2562: begin l_1 = -5;
				 l_2 = +25; end
		3717: begin l_1 = -5;
				 l_2 = -25; end
		5172: begin l_1 = +5;
				 l_2 = +26; end
		1171: begin l_1 = +5;
				 l_2 = -26; end
		5140: begin l_1 = -5;
				 l_2 = +26; end
		1139: begin l_1 = -5;
				 l_2 = -26; end
		4017: begin l_1 = +5;
				 l_2 = +27; end
		2326: begin l_1 = +5;
				 l_2 = -27; end
		3985: begin l_1 = -5;
				 l_2 = +27; end
		2294: begin l_1 = -5;
				 l_2 = -27; end
		1707: begin l_1 = +5;
				 l_2 = +28; end
		4636: begin l_1 = +5;
				 l_2 = -28; end
		1675: begin l_1 = -5;
				 l_2 = +28; end
		4604: begin l_1 = -5;
				 l_2 = -28; end
		3398: begin l_1 = +5;
				 l_2 = +29; end
		2945: begin l_1 = +5;
				 l_2 = -29; end
		3366: begin l_1 = -5;
				 l_2 = +29; end
		2913: begin l_1 = -5;
				 l_2 = -29; end
		469: begin l_1 = +5;
				 l_2 = +30; end
		5874: begin l_1 = +5;
				 l_2 = -30; end
		437: begin l_1 = -5;
				 l_2 = +30; end
		5842: begin l_1 = -5;
				 l_2 = -30; end
		922: begin l_1 = +5;
				 l_2 = +31; end
		5421: begin l_1 = +5;
				 l_2 = -31; end
		890: begin l_1 = -5;
				 l_2 = +31; end
		5389: begin l_1 = -5;
				 l_2 = -31; end
		1828: begin l_1 = +5;
				 l_2 = +32; end
		4515: begin l_1 = +5;
				 l_2 = -32; end
		1796: begin l_1 = -5;
				 l_2 = +32; end
		4483: begin l_1 = -5;
				 l_2 = -32; end
		3640: begin l_1 = +5;
				 l_2 = +33; end
		2703: begin l_1 = +5;
				 l_2 = -33; end
		3608: begin l_1 = -5;
				 l_2 = +33; end
		2671: begin l_1 = -5;
				 l_2 = -33; end
		96: begin l_1 = -6;
				 l_2 = +8; end
		6215: begin l_1 = -6;
				 l_2 = -7; end
		160: begin l_1 = +6;
				 l_2 = +8; end
		6151: begin l_1 = -6;
				 l_2 = -8; end
		288: begin l_1 = +6;
				 l_2 = +9; end
		6087: begin l_1 = +6;
				 l_2 = -9; end
		224: begin l_1 = -6;
				 l_2 = +9; end
		6023: begin l_1 = -6;
				 l_2 = -9; end
		544: begin l_1 = +6;
				 l_2 = +10; end
		5831: begin l_1 = +6;
				 l_2 = -10; end
		480: begin l_1 = -6;
				 l_2 = +10; end
		5767: begin l_1 = -6;
				 l_2 = -10; end
		1056: begin l_1 = +6;
				 l_2 = +11; end
		5319: begin l_1 = +6;
				 l_2 = -11; end
		992: begin l_1 = -6;
				 l_2 = +11; end
		5255: begin l_1 = -6;
				 l_2 = -11; end
		2080: begin l_1 = +6;
				 l_2 = +12; end
		4295: begin l_1 = +6;
				 l_2 = -12; end
		2016: begin l_1 = -6;
				 l_2 = +12; end
		4231: begin l_1 = -6;
				 l_2 = -12; end
		4128: begin l_1 = +6;
				 l_2 = +13; end
		2247: begin l_1 = +6;
				 l_2 = -13; end
		4064: begin l_1 = -6;
				 l_2 = +13; end
		2183: begin l_1 = -6;
				 l_2 = -13; end
		1913: begin l_1 = +6;
				 l_2 = +14; end
		4462: begin l_1 = +6;
				 l_2 = -14; end
		1849: begin l_1 = -6;
				 l_2 = +14; end
		4398: begin l_1 = -6;
				 l_2 = -14; end
		3794: begin l_1 = +6;
				 l_2 = +15; end
		2581: begin l_1 = +6;
				 l_2 = -15; end
		3730: begin l_1 = -6;
				 l_2 = +15; end
		2517: begin l_1 = -6;
				 l_2 = -15; end
		1245: begin l_1 = +6;
				 l_2 = +16; end
		5130: begin l_1 = +6;
				 l_2 = -16; end
		1181: begin l_1 = -6;
				 l_2 = +16; end
		5066: begin l_1 = -6;
				 l_2 = -16; end
		2458: begin l_1 = +6;
				 l_2 = +17; end
		3917: begin l_1 = +6;
				 l_2 = -17; end
		2394: begin l_1 = -6;
				 l_2 = +17; end
		3853: begin l_1 = -6;
				 l_2 = -17; end
		4884: begin l_1 = +6;
				 l_2 = +18; end
		1491: begin l_1 = +6;
				 l_2 = -18; end
		4820: begin l_1 = -6;
				 l_2 = +18; end
		1427: begin l_1 = -6;
				 l_2 = -18; end
		3425: begin l_1 = +6;
				 l_2 = +19; end
		2950: begin l_1 = +6;
				 l_2 = -19; end
		3361: begin l_1 = -6;
				 l_2 = +19; end
		2886: begin l_1 = -6;
				 l_2 = -19; end
		507: begin l_1 = +6;
				 l_2 = +20; end
		5868: begin l_1 = +6;
				 l_2 = -20; end
		443: begin l_1 = -6;
				 l_2 = +20; end
		5804: begin l_1 = -6;
				 l_2 = -20; end
		982: begin l_1 = +6;
				 l_2 = +21; end
		5393: begin l_1 = +6;
				 l_2 = -21; end
		918: begin l_1 = -6;
				 l_2 = +21; end
		5329: begin l_1 = -6;
				 l_2 = -21; end
		1932: begin l_1 = +6;
				 l_2 = +22; end
		4443: begin l_1 = +6;
				 l_2 = -22; end
		1868: begin l_1 = -6;
				 l_2 = +22; end
		4379: begin l_1 = -6;
				 l_2 = -22; end
		3832: begin l_1 = +6;
				 l_2 = +23; end
		2543: begin l_1 = +6;
				 l_2 = -23; end
		3768: begin l_1 = -6;
				 l_2 = +23; end
		2479: begin l_1 = -6;
				 l_2 = -23; end
		1321: begin l_1 = +6;
				 l_2 = +24; end
		5054: begin l_1 = +6;
				 l_2 = -24; end
		1257: begin l_1 = -6;
				 l_2 = +24; end
		4990: begin l_1 = -6;
				 l_2 = -24; end
		2610: begin l_1 = +6;
				 l_2 = +25; end
		3765: begin l_1 = +6;
				 l_2 = -25; end
		2546: begin l_1 = -6;
				 l_2 = +25; end
		3701: begin l_1 = -6;
				 l_2 = -25; end
		5188: begin l_1 = +6;
				 l_2 = +26; end
		1187: begin l_1 = +6;
				 l_2 = -26; end
		5124: begin l_1 = -6;
				 l_2 = +26; end
		1123: begin l_1 = -6;
				 l_2 = -26; end
		4033: begin l_1 = +6;
				 l_2 = +27; end
		2342: begin l_1 = +6;
				 l_2 = -27; end
		3969: begin l_1 = -6;
				 l_2 = +27; end
		2278: begin l_1 = -6;
				 l_2 = -27; end
		1723: begin l_1 = +6;
				 l_2 = +28; end
		4652: begin l_1 = +6;
				 l_2 = -28; end
		1659: begin l_1 = -6;
				 l_2 = +28; end
		4588: begin l_1 = -6;
				 l_2 = -28; end
		3414: begin l_1 = +6;
				 l_2 = +29; end
		2961: begin l_1 = +6;
				 l_2 = -29; end
		3350: begin l_1 = -6;
				 l_2 = +29; end
		2897: begin l_1 = -6;
				 l_2 = -29; end
		485: begin l_1 = +6;
				 l_2 = +30; end
		5890: begin l_1 = +6;
				 l_2 = -30; end
		421: begin l_1 = -6;
				 l_2 = +30; end
		5826: begin l_1 = -6;
				 l_2 = -30; end
		938: begin l_1 = +6;
				 l_2 = +31; end
		5437: begin l_1 = +6;
				 l_2 = -31; end
		874: begin l_1 = -6;
				 l_2 = +31; end
		5373: begin l_1 = -6;
				 l_2 = -31; end
		1844: begin l_1 = +6;
				 l_2 = +32; end
		4531: begin l_1 = +6;
				 l_2 = -32; end
		1780: begin l_1 = -6;
				 l_2 = +32; end
		4467: begin l_1 = -6;
				 l_2 = -32; end
		3656: begin l_1 = +6;
				 l_2 = +33; end
		2719: begin l_1 = +6;
				 l_2 = -33; end
		3592: begin l_1 = -6;
				 l_2 = +33; end
		2655: begin l_1 = -6;
				 l_2 = -33; end
		192: begin l_1 = -7;
				 l_2 = +9; end
		6119: begin l_1 = -7;
				 l_2 = -8; end
		320: begin l_1 = +7;
				 l_2 = +9; end
		5991: begin l_1 = -7;
				 l_2 = -9; end
		576: begin l_1 = +7;
				 l_2 = +10; end
		5863: begin l_1 = +7;
				 l_2 = -10; end
		448: begin l_1 = -7;
				 l_2 = +10; end
		5735: begin l_1 = -7;
				 l_2 = -10; end
		1088: begin l_1 = +7;
				 l_2 = +11; end
		5351: begin l_1 = +7;
				 l_2 = -11; end
		960: begin l_1 = -7;
				 l_2 = +11; end
		5223: begin l_1 = -7;
				 l_2 = -11; end
		2112: begin l_1 = +7;
				 l_2 = +12; end
		4327: begin l_1 = +7;
				 l_2 = -12; end
		1984: begin l_1 = -7;
				 l_2 = +12; end
		4199: begin l_1 = -7;
				 l_2 = -12; end
		4160: begin l_1 = +7;
				 l_2 = +13; end
		2279: begin l_1 = +7;
				 l_2 = -13; end
		4032: begin l_1 = -7;
				 l_2 = +13; end
		2151: begin l_1 = -7;
				 l_2 = -13; end
		1945: begin l_1 = +7;
				 l_2 = +14; end
		4494: begin l_1 = +7;
				 l_2 = -14; end
		1817: begin l_1 = -7;
				 l_2 = +14; end
		4366: begin l_1 = -7;
				 l_2 = -14; end
		3826: begin l_1 = +7;
				 l_2 = +15; end
		2613: begin l_1 = +7;
				 l_2 = -15; end
		3698: begin l_1 = -7;
				 l_2 = +15; end
		2485: begin l_1 = -7;
				 l_2 = -15; end
		1277: begin l_1 = +7;
				 l_2 = +16; end
		5162: begin l_1 = +7;
				 l_2 = -16; end
		1149: begin l_1 = -7;
				 l_2 = +16; end
		5034: begin l_1 = -7;
				 l_2 = -16; end
		2490: begin l_1 = +7;
				 l_2 = +17; end
		3949: begin l_1 = +7;
				 l_2 = -17; end
		2362: begin l_1 = -7;
				 l_2 = +17; end
		3821: begin l_1 = -7;
				 l_2 = -17; end
		4916: begin l_1 = +7;
				 l_2 = +18; end
		1523: begin l_1 = +7;
				 l_2 = -18; end
		4788: begin l_1 = -7;
				 l_2 = +18; end
		1395: begin l_1 = -7;
				 l_2 = -18; end
		3457: begin l_1 = +7;
				 l_2 = +19; end
		2982: begin l_1 = +7;
				 l_2 = -19; end
		3329: begin l_1 = -7;
				 l_2 = +19; end
		2854: begin l_1 = -7;
				 l_2 = -19; end
		539: begin l_1 = +7;
				 l_2 = +20; end
		5900: begin l_1 = +7;
				 l_2 = -20; end
		411: begin l_1 = -7;
				 l_2 = +20; end
		5772: begin l_1 = -7;
				 l_2 = -20; end
		1014: begin l_1 = +7;
				 l_2 = +21; end
		5425: begin l_1 = +7;
				 l_2 = -21; end
		886: begin l_1 = -7;
				 l_2 = +21; end
		5297: begin l_1 = -7;
				 l_2 = -21; end
		1964: begin l_1 = +7;
				 l_2 = +22; end
		4475: begin l_1 = +7;
				 l_2 = -22; end
		1836: begin l_1 = -7;
				 l_2 = +22; end
		4347: begin l_1 = -7;
				 l_2 = -22; end
		3864: begin l_1 = +7;
				 l_2 = +23; end
		2575: begin l_1 = +7;
				 l_2 = -23; end
		3736: begin l_1 = -7;
				 l_2 = +23; end
		2447: begin l_1 = -7;
				 l_2 = -23; end
		1353: begin l_1 = +7;
				 l_2 = +24; end
		5086: begin l_1 = +7;
				 l_2 = -24; end
		1225: begin l_1 = -7;
				 l_2 = +24; end
		4958: begin l_1 = -7;
				 l_2 = -24; end
		2642: begin l_1 = +7;
				 l_2 = +25; end
		3797: begin l_1 = +7;
				 l_2 = -25; end
		2514: begin l_1 = -7;
				 l_2 = +25; end
		3669: begin l_1 = -7;
				 l_2 = -25; end
		5220: begin l_1 = +7;
				 l_2 = +26; end
		1219: begin l_1 = +7;
				 l_2 = -26; end
		5092: begin l_1 = -7;
				 l_2 = +26; end
		1091: begin l_1 = -7;
				 l_2 = -26; end
		4065: begin l_1 = +7;
				 l_2 = +27; end
		2374: begin l_1 = +7;
				 l_2 = -27; end
		3937: begin l_1 = -7;
				 l_2 = +27; end
		2246: begin l_1 = -7;
				 l_2 = -27; end
		1755: begin l_1 = +7;
				 l_2 = +28; end
		4684: begin l_1 = +7;
				 l_2 = -28; end
		1627: begin l_1 = -7;
				 l_2 = +28; end
		4556: begin l_1 = -7;
				 l_2 = -28; end
		3446: begin l_1 = +7;
				 l_2 = +29; end
		2993: begin l_1 = +7;
				 l_2 = -29; end
		3318: begin l_1 = -7;
				 l_2 = +29; end
		2865: begin l_1 = -7;
				 l_2 = -29; end
		517: begin l_1 = +7;
				 l_2 = +30; end
		5922: begin l_1 = +7;
				 l_2 = -30; end
		389: begin l_1 = -7;
				 l_2 = +30; end
		5794: begin l_1 = -7;
				 l_2 = -30; end
		970: begin l_1 = +7;
				 l_2 = +31; end
		5469: begin l_1 = +7;
				 l_2 = -31; end
		842: begin l_1 = -7;
				 l_2 = +31; end
		5341: begin l_1 = -7;
				 l_2 = -31; end
		1876: begin l_1 = +7;
				 l_2 = +32; end
		4563: begin l_1 = +7;
				 l_2 = -32; end
		1748: begin l_1 = -7;
				 l_2 = +32; end
		4435: begin l_1 = -7;
				 l_2 = -32; end
		3688: begin l_1 = +7;
				 l_2 = +33; end
		2751: begin l_1 = +7;
				 l_2 = -33; end
		3560: begin l_1 = -7;
				 l_2 = +33; end
		2623: begin l_1 = -7;
				 l_2 = -33; end
		384: begin l_1 = -8;
				 l_2 = +10; end
		5927: begin l_1 = -8;
				 l_2 = -9; end
		640: begin l_1 = +8;
				 l_2 = +10; end
		5671: begin l_1 = -8;
				 l_2 = -10; end
		1152: begin l_1 = +8;
				 l_2 = +11; end
		5415: begin l_1 = +8;
				 l_2 = -11; end
		896: begin l_1 = -8;
				 l_2 = +11; end
		5159: begin l_1 = -8;
				 l_2 = -11; end
		2176: begin l_1 = +8;
				 l_2 = +12; end
		4391: begin l_1 = +8;
				 l_2 = -12; end
		1920: begin l_1 = -8;
				 l_2 = +12; end
		4135: begin l_1 = -8;
				 l_2 = -12; end
		4224: begin l_1 = +8;
				 l_2 = +13; end
		2343: begin l_1 = +8;
				 l_2 = -13; end
		3968: begin l_1 = -8;
				 l_2 = +13; end
		2087: begin l_1 = -8;
				 l_2 = -13; end
		2009: begin l_1 = +8;
				 l_2 = +14; end
		4558: begin l_1 = +8;
				 l_2 = -14; end
		1753: begin l_1 = -8;
				 l_2 = +14; end
		4302: begin l_1 = -8;
				 l_2 = -14; end
		3890: begin l_1 = +8;
				 l_2 = +15; end
		2677: begin l_1 = +8;
				 l_2 = -15; end
		3634: begin l_1 = -8;
				 l_2 = +15; end
		2421: begin l_1 = -8;
				 l_2 = -15; end
		1341: begin l_1 = +8;
				 l_2 = +16; end
		5226: begin l_1 = +8;
				 l_2 = -16; end
		1085: begin l_1 = -8;
				 l_2 = +16; end
		4970: begin l_1 = -8;
				 l_2 = -16; end
		2554: begin l_1 = +8;
				 l_2 = +17; end
		4013: begin l_1 = +8;
				 l_2 = -17; end
		2298: begin l_1 = -8;
				 l_2 = +17; end
		3757: begin l_1 = -8;
				 l_2 = -17; end
		4980: begin l_1 = +8;
				 l_2 = +18; end
		1587: begin l_1 = +8;
				 l_2 = -18; end
		4724: begin l_1 = -8;
				 l_2 = +18; end
		1331: begin l_1 = -8;
				 l_2 = -18; end
		3521: begin l_1 = +8;
				 l_2 = +19; end
		3046: begin l_1 = +8;
				 l_2 = -19; end
		3265: begin l_1 = -8;
				 l_2 = +19; end
		2790: begin l_1 = -8;
				 l_2 = -19; end
		603: begin l_1 = +8;
				 l_2 = +20; end
		5964: begin l_1 = +8;
				 l_2 = -20; end
		347: begin l_1 = -8;
				 l_2 = +20; end
		5708: begin l_1 = -8;
				 l_2 = -20; end
		1078: begin l_1 = +8;
				 l_2 = +21; end
		5489: begin l_1 = +8;
				 l_2 = -21; end
		822: begin l_1 = -8;
				 l_2 = +21; end
		5233: begin l_1 = -8;
				 l_2 = -21; end
		2028: begin l_1 = +8;
				 l_2 = +22; end
		4539: begin l_1 = +8;
				 l_2 = -22; end
		1772: begin l_1 = -8;
				 l_2 = +22; end
		4283: begin l_1 = -8;
				 l_2 = -22; end
		3928: begin l_1 = +8;
				 l_2 = +23; end
		2639: begin l_1 = +8;
				 l_2 = -23; end
		3672: begin l_1 = -8;
				 l_2 = +23; end
		2383: begin l_1 = -8;
				 l_2 = -23; end
		1417: begin l_1 = +8;
				 l_2 = +24; end
		5150: begin l_1 = +8;
				 l_2 = -24; end
		1161: begin l_1 = -8;
				 l_2 = +24; end
		4894: begin l_1 = -8;
				 l_2 = -24; end
		2706: begin l_1 = +8;
				 l_2 = +25; end
		3861: begin l_1 = +8;
				 l_2 = -25; end
		2450: begin l_1 = -8;
				 l_2 = +25; end
		3605: begin l_1 = -8;
				 l_2 = -25; end
		5284: begin l_1 = +8;
				 l_2 = +26; end
		1283: begin l_1 = +8;
				 l_2 = -26; end
		5028: begin l_1 = -8;
				 l_2 = +26; end
		1027: begin l_1 = -8;
				 l_2 = -26; end
		4129: begin l_1 = +8;
				 l_2 = +27; end
		2438: begin l_1 = +8;
				 l_2 = -27; end
		3873: begin l_1 = -8;
				 l_2 = +27; end
		2182: begin l_1 = -8;
				 l_2 = -27; end
		1819: begin l_1 = +8;
				 l_2 = +28; end
		4748: begin l_1 = +8;
				 l_2 = -28; end
		1563: begin l_1 = -8;
				 l_2 = +28; end
		4492: begin l_1 = -8;
				 l_2 = -28; end
		3510: begin l_1 = +8;
				 l_2 = +29; end
		3057: begin l_1 = +8;
				 l_2 = -29; end
		3254: begin l_1 = -8;
				 l_2 = +29; end
		2801: begin l_1 = -8;
				 l_2 = -29; end
		581: begin l_1 = +8;
				 l_2 = +30; end
		5986: begin l_1 = +8;
				 l_2 = -30; end
		325: begin l_1 = -8;
				 l_2 = +30; end
		5730: begin l_1 = -8;
				 l_2 = -30; end
		1034: begin l_1 = +8;
				 l_2 = +31; end
		5533: begin l_1 = +8;
				 l_2 = -31; end
		778: begin l_1 = -8;
				 l_2 = +31; end
		5277: begin l_1 = -8;
				 l_2 = -31; end
		1940: begin l_1 = +8;
				 l_2 = +32; end
		4627: begin l_1 = +8;
				 l_2 = -32; end
		1684: begin l_1 = -8;
				 l_2 = +32; end
		4371: begin l_1 = -8;
				 l_2 = -32; end
		3752: begin l_1 = +8;
				 l_2 = +33; end
		2815: begin l_1 = +8;
				 l_2 = -33; end
		3496: begin l_1 = -8;
				 l_2 = +33; end
		2559: begin l_1 = -8;
				 l_2 = -33; end
		768: begin l_1 = -9;
				 l_2 = +11; end
		5543: begin l_1 = -9;
				 l_2 = -10; end
		1280: begin l_1 = +9;
				 l_2 = +11; end
		5031: begin l_1 = -9;
				 l_2 = -11; end
		2304: begin l_1 = +9;
				 l_2 = +12; end
		4519: begin l_1 = +9;
				 l_2 = -12; end
		1792: begin l_1 = -9;
				 l_2 = +12; end
		4007: begin l_1 = -9;
				 l_2 = -12; end
		4352: begin l_1 = +9;
				 l_2 = +13; end
		2471: begin l_1 = +9;
				 l_2 = -13; end
		3840: begin l_1 = -9;
				 l_2 = +13; end
		1959: begin l_1 = -9;
				 l_2 = -13; end
		2137: begin l_1 = +9;
				 l_2 = +14; end
		4686: begin l_1 = +9;
				 l_2 = -14; end
		1625: begin l_1 = -9;
				 l_2 = +14; end
		4174: begin l_1 = -9;
				 l_2 = -14; end
		4018: begin l_1 = +9;
				 l_2 = +15; end
		2805: begin l_1 = +9;
				 l_2 = -15; end
		3506: begin l_1 = -9;
				 l_2 = +15; end
		2293: begin l_1 = -9;
				 l_2 = -15; end
		1469: begin l_1 = +9;
				 l_2 = +16; end
		5354: begin l_1 = +9;
				 l_2 = -16; end
		957: begin l_1 = -9;
				 l_2 = +16; end
		4842: begin l_1 = -9;
				 l_2 = -16; end
		2682: begin l_1 = +9;
				 l_2 = +17; end
		4141: begin l_1 = +9;
				 l_2 = -17; end
		2170: begin l_1 = -9;
				 l_2 = +17; end
		3629: begin l_1 = -9;
				 l_2 = -17; end
		5108: begin l_1 = +9;
				 l_2 = +18; end
		1715: begin l_1 = +9;
				 l_2 = -18; end
		4596: begin l_1 = -9;
				 l_2 = +18; end
		1203: begin l_1 = -9;
				 l_2 = -18; end
		3649: begin l_1 = +9;
				 l_2 = +19; end
		3174: begin l_1 = +9;
				 l_2 = -19; end
		3137: begin l_1 = -9;
				 l_2 = +19; end
		2662: begin l_1 = -9;
				 l_2 = -19; end
		731: begin l_1 = +9;
				 l_2 = +20; end
		6092: begin l_1 = +9;
				 l_2 = -20; end
		219: begin l_1 = -9;
				 l_2 = +20; end
		5580: begin l_1 = -9;
				 l_2 = -20; end
		1206: begin l_1 = +9;
				 l_2 = +21; end
		5617: begin l_1 = +9;
				 l_2 = -21; end
		694: begin l_1 = -9;
				 l_2 = +21; end
		5105: begin l_1 = -9;
				 l_2 = -21; end
		2156: begin l_1 = +9;
				 l_2 = +22; end
		4667: begin l_1 = +9;
				 l_2 = -22; end
		1644: begin l_1 = -9;
				 l_2 = +22; end
		4155: begin l_1 = -9;
				 l_2 = -22; end
		4056: begin l_1 = +9;
				 l_2 = +23; end
		2767: begin l_1 = +9;
				 l_2 = -23; end
		3544: begin l_1 = -9;
				 l_2 = +23; end
		2255: begin l_1 = -9;
				 l_2 = -23; end
		1545: begin l_1 = +9;
				 l_2 = +24; end
		5278: begin l_1 = +9;
				 l_2 = -24; end
		1033: begin l_1 = -9;
				 l_2 = +24; end
		4766: begin l_1 = -9;
				 l_2 = -24; end
		2834: begin l_1 = +9;
				 l_2 = +25; end
		3989: begin l_1 = +9;
				 l_2 = -25; end
		2322: begin l_1 = -9;
				 l_2 = +25; end
		3477: begin l_1 = -9;
				 l_2 = -25; end
		5412: begin l_1 = +9;
				 l_2 = +26; end
		1411: begin l_1 = +9;
				 l_2 = -26; end
		4900: begin l_1 = -9;
				 l_2 = +26; end
		899: begin l_1 = -9;
				 l_2 = -26; end
		4257: begin l_1 = +9;
				 l_2 = +27; end
		2566: begin l_1 = +9;
				 l_2 = -27; end
		3745: begin l_1 = -9;
				 l_2 = +27; end
		2054: begin l_1 = -9;
				 l_2 = -27; end
		1947: begin l_1 = +9;
				 l_2 = +28; end
		4876: begin l_1 = +9;
				 l_2 = -28; end
		1435: begin l_1 = -9;
				 l_2 = +28; end
		4364: begin l_1 = -9;
				 l_2 = -28; end
		3638: begin l_1 = +9;
				 l_2 = +29; end
		3185: begin l_1 = +9;
				 l_2 = -29; end
		3126: begin l_1 = -9;
				 l_2 = +29; end
		2673: begin l_1 = -9;
				 l_2 = -29; end
		709: begin l_1 = +9;
				 l_2 = +30; end
		6114: begin l_1 = +9;
				 l_2 = -30; end
		197: begin l_1 = -9;
				 l_2 = +30; end
		5602: begin l_1 = -9;
				 l_2 = -30; end
		1162: begin l_1 = +9;
				 l_2 = +31; end
		5661: begin l_1 = +9;
				 l_2 = -31; end
		650: begin l_1 = -9;
				 l_2 = +31; end
		5149: begin l_1 = -9;
				 l_2 = -31; end
		2068: begin l_1 = +9;
				 l_2 = +32; end
		4755: begin l_1 = +9;
				 l_2 = -32; end
		1556: begin l_1 = -9;
				 l_2 = +32; end
		4243: begin l_1 = -9;
				 l_2 = -32; end
		3880: begin l_1 = +9;
				 l_2 = +33; end
		2943: begin l_1 = +9;
				 l_2 = -33; end
		3368: begin l_1 = -9;
				 l_2 = +33; end
		2431: begin l_1 = -9;
				 l_2 = -33; end
		1536: begin l_1 = -10;
				 l_2 = +12; end
		4775: begin l_1 = -10;
				 l_2 = -11; end
		2560: begin l_1 = +10;
				 l_2 = +12; end
		3751: begin l_1 = -10;
				 l_2 = -12; end
		4608: begin l_1 = +10;
				 l_2 = +13; end
		2727: begin l_1 = +10;
				 l_2 = -13; end
		3584: begin l_1 = -10;
				 l_2 = +13; end
		1703: begin l_1 = -10;
				 l_2 = -13; end
		2393: begin l_1 = +10;
				 l_2 = +14; end
		4942: begin l_1 = +10;
				 l_2 = -14; end
		1369: begin l_1 = -10;
				 l_2 = +14; end
		3918: begin l_1 = -10;
				 l_2 = -14; end
		4274: begin l_1 = +10;
				 l_2 = +15; end
		3061: begin l_1 = +10;
				 l_2 = -15; end
		3250: begin l_1 = -10;
				 l_2 = +15; end
		2037: begin l_1 = -10;
				 l_2 = -15; end
		1725: begin l_1 = +10;
				 l_2 = +16; end
		5610: begin l_1 = +10;
				 l_2 = -16; end
		701: begin l_1 = -10;
				 l_2 = +16; end
		4586: begin l_1 = -10;
				 l_2 = -16; end
		2938: begin l_1 = +10;
				 l_2 = +17; end
		4397: begin l_1 = +10;
				 l_2 = -17; end
		1914: begin l_1 = -10;
				 l_2 = +17; end
		3373: begin l_1 = -10;
				 l_2 = -17; end
		5364: begin l_1 = +10;
				 l_2 = +18; end
		1971: begin l_1 = +10;
				 l_2 = -18; end
		4340: begin l_1 = -10;
				 l_2 = +18; end
		947: begin l_1 = -10;
				 l_2 = -18; end
		3905: begin l_1 = +10;
				 l_2 = +19; end
		3430: begin l_1 = +10;
				 l_2 = -19; end
		2881: begin l_1 = -10;
				 l_2 = +19; end
		2406: begin l_1 = -10;
				 l_2 = -19; end
		987: begin l_1 = +10;
				 l_2 = +20; end
		37: begin l_1 = +10;
				 l_2 = -20; end
		6274: begin l_1 = -10;
				 l_2 = +20; end
		5324: begin l_1 = -10;
				 l_2 = -20; end
		1462: begin l_1 = +10;
				 l_2 = +21; end
		5873: begin l_1 = +10;
				 l_2 = -21; end
		438: begin l_1 = -10;
				 l_2 = +21; end
		4849: begin l_1 = -10;
				 l_2 = -21; end
		2412: begin l_1 = +10;
				 l_2 = +22; end
		4923: begin l_1 = +10;
				 l_2 = -22; end
		1388: begin l_1 = -10;
				 l_2 = +22; end
		3899: begin l_1 = -10;
				 l_2 = -22; end
		4312: begin l_1 = +10;
				 l_2 = +23; end
		3023: begin l_1 = +10;
				 l_2 = -23; end
		3288: begin l_1 = -10;
				 l_2 = +23; end
		1999: begin l_1 = -10;
				 l_2 = -23; end
		1801: begin l_1 = +10;
				 l_2 = +24; end
		5534: begin l_1 = +10;
				 l_2 = -24; end
		777: begin l_1 = -10;
				 l_2 = +24; end
		4510: begin l_1 = -10;
				 l_2 = -24; end
		3090: begin l_1 = +10;
				 l_2 = +25; end
		4245: begin l_1 = +10;
				 l_2 = -25; end
		2066: begin l_1 = -10;
				 l_2 = +25; end
		3221: begin l_1 = -10;
				 l_2 = -25; end
		5668: begin l_1 = +10;
				 l_2 = +26; end
		1667: begin l_1 = +10;
				 l_2 = -26; end
		4644: begin l_1 = -10;
				 l_2 = +26; end
		643: begin l_1 = -10;
				 l_2 = -26; end
		4513: begin l_1 = +10;
				 l_2 = +27; end
		2822: begin l_1 = +10;
				 l_2 = -27; end
		3489: begin l_1 = -10;
				 l_2 = +27; end
		1798: begin l_1 = -10;
				 l_2 = -27; end
		2203: begin l_1 = +10;
				 l_2 = +28; end
		5132: begin l_1 = +10;
				 l_2 = -28; end
		1179: begin l_1 = -10;
				 l_2 = +28; end
		4108: begin l_1 = -10;
				 l_2 = -28; end
		3894: begin l_1 = +10;
				 l_2 = +29; end
		3441: begin l_1 = +10;
				 l_2 = -29; end
		2870: begin l_1 = -10;
				 l_2 = +29; end
		2417: begin l_1 = -10;
				 l_2 = -29; end
		965: begin l_1 = +10;
				 l_2 = +30; end
		59: begin l_1 = +10;
				 l_2 = -30; end
		6252: begin l_1 = -10;
				 l_2 = +30; end
		5346: begin l_1 = -10;
				 l_2 = -30; end
		1418: begin l_1 = +10;
				 l_2 = +31; end
		5917: begin l_1 = +10;
				 l_2 = -31; end
		394: begin l_1 = -10;
				 l_2 = +31; end
		4893: begin l_1 = -10;
				 l_2 = -31; end
		2324: begin l_1 = +10;
				 l_2 = +32; end
		5011: begin l_1 = +10;
				 l_2 = -32; end
		1300: begin l_1 = -10;
				 l_2 = +32; end
		3987: begin l_1 = -10;
				 l_2 = -32; end
		4136: begin l_1 = +10;
				 l_2 = +33; end
		3199: begin l_1 = +10;
				 l_2 = -33; end
		3112: begin l_1 = -10;
				 l_2 = +33; end
		2175: begin l_1 = -10;
				 l_2 = -33; end
		3072: begin l_1 = -11;
				 l_2 = +13; end
		3239: begin l_1 = -11;
				 l_2 = -12; end
		5120: begin l_1 = +11;
				 l_2 = +13; end
		1191: begin l_1 = -11;
				 l_2 = -13; end
		2905: begin l_1 = +11;
				 l_2 = +14; end
		5454: begin l_1 = +11;
				 l_2 = -14; end
		857: begin l_1 = -11;
				 l_2 = +14; end
		3406: begin l_1 = -11;
				 l_2 = -14; end
		4786: begin l_1 = +11;
				 l_2 = +15; end
		3573: begin l_1 = +11;
				 l_2 = -15; end
		2738: begin l_1 = -11;
				 l_2 = +15; end
		1525: begin l_1 = -11;
				 l_2 = -15; end
		2237: begin l_1 = +11;
				 l_2 = +16; end
		6122: begin l_1 = +11;
				 l_2 = -16; end
		189: begin l_1 = -11;
				 l_2 = +16; end
		4074: begin l_1 = -11;
				 l_2 = -16; end
		3450: begin l_1 = +11;
				 l_2 = +17; end
		4909: begin l_1 = +11;
				 l_2 = -17; end
		1402: begin l_1 = -11;
				 l_2 = +17; end
		2861: begin l_1 = -11;
				 l_2 = -17; end
		5876: begin l_1 = +11;
				 l_2 = +18; end
		2483: begin l_1 = +11;
				 l_2 = -18; end
		3828: begin l_1 = -11;
				 l_2 = +18; end
		435: begin l_1 = -11;
				 l_2 = -18; end
		4417: begin l_1 = +11;
				 l_2 = +19; end
		3942: begin l_1 = +11;
				 l_2 = -19; end
		2369: begin l_1 = -11;
				 l_2 = +19; end
		1894: begin l_1 = -11;
				 l_2 = -19; end
		1499: begin l_1 = +11;
				 l_2 = +20; end
		549: begin l_1 = +11;
				 l_2 = -20; end
		5762: begin l_1 = -11;
				 l_2 = +20; end
		4812: begin l_1 = -11;
				 l_2 = -20; end
		1974: begin l_1 = +11;
				 l_2 = +21; end
		74: begin l_1 = +11;
				 l_2 = -21; end
		6237: begin l_1 = -11;
				 l_2 = +21; end
		4337: begin l_1 = -11;
				 l_2 = -21; end
		2924: begin l_1 = +11;
				 l_2 = +22; end
		5435: begin l_1 = +11;
				 l_2 = -22; end
		876: begin l_1 = -11;
				 l_2 = +22; end
		3387: begin l_1 = -11;
				 l_2 = -22; end
		4824: begin l_1 = +11;
				 l_2 = +23; end
		3535: begin l_1 = +11;
				 l_2 = -23; end
		2776: begin l_1 = -11;
				 l_2 = +23; end
		1487: begin l_1 = -11;
				 l_2 = -23; end
		2313: begin l_1 = +11;
				 l_2 = +24; end
		6046: begin l_1 = +11;
				 l_2 = -24; end
		265: begin l_1 = -11;
				 l_2 = +24; end
		3998: begin l_1 = -11;
				 l_2 = -24; end
		3602: begin l_1 = +11;
				 l_2 = +25; end
		4757: begin l_1 = +11;
				 l_2 = -25; end
		1554: begin l_1 = -11;
				 l_2 = +25; end
		2709: begin l_1 = -11;
				 l_2 = -25; end
		6180: begin l_1 = +11;
				 l_2 = +26; end
		2179: begin l_1 = +11;
				 l_2 = -26; end
		4132: begin l_1 = -11;
				 l_2 = +26; end
		131: begin l_1 = -11;
				 l_2 = -26; end
		5025: begin l_1 = +11;
				 l_2 = +27; end
		3334: begin l_1 = +11;
				 l_2 = -27; end
		2977: begin l_1 = -11;
				 l_2 = +27; end
		1286: begin l_1 = -11;
				 l_2 = -27; end
		2715: begin l_1 = +11;
				 l_2 = +28; end
		5644: begin l_1 = +11;
				 l_2 = -28; end
		667: begin l_1 = -11;
				 l_2 = +28; end
		3596: begin l_1 = -11;
				 l_2 = -28; end
		4406: begin l_1 = +11;
				 l_2 = +29; end
		3953: begin l_1 = +11;
				 l_2 = -29; end
		2358: begin l_1 = -11;
				 l_2 = +29; end
		1905: begin l_1 = -11;
				 l_2 = -29; end
		1477: begin l_1 = +11;
				 l_2 = +30; end
		571: begin l_1 = +11;
				 l_2 = -30; end
		5740: begin l_1 = -11;
				 l_2 = +30; end
		4834: begin l_1 = -11;
				 l_2 = -30; end
		1930: begin l_1 = +11;
				 l_2 = +31; end
		118: begin l_1 = +11;
				 l_2 = -31; end
		6193: begin l_1 = -11;
				 l_2 = +31; end
		4381: begin l_1 = -11;
				 l_2 = -31; end
		2836: begin l_1 = +11;
				 l_2 = +32; end
		5523: begin l_1 = +11;
				 l_2 = -32; end
		788: begin l_1 = -11;
				 l_2 = +32; end
		3475: begin l_1 = -11;
				 l_2 = -32; end
		4648: begin l_1 = +11;
				 l_2 = +33; end
		3711: begin l_1 = +11;
				 l_2 = -33; end
		2600: begin l_1 = -11;
				 l_2 = +33; end
		1663: begin l_1 = -11;
				 l_2 = -33; end
		6144: begin l_1 = -12;
				 l_2 = +14; end
		167: begin l_1 = -12;
				 l_2 = -13; end
		3929: begin l_1 = +12;
				 l_2 = +14; end
		2382: begin l_1 = -12;
				 l_2 = -14; end
		5810: begin l_1 = +12;
				 l_2 = +15; end
		4597: begin l_1 = +12;
				 l_2 = -15; end
		1714: begin l_1 = -12;
				 l_2 = +15; end
		501: begin l_1 = -12;
				 l_2 = -15; end
		3261: begin l_1 = +12;
				 l_2 = +16; end
		835: begin l_1 = +12;
				 l_2 = -16; end
		5476: begin l_1 = -12;
				 l_2 = +16; end
		3050: begin l_1 = -12;
				 l_2 = -16; end
		4474: begin l_1 = +12;
				 l_2 = +17; end
		5933: begin l_1 = +12;
				 l_2 = -17; end
		378: begin l_1 = -12;
				 l_2 = +17; end
		1837: begin l_1 = -12;
				 l_2 = -17; end
		589: begin l_1 = +12;
				 l_2 = +18; end
		3507: begin l_1 = +12;
				 l_2 = -18; end
		2804: begin l_1 = -12;
				 l_2 = +18; end
		5722: begin l_1 = -12;
				 l_2 = -18; end
		5441: begin l_1 = +12;
				 l_2 = +19; end
		4966: begin l_1 = +12;
				 l_2 = -19; end
		1345: begin l_1 = -12;
				 l_2 = +19; end
		870: begin l_1 = -12;
				 l_2 = -19; end
		2523: begin l_1 = +12;
				 l_2 = +20; end
		1573: begin l_1 = +12;
				 l_2 = -20; end
		4738: begin l_1 = -12;
				 l_2 = +20; end
		3788: begin l_1 = -12;
				 l_2 = -20; end
		2998: begin l_1 = +12;
				 l_2 = +21; end
		1098: begin l_1 = +12;
				 l_2 = -21; end
		5213: begin l_1 = -12;
				 l_2 = +21; end
		3313: begin l_1 = -12;
				 l_2 = -21; end
		3948: begin l_1 = +12;
				 l_2 = +22; end
		148: begin l_1 = +12;
				 l_2 = -22; end
		6163: begin l_1 = -12;
				 l_2 = +22; end
		2363: begin l_1 = -12;
				 l_2 = -22; end
		5848: begin l_1 = +12;
				 l_2 = +23; end
		4559: begin l_1 = +12;
				 l_2 = -23; end
		1752: begin l_1 = -12;
				 l_2 = +23; end
		463: begin l_1 = -12;
				 l_2 = -23; end
		3337: begin l_1 = +12;
				 l_2 = +24; end
		759: begin l_1 = +12;
				 l_2 = -24; end
		5552: begin l_1 = -12;
				 l_2 = +24; end
		2974: begin l_1 = -12;
				 l_2 = -24; end
		4626: begin l_1 = +12;
				 l_2 = +25; end
		5781: begin l_1 = +12;
				 l_2 = -25; end
		530: begin l_1 = -12;
				 l_2 = +25; end
		1685: begin l_1 = -12;
				 l_2 = -25; end
		893: begin l_1 = +12;
				 l_2 = +26; end
		3203: begin l_1 = +12;
				 l_2 = -26; end
		3108: begin l_1 = -12;
				 l_2 = +26; end
		5418: begin l_1 = -12;
				 l_2 = -26; end
		6049: begin l_1 = +12;
				 l_2 = +27; end
		4358: begin l_1 = +12;
				 l_2 = -27; end
		1953: begin l_1 = -12;
				 l_2 = +27; end
		262: begin l_1 = -12;
				 l_2 = -27; end
		3739: begin l_1 = +12;
				 l_2 = +28; end
		357: begin l_1 = +12;
				 l_2 = -28; end
		5954: begin l_1 = -12;
				 l_2 = +28; end
		2572: begin l_1 = -12;
				 l_2 = -28; end
		5430: begin l_1 = +12;
				 l_2 = +29; end
		4977: begin l_1 = +12;
				 l_2 = -29; end
		1334: begin l_1 = -12;
				 l_2 = +29; end
		881: begin l_1 = -12;
				 l_2 = -29; end
		2501: begin l_1 = +12;
				 l_2 = +30; end
		1595: begin l_1 = +12;
				 l_2 = -30; end
		4716: begin l_1 = -12;
				 l_2 = +30; end
		3810: begin l_1 = -12;
				 l_2 = -30; end
		2954: begin l_1 = +12;
				 l_2 = +31; end
		1142: begin l_1 = +12;
				 l_2 = -31; end
		5169: begin l_1 = -12;
				 l_2 = +31; end
		3357: begin l_1 = -12;
				 l_2 = -31; end
		3860: begin l_1 = +12;
				 l_2 = +32; end
		236: begin l_1 = +12;
				 l_2 = -32; end
		6075: begin l_1 = -12;
				 l_2 = +32; end
		2451: begin l_1 = -12;
				 l_2 = -32; end
		5672: begin l_1 = +12;
				 l_2 = +33; end
		4735: begin l_1 = +12;
				 l_2 = -33; end
		1576: begin l_1 = -12;
				 l_2 = +33; end
		639: begin l_1 = -12;
				 l_2 = -33; end
		5977: begin l_1 = -13;
				 l_2 = +15; end
		334: begin l_1 = -13;
				 l_2 = -14; end
		1547: begin l_1 = +13;
				 l_2 = +15; end
		4764: begin l_1 = -13;
				 l_2 = -15; end
		5309: begin l_1 = +13;
				 l_2 = +16; end
		2883: begin l_1 = +13;
				 l_2 = -16; end
		3428: begin l_1 = -13;
				 l_2 = +16; end
		1002: begin l_1 = -13;
				 l_2 = -16; end
		211: begin l_1 = +13;
				 l_2 = +17; end
		1670: begin l_1 = +13;
				 l_2 = -17; end
		4641: begin l_1 = -13;
				 l_2 = +17; end
		6100: begin l_1 = -13;
				 l_2 = -17; end
		2637: begin l_1 = +13;
				 l_2 = +18; end
		5555: begin l_1 = +13;
				 l_2 = -18; end
		756: begin l_1 = -13;
				 l_2 = +18; end
		3674: begin l_1 = -13;
				 l_2 = -18; end
		1178: begin l_1 = +13;
				 l_2 = +19; end
		703: begin l_1 = +13;
				 l_2 = -19; end
		5608: begin l_1 = -13;
				 l_2 = +19; end
		5133: begin l_1 = -13;
				 l_2 = -19; end
		4571: begin l_1 = +13;
				 l_2 = +20; end
		3621: begin l_1 = +13;
				 l_2 = -20; end
		2690: begin l_1 = -13;
				 l_2 = +20; end
		1740: begin l_1 = -13;
				 l_2 = -20; end
		5046: begin l_1 = +13;
				 l_2 = +21; end
		3146: begin l_1 = +13;
				 l_2 = -21; end
		3165: begin l_1 = -13;
				 l_2 = +21; end
		1265: begin l_1 = -13;
				 l_2 = -21; end
		5996: begin l_1 = +13;
				 l_2 = +22; end
		2196: begin l_1 = +13;
				 l_2 = -22; end
		4115: begin l_1 = -13;
				 l_2 = +22; end
		315: begin l_1 = -13;
				 l_2 = -22; end
		1585: begin l_1 = +13;
				 l_2 = +23; end
		296: begin l_1 = +13;
				 l_2 = -23; end
		6015: begin l_1 = -13;
				 l_2 = +23; end
		4726: begin l_1 = -13;
				 l_2 = -23; end
		5385: begin l_1 = +13;
				 l_2 = +24; end
		2807: begin l_1 = +13;
				 l_2 = -24; end
		3504: begin l_1 = -13;
				 l_2 = +24; end
		926: begin l_1 = -13;
				 l_2 = -24; end
		363: begin l_1 = +13;
				 l_2 = +25; end
		1518: begin l_1 = +13;
				 l_2 = -25; end
		4793: begin l_1 = -13;
				 l_2 = +25; end
		5948: begin l_1 = -13;
				 l_2 = -25; end
		2941: begin l_1 = +13;
				 l_2 = +26; end
		5251: begin l_1 = +13;
				 l_2 = -26; end
		1060: begin l_1 = -13;
				 l_2 = +26; end
		3370: begin l_1 = -13;
				 l_2 = -26; end
		1786: begin l_1 = +13;
				 l_2 = +27; end
		95: begin l_1 = +13;
				 l_2 = -27; end
		6216: begin l_1 = -13;
				 l_2 = +27; end
		4525: begin l_1 = -13;
				 l_2 = -27; end
		5787: begin l_1 = +13;
				 l_2 = +28; end
		2405: begin l_1 = +13;
				 l_2 = -28; end
		3906: begin l_1 = -13;
				 l_2 = +28; end
		524: begin l_1 = -13;
				 l_2 = -28; end
		1167: begin l_1 = +13;
				 l_2 = +29; end
		714: begin l_1 = +13;
				 l_2 = -29; end
		5597: begin l_1 = -13;
				 l_2 = +29; end
		5144: begin l_1 = -13;
				 l_2 = -29; end
		4549: begin l_1 = +13;
				 l_2 = +30; end
		3643: begin l_1 = +13;
				 l_2 = -30; end
		2668: begin l_1 = -13;
				 l_2 = +30; end
		1762: begin l_1 = -13;
				 l_2 = -30; end
		5002: begin l_1 = +13;
				 l_2 = +31; end
		3190: begin l_1 = +13;
				 l_2 = -31; end
		3121: begin l_1 = -13;
				 l_2 = +31; end
		1309: begin l_1 = -13;
				 l_2 = -31; end
		5908: begin l_1 = +13;
				 l_2 = +32; end
		2284: begin l_1 = +13;
				 l_2 = -32; end
		4027: begin l_1 = -13;
				 l_2 = +32; end
		403: begin l_1 = -13;
				 l_2 = -32; end
		1409: begin l_1 = +13;
				 l_2 = +33; end
		472: begin l_1 = +13;
				 l_2 = -33; end
		5839: begin l_1 = -13;
				 l_2 = +33; end
		4902: begin l_1 = -13;
				 l_2 = -33; end
		5643: begin l_1 = -14;
				 l_2 = +16; end
		668: begin l_1 = -14;
				 l_2 = -15; end
		3094: begin l_1 = +14;
				 l_2 = +16; end
		3217: begin l_1 = -14;
				 l_2 = -16; end
		4307: begin l_1 = +14;
				 l_2 = +17; end
		5766: begin l_1 = +14;
				 l_2 = -17; end
		545: begin l_1 = -14;
				 l_2 = +17; end
		2004: begin l_1 = -14;
				 l_2 = -17; end
		422: begin l_1 = +14;
				 l_2 = +18; end
		3340: begin l_1 = +14;
				 l_2 = -18; end
		2971: begin l_1 = -14;
				 l_2 = +18; end
		5889: begin l_1 = -14;
				 l_2 = -18; end
		5274: begin l_1 = +14;
				 l_2 = +19; end
		4799: begin l_1 = +14;
				 l_2 = -19; end
		1512: begin l_1 = -14;
				 l_2 = +19; end
		1037: begin l_1 = -14;
				 l_2 = -19; end
		2356: begin l_1 = +14;
				 l_2 = +20; end
		1406: begin l_1 = +14;
				 l_2 = -20; end
		4905: begin l_1 = -14;
				 l_2 = +20; end
		3955: begin l_1 = -14;
				 l_2 = -20; end
		2831: begin l_1 = +14;
				 l_2 = +21; end
		931: begin l_1 = +14;
				 l_2 = -21; end
		5380: begin l_1 = -14;
				 l_2 = +21; end
		3480: begin l_1 = -14;
				 l_2 = -21; end
		3781: begin l_1 = +14;
				 l_2 = +22; end
		6292: begin l_1 = +14;
				 l_2 = -22; end
		19: begin l_1 = -14;
				 l_2 = +22; end
		2530: begin l_1 = -14;
				 l_2 = -22; end
		5681: begin l_1 = +14;
				 l_2 = +23; end
		4392: begin l_1 = +14;
				 l_2 = -23; end
		1919: begin l_1 = -14;
				 l_2 = +23; end
		630: begin l_1 = -14;
				 l_2 = -23; end
		3170: begin l_1 = +14;
				 l_2 = +24; end
		592: begin l_1 = +14;
				 l_2 = -24; end
		5719: begin l_1 = -14;
				 l_2 = +24; end
		3141: begin l_1 = -14;
				 l_2 = -24; end
		4459: begin l_1 = +14;
				 l_2 = +25; end
		5614: begin l_1 = +14;
				 l_2 = -25; end
		697: begin l_1 = -14;
				 l_2 = +25; end
		1852: begin l_1 = -14;
				 l_2 = -25; end
		726: begin l_1 = +14;
				 l_2 = +26; end
		3036: begin l_1 = +14;
				 l_2 = -26; end
		3275: begin l_1 = -14;
				 l_2 = +26; end
		5585: begin l_1 = -14;
				 l_2 = -26; end
		5882: begin l_1 = +14;
				 l_2 = +27; end
		4191: begin l_1 = +14;
				 l_2 = -27; end
		2120: begin l_1 = -14;
				 l_2 = +27; end
		429: begin l_1 = -14;
				 l_2 = -27; end
		3572: begin l_1 = +14;
				 l_2 = +28; end
		190: begin l_1 = +14;
				 l_2 = -28; end
		6121: begin l_1 = -14;
				 l_2 = +28; end
		2739: begin l_1 = -14;
				 l_2 = -28; end
		5263: begin l_1 = +14;
				 l_2 = +29; end
		4810: begin l_1 = +14;
				 l_2 = -29; end
		1501: begin l_1 = -14;
				 l_2 = +29; end
		1048: begin l_1 = -14;
				 l_2 = -29; end
		2334: begin l_1 = +14;
				 l_2 = +30; end
		1428: begin l_1 = +14;
				 l_2 = -30; end
		4883: begin l_1 = -14;
				 l_2 = +30; end
		3977: begin l_1 = -14;
				 l_2 = -30; end
		2787: begin l_1 = +14;
				 l_2 = +31; end
		975: begin l_1 = +14;
				 l_2 = -31; end
		5336: begin l_1 = -14;
				 l_2 = +31; end
		3524: begin l_1 = -14;
				 l_2 = -31; end
		3693: begin l_1 = +14;
				 l_2 = +32; end
		69: begin l_1 = +14;
				 l_2 = -32; end
		6242: begin l_1 = -14;
				 l_2 = +32; end
		2618: begin l_1 = -14;
				 l_2 = -32; end
		5505: begin l_1 = +14;
				 l_2 = +33; end
		4568: begin l_1 = +14;
				 l_2 = -33; end
		1743: begin l_1 = -14;
				 l_2 = +33; end
		806: begin l_1 = -14;
				 l_2 = -33; end
		4975: begin l_1 = -15;
				 l_2 = +17; end
		1336: begin l_1 = -15;
				 l_2 = -16; end
		6188: begin l_1 = +15;
				 l_2 = +17; end
		123: begin l_1 = -15;
				 l_2 = -17; end
		2303: begin l_1 = +15;
				 l_2 = +18; end
		5221: begin l_1 = +15;
				 l_2 = -18; end
		1090: begin l_1 = -15;
				 l_2 = +18; end
		4008: begin l_1 = -15;
				 l_2 = -18; end
		844: begin l_1 = +15;
				 l_2 = +19; end
		369: begin l_1 = +15;
				 l_2 = -19; end
		5942: begin l_1 = -15;
				 l_2 = +19; end
		5467: begin l_1 = -15;
				 l_2 = -19; end
		4237: begin l_1 = +15;
				 l_2 = +20; end
		3287: begin l_1 = +15;
				 l_2 = -20; end
		3024: begin l_1 = -15;
				 l_2 = +20; end
		2074: begin l_1 = -15;
				 l_2 = -20; end
		4712: begin l_1 = +15;
				 l_2 = +21; end
		2812: begin l_1 = +15;
				 l_2 = -21; end
		3499: begin l_1 = -15;
				 l_2 = +21; end
		1599: begin l_1 = -15;
				 l_2 = -21; end
		5662: begin l_1 = +15;
				 l_2 = +22; end
		1862: begin l_1 = +15;
				 l_2 = -22; end
		4449: begin l_1 = -15;
				 l_2 = +22; end
		649: begin l_1 = -15;
				 l_2 = -22; end
		1251: begin l_1 = +15;
				 l_2 = +23; end
		6273: begin l_1 = +15;
				 l_2 = -23; end
		38: begin l_1 = -15;
				 l_2 = +23; end
		5060: begin l_1 = -15;
				 l_2 = -23; end
		5051: begin l_1 = +15;
				 l_2 = +24; end
		2473: begin l_1 = +15;
				 l_2 = -24; end
		3838: begin l_1 = -15;
				 l_2 = +24; end
		1260: begin l_1 = -15;
				 l_2 = -24; end
		29: begin l_1 = +15;
				 l_2 = +25; end
		1184: begin l_1 = +15;
				 l_2 = -25; end
		5127: begin l_1 = -15;
				 l_2 = +25; end
		6282: begin l_1 = -15;
				 l_2 = -25; end
		2607: begin l_1 = +15;
				 l_2 = +26; end
		4917: begin l_1 = +15;
				 l_2 = -26; end
		1394: begin l_1 = -15;
				 l_2 = +26; end
		3704: begin l_1 = -15;
				 l_2 = -26; end
		1452: begin l_1 = +15;
				 l_2 = +27; end
		6072: begin l_1 = +15;
				 l_2 = -27; end
		239: begin l_1 = -15;
				 l_2 = +27; end
		4859: begin l_1 = -15;
				 l_2 = -27; end
		5453: begin l_1 = +15;
				 l_2 = +28; end
		2071: begin l_1 = +15;
				 l_2 = -28; end
		4240: begin l_1 = -15;
				 l_2 = +28; end
		858: begin l_1 = -15;
				 l_2 = -28; end
		833: begin l_1 = +15;
				 l_2 = +29; end
		380: begin l_1 = +15;
				 l_2 = -29; end
		5931: begin l_1 = -15;
				 l_2 = +29; end
		5478: begin l_1 = -15;
				 l_2 = -29; end
		4215: begin l_1 = +15;
				 l_2 = +30; end
		3309: begin l_1 = +15;
				 l_2 = -30; end
		3002: begin l_1 = -15;
				 l_2 = +30; end
		2096: begin l_1 = -15;
				 l_2 = -30; end
		4668: begin l_1 = +15;
				 l_2 = +31; end
		2856: begin l_1 = +15;
				 l_2 = -31; end
		3455: begin l_1 = -15;
				 l_2 = +31; end
		1643: begin l_1 = -15;
				 l_2 = -31; end
		5574: begin l_1 = +15;
				 l_2 = +32; end
		1950: begin l_1 = +15;
				 l_2 = -32; end
		4361: begin l_1 = -15;
				 l_2 = +32; end
		737: begin l_1 = -15;
				 l_2 = -32; end
		1075: begin l_1 = +15;
				 l_2 = +33; end
		138: begin l_1 = +15;
				 l_2 = -33; end
		6173: begin l_1 = -15;
				 l_2 = +33; end
		5236: begin l_1 = -15;
				 l_2 = -33; end
		3639: begin l_1 = -16;
				 l_2 = +18; end
		2672: begin l_1 = -16;
				 l_2 = -17; end
		6065: begin l_1 = +16;
				 l_2 = +18; end
		246: begin l_1 = -16;
				 l_2 = -18; end
		4606: begin l_1 = +16;
				 l_2 = +19; end
		4131: begin l_1 = +16;
				 l_2 = -19; end
		2180: begin l_1 = -16;
				 l_2 = +19; end
		1705: begin l_1 = -16;
				 l_2 = -19; end
		1688: begin l_1 = +16;
				 l_2 = +20; end
		738: begin l_1 = +16;
				 l_2 = -20; end
		5573: begin l_1 = -16;
				 l_2 = +20; end
		4623: begin l_1 = -16;
				 l_2 = -20; end
		2163: begin l_1 = +16;
				 l_2 = +21; end
		263: begin l_1 = +16;
				 l_2 = -21; end
		6048: begin l_1 = -16;
				 l_2 = +21; end
		4148: begin l_1 = -16;
				 l_2 = -21; end
		3113: begin l_1 = +16;
				 l_2 = +22; end
		5624: begin l_1 = +16;
				 l_2 = -22; end
		687: begin l_1 = -16;
				 l_2 = +22; end
		3198: begin l_1 = -16;
				 l_2 = -22; end
		5013: begin l_1 = +16;
				 l_2 = +23; end
		3724: begin l_1 = +16;
				 l_2 = -23; end
		2587: begin l_1 = -16;
				 l_2 = +23; end
		1298: begin l_1 = -16;
				 l_2 = -23; end
		2502: begin l_1 = +16;
				 l_2 = +24; end
		6235: begin l_1 = +16;
				 l_2 = -24; end
		76: begin l_1 = -16;
				 l_2 = +24; end
		3809: begin l_1 = -16;
				 l_2 = -24; end
		3791: begin l_1 = +16;
				 l_2 = +25; end
		4946: begin l_1 = +16;
				 l_2 = -25; end
		1365: begin l_1 = -16;
				 l_2 = +25; end
		2520: begin l_1 = -16;
				 l_2 = -25; end
		58: begin l_1 = +16;
				 l_2 = +26; end
		2368: begin l_1 = +16;
				 l_2 = -26; end
		3943: begin l_1 = -16;
				 l_2 = +26; end
		6253: begin l_1 = -16;
				 l_2 = -26; end
		5214: begin l_1 = +16;
				 l_2 = +27; end
		3523: begin l_1 = +16;
				 l_2 = -27; end
		2788: begin l_1 = -16;
				 l_2 = +27; end
		1097: begin l_1 = -16;
				 l_2 = -27; end
		2904: begin l_1 = +16;
				 l_2 = +28; end
		5833: begin l_1 = +16;
				 l_2 = -28; end
		478: begin l_1 = -16;
				 l_2 = +28; end
		3407: begin l_1 = -16;
				 l_2 = -28; end
		4595: begin l_1 = +16;
				 l_2 = +29; end
		4142: begin l_1 = +16;
				 l_2 = -29; end
		2169: begin l_1 = -16;
				 l_2 = +29; end
		1716: begin l_1 = -16;
				 l_2 = -29; end
		1666: begin l_1 = +16;
				 l_2 = +30; end
		760: begin l_1 = +16;
				 l_2 = -30; end
		5551: begin l_1 = -16;
				 l_2 = +30; end
		4645: begin l_1 = -16;
				 l_2 = -30; end
		2119: begin l_1 = +16;
				 l_2 = +31; end
		307: begin l_1 = +16;
				 l_2 = -31; end
		6004: begin l_1 = -16;
				 l_2 = +31; end
		4192: begin l_1 = -16;
				 l_2 = -31; end
		3025: begin l_1 = +16;
				 l_2 = +32; end
		5712: begin l_1 = +16;
				 l_2 = -32; end
		599: begin l_1 = -16;
				 l_2 = +32; end
		3286: begin l_1 = -16;
				 l_2 = -32; end
		4837: begin l_1 = +16;
				 l_2 = +33; end
		3900: begin l_1 = +16;
				 l_2 = -33; end
		2411: begin l_1 = -16;
				 l_2 = +33; end
		1474: begin l_1 = -16;
				 l_2 = -33; end
		967: begin l_1 = -17;
				 l_2 = +19; end
		5344: begin l_1 = -17;
				 l_2 = -18; end
		5819: begin l_1 = +17;
				 l_2 = +19; end
		492: begin l_1 = -17;
				 l_2 = -19; end
		2901: begin l_1 = +17;
				 l_2 = +20; end
		1951: begin l_1 = +17;
				 l_2 = -20; end
		4360: begin l_1 = -17;
				 l_2 = +20; end
		3410: begin l_1 = -17;
				 l_2 = -20; end
		3376: begin l_1 = +17;
				 l_2 = +21; end
		1476: begin l_1 = +17;
				 l_2 = -21; end
		4835: begin l_1 = -17;
				 l_2 = +21; end
		2935: begin l_1 = -17;
				 l_2 = -21; end
		4326: begin l_1 = +17;
				 l_2 = +22; end
		526: begin l_1 = +17;
				 l_2 = -22; end
		5785: begin l_1 = -17;
				 l_2 = +22; end
		1985: begin l_1 = -17;
				 l_2 = -22; end
		6226: begin l_1 = +17;
				 l_2 = +23; end
		4937: begin l_1 = +17;
				 l_2 = -23; end
		1374: begin l_1 = -17;
				 l_2 = +23; end
		85: begin l_1 = -17;
				 l_2 = -23; end
		3715: begin l_1 = +17;
				 l_2 = +24; end
		1137: begin l_1 = +17;
				 l_2 = -24; end
		5174: begin l_1 = -17;
				 l_2 = +24; end
		2596: begin l_1 = -17;
				 l_2 = -24; end
		5004: begin l_1 = +17;
				 l_2 = +25; end
		6159: begin l_1 = +17;
				 l_2 = -25; end
		152: begin l_1 = -17;
				 l_2 = +25; end
		1307: begin l_1 = -17;
				 l_2 = -25; end
		1271: begin l_1 = +17;
				 l_2 = +26; end
		3581: begin l_1 = +17;
				 l_2 = -26; end
		2730: begin l_1 = -17;
				 l_2 = +26; end
		5040: begin l_1 = -17;
				 l_2 = -26; end
		116: begin l_1 = +17;
				 l_2 = +27; end
		4736: begin l_1 = +17;
				 l_2 = -27; end
		1575: begin l_1 = -17;
				 l_2 = +27; end
		6195: begin l_1 = -17;
				 l_2 = -27; end
		4117: begin l_1 = +17;
				 l_2 = +28; end
		735: begin l_1 = +17;
				 l_2 = -28; end
		5576: begin l_1 = -17;
				 l_2 = +28; end
		2194: begin l_1 = -17;
				 l_2 = -28; end
		5808: begin l_1 = +17;
				 l_2 = +29; end
		5355: begin l_1 = +17;
				 l_2 = -29; end
		956: begin l_1 = -17;
				 l_2 = +29; end
		503: begin l_1 = -17;
				 l_2 = -29; end
		2879: begin l_1 = +17;
				 l_2 = +30; end
		1973: begin l_1 = +17;
				 l_2 = -30; end
		4338: begin l_1 = -17;
				 l_2 = +30; end
		3432: begin l_1 = -17;
				 l_2 = -30; end
		3332: begin l_1 = +17;
				 l_2 = +31; end
		1520: begin l_1 = +17;
				 l_2 = -31; end
		4791: begin l_1 = -17;
				 l_2 = +31; end
		2979: begin l_1 = -17;
				 l_2 = -31; end
		4238: begin l_1 = +17;
				 l_2 = +32; end
		614: begin l_1 = +17;
				 l_2 = -32; end
		5697: begin l_1 = -17;
				 l_2 = +32; end
		2073: begin l_1 = -17;
				 l_2 = -32; end
		6050: begin l_1 = +17;
				 l_2 = +33; end
		5113: begin l_1 = +17;
				 l_2 = -33; end
		1198: begin l_1 = -17;
				 l_2 = +33; end
		261: begin l_1 = -17;
				 l_2 = -33; end
		1934: begin l_1 = -18;
				 l_2 = +20; end
		4377: begin l_1 = -18;
				 l_2 = -19; end
		5327: begin l_1 = +18;
				 l_2 = +20; end
		984: begin l_1 = -18;
				 l_2 = -20; end
		5802: begin l_1 = +18;
				 l_2 = +21; end
		3902: begin l_1 = +18;
				 l_2 = -21; end
		2409: begin l_1 = -18;
				 l_2 = +21; end
		509: begin l_1 = -18;
				 l_2 = -21; end
		441: begin l_1 = +18;
				 l_2 = +22; end
		2952: begin l_1 = +18;
				 l_2 = -22; end
		3359: begin l_1 = -18;
				 l_2 = +22; end
		5870: begin l_1 = -18;
				 l_2 = -22; end
		2341: begin l_1 = +18;
				 l_2 = +23; end
		1052: begin l_1 = +18;
				 l_2 = -23; end
		5259: begin l_1 = -18;
				 l_2 = +23; end
		3970: begin l_1 = -18;
				 l_2 = -23; end
		6141: begin l_1 = +18;
				 l_2 = +24; end
		3563: begin l_1 = +18;
				 l_2 = -24; end
		2748: begin l_1 = -18;
				 l_2 = +24; end
		170: begin l_1 = -18;
				 l_2 = -24; end
		1119: begin l_1 = +18;
				 l_2 = +25; end
		2274: begin l_1 = +18;
				 l_2 = -25; end
		4037: begin l_1 = -18;
				 l_2 = +25; end
		5192: begin l_1 = -18;
				 l_2 = -25; end
		3697: begin l_1 = +18;
				 l_2 = +26; end
		6007: begin l_1 = +18;
				 l_2 = -26; end
		304: begin l_1 = -18;
				 l_2 = +26; end
		2614: begin l_1 = -18;
				 l_2 = -26; end
		2542: begin l_1 = +18;
				 l_2 = +27; end
		851: begin l_1 = +18;
				 l_2 = -27; end
		5460: begin l_1 = -18;
				 l_2 = +27; end
		3769: begin l_1 = -18;
				 l_2 = -27; end
		232: begin l_1 = +18;
				 l_2 = +28; end
		3161: begin l_1 = +18;
				 l_2 = -28; end
		3150: begin l_1 = -18;
				 l_2 = +28; end
		6079: begin l_1 = -18;
				 l_2 = -28; end
		1923: begin l_1 = +18;
				 l_2 = +29; end
		1470: begin l_1 = +18;
				 l_2 = -29; end
		4841: begin l_1 = -18;
				 l_2 = +29; end
		4388: begin l_1 = -18;
				 l_2 = -29; end
		5305: begin l_1 = +18;
				 l_2 = +30; end
		4399: begin l_1 = +18;
				 l_2 = -30; end
		1912: begin l_1 = -18;
				 l_2 = +30; end
		1006: begin l_1 = -18;
				 l_2 = -30; end
		5758: begin l_1 = +18;
				 l_2 = +31; end
		3946: begin l_1 = +18;
				 l_2 = -31; end
		2365: begin l_1 = -18;
				 l_2 = +31; end
		553: begin l_1 = -18;
				 l_2 = -31; end
		353: begin l_1 = +18;
				 l_2 = +32; end
		3040: begin l_1 = +18;
				 l_2 = -32; end
		3271: begin l_1 = -18;
				 l_2 = +32; end
		5958: begin l_1 = -18;
				 l_2 = -32; end
		2165: begin l_1 = +18;
				 l_2 = +33; end
		1228: begin l_1 = +18;
				 l_2 = -33; end
		5083: begin l_1 = -18;
				 l_2 = +33; end
		4146: begin l_1 = -18;
				 l_2 = -33; end
		3868: begin l_1 = -19;
				 l_2 = +21; end
		2443: begin l_1 = -19;
				 l_2 = -20; end
		4343: begin l_1 = +19;
				 l_2 = +21; end
		1968: begin l_1 = -19;
				 l_2 = -21; end
		5293: begin l_1 = +19;
				 l_2 = +22; end
		1493: begin l_1 = +19;
				 l_2 = -22; end
		4818: begin l_1 = -19;
				 l_2 = +22; end
		1018: begin l_1 = -19;
				 l_2 = -22; end
		882: begin l_1 = +19;
				 l_2 = +23; end
		5904: begin l_1 = +19;
				 l_2 = -23; end
		407: begin l_1 = -19;
				 l_2 = +23; end
		5429: begin l_1 = -19;
				 l_2 = -23; end
		4682: begin l_1 = +19;
				 l_2 = +24; end
		2104: begin l_1 = +19;
				 l_2 = -24; end
		4207: begin l_1 = -19;
				 l_2 = +24; end
		1629: begin l_1 = -19;
				 l_2 = -24; end
		5971: begin l_1 = +19;
				 l_2 = +25; end
		815: begin l_1 = +19;
				 l_2 = -25; end
		5496: begin l_1 = -19;
				 l_2 = +25; end
		340: begin l_1 = -19;
				 l_2 = -25; end
		2238: begin l_1 = +19;
				 l_2 = +26; end
		4548: begin l_1 = +19;
				 l_2 = -26; end
		1763: begin l_1 = -19;
				 l_2 = +26; end
		4073: begin l_1 = -19;
				 l_2 = -26; end
		1083: begin l_1 = +19;
				 l_2 = +27; end
		5703: begin l_1 = +19;
				 l_2 = -27; end
		608: begin l_1 = -19;
				 l_2 = +27; end
		5228: begin l_1 = -19;
				 l_2 = -27; end
		5084: begin l_1 = +19;
				 l_2 = +28; end
		1702: begin l_1 = +19;
				 l_2 = -28; end
		4609: begin l_1 = -19;
				 l_2 = +28; end
		1227: begin l_1 = -19;
				 l_2 = -28; end
		464: begin l_1 = +19;
				 l_2 = +29; end
		11: begin l_1 = +19;
				 l_2 = -29; end
		6300: begin l_1 = -19;
				 l_2 = +29; end
		5847: begin l_1 = -19;
				 l_2 = -29; end
		3846: begin l_1 = +19;
				 l_2 = +30; end
		2940: begin l_1 = +19;
				 l_2 = -30; end
		3371: begin l_1 = -19;
				 l_2 = +30; end
		2465: begin l_1 = -19;
				 l_2 = -30; end
		4299: begin l_1 = +19;
				 l_2 = +31; end
		2487: begin l_1 = +19;
				 l_2 = -31; end
		3824: begin l_1 = -19;
				 l_2 = +31; end
		2012: begin l_1 = -19;
				 l_2 = -31; end
		5205: begin l_1 = +19;
				 l_2 = +32; end
		1581: begin l_1 = +19;
				 l_2 = -32; end
		4730: begin l_1 = -19;
				 l_2 = +32; end
		1106: begin l_1 = -19;
				 l_2 = -32; end
		706: begin l_1 = +19;
				 l_2 = +33; end
		6080: begin l_1 = +19;
				 l_2 = -33; end
		231: begin l_1 = -19;
				 l_2 = +33; end
		5605: begin l_1 = -19;
				 l_2 = -33; end
		1425: begin l_1 = -20;
				 l_2 = +22; end
		4886: begin l_1 = -20;
				 l_2 = -21; end
		2375: begin l_1 = +20;
				 l_2 = +22; end
		3936: begin l_1 = -20;
				 l_2 = -22; end
		4275: begin l_1 = +20;
				 l_2 = +23; end
		2986: begin l_1 = +20;
				 l_2 = -23; end
		3325: begin l_1 = -20;
				 l_2 = +23; end
		2036: begin l_1 = -20;
				 l_2 = -23; end
		1764: begin l_1 = +20;
				 l_2 = +24; end
		5497: begin l_1 = +20;
				 l_2 = -24; end
		814: begin l_1 = -20;
				 l_2 = +24; end
		4547: begin l_1 = -20;
				 l_2 = -24; end
		3053: begin l_1 = +20;
				 l_2 = +25; end
		4208: begin l_1 = +20;
				 l_2 = -25; end
		2103: begin l_1 = -20;
				 l_2 = +25; end
		3258: begin l_1 = -20;
				 l_2 = -25; end
		5631: begin l_1 = +20;
				 l_2 = +26; end
		1630: begin l_1 = +20;
				 l_2 = -26; end
		4681: begin l_1 = -20;
				 l_2 = +26; end
		680: begin l_1 = -20;
				 l_2 = -26; end
		4476: begin l_1 = +20;
				 l_2 = +27; end
		2785: begin l_1 = +20;
				 l_2 = -27; end
		3526: begin l_1 = -20;
				 l_2 = +27; end
		1835: begin l_1 = -20;
				 l_2 = -27; end
		2166: begin l_1 = +20;
				 l_2 = +28; end
		5095: begin l_1 = +20;
				 l_2 = -28; end
		1216: begin l_1 = -20;
				 l_2 = +28; end
		4145: begin l_1 = -20;
				 l_2 = -28; end
		3857: begin l_1 = +20;
				 l_2 = +29; end
		3404: begin l_1 = +20;
				 l_2 = -29; end
		2907: begin l_1 = -20;
				 l_2 = +29; end
		2454: begin l_1 = -20;
				 l_2 = -29; end
		928: begin l_1 = +20;
				 l_2 = +30; end
		22: begin l_1 = +20;
				 l_2 = -30; end
		6289: begin l_1 = -20;
				 l_2 = +30; end
		5383: begin l_1 = -20;
				 l_2 = -30; end
		1381: begin l_1 = +20;
				 l_2 = +31; end
		5880: begin l_1 = +20;
				 l_2 = -31; end
		431: begin l_1 = -20;
				 l_2 = +31; end
		4930: begin l_1 = -20;
				 l_2 = -31; end
		2287: begin l_1 = +20;
				 l_2 = +32; end
		4974: begin l_1 = +20;
				 l_2 = -32; end
		1337: begin l_1 = -20;
				 l_2 = +32; end
		4024: begin l_1 = -20;
				 l_2 = -32; end
		4099: begin l_1 = +20;
				 l_2 = +33; end
		3162: begin l_1 = +20;
				 l_2 = -33; end
		3149: begin l_1 = -20;
				 l_2 = +33; end
		2212: begin l_1 = -20;
				 l_2 = -33; end
		2850: begin l_1 = -21;
				 l_2 = +23; end
		3461: begin l_1 = -21;
				 l_2 = -22; end
		4750: begin l_1 = +21;
				 l_2 = +23; end
		1561: begin l_1 = -21;
				 l_2 = -23; end
		2239: begin l_1 = +21;
				 l_2 = +24; end
		5972: begin l_1 = +21;
				 l_2 = -24; end
		339: begin l_1 = -21;
				 l_2 = +24; end
		4072: begin l_1 = -21;
				 l_2 = -24; end
		3528: begin l_1 = +21;
				 l_2 = +25; end
		4683: begin l_1 = +21;
				 l_2 = -25; end
		1628: begin l_1 = -21;
				 l_2 = +25; end
		2783: begin l_1 = -21;
				 l_2 = -25; end
		6106: begin l_1 = +21;
				 l_2 = +26; end
		2105: begin l_1 = +21;
				 l_2 = -26; end
		4206: begin l_1 = -21;
				 l_2 = +26; end
		205: begin l_1 = -21;
				 l_2 = -26; end
		4951: begin l_1 = +21;
				 l_2 = +27; end
		3260: begin l_1 = +21;
				 l_2 = -27; end
		3051: begin l_1 = -21;
				 l_2 = +27; end
		1360: begin l_1 = -21;
				 l_2 = -27; end
		2641: begin l_1 = +21;
				 l_2 = +28; end
		5570: begin l_1 = +21;
				 l_2 = -28; end
		741: begin l_1 = -21;
				 l_2 = +28; end
		3670: begin l_1 = -21;
				 l_2 = -28; end
		4332: begin l_1 = +21;
				 l_2 = +29; end
		3879: begin l_1 = +21;
				 l_2 = -29; end
		2432: begin l_1 = -21;
				 l_2 = +29; end
		1979: begin l_1 = -21;
				 l_2 = -29; end
		1403: begin l_1 = +21;
				 l_2 = +30; end
		497: begin l_1 = +21;
				 l_2 = -30; end
		5814: begin l_1 = -21;
				 l_2 = +30; end
		4908: begin l_1 = -21;
				 l_2 = -30; end
		1856: begin l_1 = +21;
				 l_2 = +31; end
		44: begin l_1 = +21;
				 l_2 = -31; end
		6267: begin l_1 = -21;
				 l_2 = +31; end
		4455: begin l_1 = -21;
				 l_2 = -31; end
		2762: begin l_1 = +21;
				 l_2 = +32; end
		5449: begin l_1 = +21;
				 l_2 = -32; end
		862: begin l_1 = -21;
				 l_2 = +32; end
		3549: begin l_1 = -21;
				 l_2 = -32; end
		4574: begin l_1 = +21;
				 l_2 = +33; end
		3637: begin l_1 = +21;
				 l_2 = -33; end
		2674: begin l_1 = -21;
				 l_2 = +33; end
		1737: begin l_1 = -21;
				 l_2 = -33; end
		5700: begin l_1 = -22;
				 l_2 = +24; end
		611: begin l_1 = -22;
				 l_2 = -23; end
		3189: begin l_1 = +22;
				 l_2 = +24; end
		3122: begin l_1 = -22;
				 l_2 = -24; end
		4478: begin l_1 = +22;
				 l_2 = +25; end
		5633: begin l_1 = +22;
				 l_2 = -25; end
		678: begin l_1 = -22;
				 l_2 = +25; end
		1833: begin l_1 = -22;
				 l_2 = -25; end
		745: begin l_1 = +22;
				 l_2 = +26; end
		3055: begin l_1 = +22;
				 l_2 = -26; end
		3256: begin l_1 = -22;
				 l_2 = +26; end
		5566: begin l_1 = -22;
				 l_2 = -26; end
		5901: begin l_1 = +22;
				 l_2 = +27; end
		4210: begin l_1 = +22;
				 l_2 = -27; end
		2101: begin l_1 = -22;
				 l_2 = +27; end
		410: begin l_1 = -22;
				 l_2 = -27; end
		3591: begin l_1 = +22;
				 l_2 = +28; end
		209: begin l_1 = +22;
				 l_2 = -28; end
		6102: begin l_1 = -22;
				 l_2 = +28; end
		2720: begin l_1 = -22;
				 l_2 = -28; end
		5282: begin l_1 = +22;
				 l_2 = +29; end
		4829: begin l_1 = +22;
				 l_2 = -29; end
		1482: begin l_1 = -22;
				 l_2 = +29; end
		1029: begin l_1 = -22;
				 l_2 = -29; end
		2353: begin l_1 = +22;
				 l_2 = +30; end
		1447: begin l_1 = +22;
				 l_2 = -30; end
		4864: begin l_1 = -22;
				 l_2 = +30; end
		3958: begin l_1 = -22;
				 l_2 = -30; end
		2806: begin l_1 = +22;
				 l_2 = +31; end
		994: begin l_1 = +22;
				 l_2 = -31; end
		5317: begin l_1 = -22;
				 l_2 = +31; end
		3505: begin l_1 = -22;
				 l_2 = -31; end
		3712: begin l_1 = +22;
				 l_2 = +32; end
		88: begin l_1 = +22;
				 l_2 = -32; end
		6223: begin l_1 = -22;
				 l_2 = +32; end
		2599: begin l_1 = -22;
				 l_2 = -32; end
		5524: begin l_1 = +22;
				 l_2 = +33; end
		4587: begin l_1 = +22;
				 l_2 = -33; end
		1724: begin l_1 = -22;
				 l_2 = +33; end
		787: begin l_1 = -22;
				 l_2 = -33; end
		5089: begin l_1 = -23;
				 l_2 = +25; end
		1222: begin l_1 = -23;
				 l_2 = -24; end
		67: begin l_1 = +23;
				 l_2 = +25; end
		6244: begin l_1 = -23;
				 l_2 = -25; end
		2645: begin l_1 = +23;
				 l_2 = +26; end
		4955: begin l_1 = +23;
				 l_2 = -26; end
		1356: begin l_1 = -23;
				 l_2 = +26; end
		3666: begin l_1 = -23;
				 l_2 = -26; end
		1490: begin l_1 = +23;
				 l_2 = +27; end
		6110: begin l_1 = +23;
				 l_2 = -27; end
		201: begin l_1 = -23;
				 l_2 = +27; end
		4821: begin l_1 = -23;
				 l_2 = -27; end
		5491: begin l_1 = +23;
				 l_2 = +28; end
		2109: begin l_1 = +23;
				 l_2 = -28; end
		4202: begin l_1 = -23;
				 l_2 = +28; end
		820: begin l_1 = -23;
				 l_2 = -28; end
		871: begin l_1 = +23;
				 l_2 = +29; end
		418: begin l_1 = +23;
				 l_2 = -29; end
		5893: begin l_1 = -23;
				 l_2 = +29; end
		5440: begin l_1 = -23;
				 l_2 = -29; end
		4253: begin l_1 = +23;
				 l_2 = +30; end
		3347: begin l_1 = +23;
				 l_2 = -30; end
		2964: begin l_1 = -23;
				 l_2 = +30; end
		2058: begin l_1 = -23;
				 l_2 = -30; end
		4706: begin l_1 = +23;
				 l_2 = +31; end
		2894: begin l_1 = +23;
				 l_2 = -31; end
		3417: begin l_1 = -23;
				 l_2 = +31; end
		1605: begin l_1 = -23;
				 l_2 = -31; end
		5612: begin l_1 = +23;
				 l_2 = +32; end
		1988: begin l_1 = +23;
				 l_2 = -32; end
		4323: begin l_1 = -23;
				 l_2 = +32; end
		699: begin l_1 = -23;
				 l_2 = -32; end
		1113: begin l_1 = +23;
				 l_2 = +33; end
		176: begin l_1 = +23;
				 l_2 = -33; end
		6135: begin l_1 = -23;
				 l_2 = +33; end
		5198: begin l_1 = -23;
				 l_2 = -33; end
		3867: begin l_1 = -24;
				 l_2 = +26; end
		2444: begin l_1 = -24;
				 l_2 = -25; end
		134: begin l_1 = +24;
				 l_2 = +26; end
		6177: begin l_1 = -24;
				 l_2 = -26; end
		5290: begin l_1 = +24;
				 l_2 = +27; end
		3599: begin l_1 = +24;
				 l_2 = -27; end
		2712: begin l_1 = -24;
				 l_2 = +27; end
		1021: begin l_1 = -24;
				 l_2 = -27; end
		2980: begin l_1 = +24;
				 l_2 = +28; end
		5909: begin l_1 = +24;
				 l_2 = -28; end
		402: begin l_1 = -24;
				 l_2 = +28; end
		3331: begin l_1 = -24;
				 l_2 = -28; end
		4671: begin l_1 = +24;
				 l_2 = +29; end
		4218: begin l_1 = +24;
				 l_2 = -29; end
		2093: begin l_1 = -24;
				 l_2 = +29; end
		1640: begin l_1 = -24;
				 l_2 = -29; end
		1742: begin l_1 = +24;
				 l_2 = +30; end
		836: begin l_1 = +24;
				 l_2 = -30; end
		5475: begin l_1 = -24;
				 l_2 = +30; end
		4569: begin l_1 = -24;
				 l_2 = -30; end
		2195: begin l_1 = +24;
				 l_2 = +31; end
		383: begin l_1 = +24;
				 l_2 = -31; end
		5928: begin l_1 = -24;
				 l_2 = +31; end
		4116: begin l_1 = -24;
				 l_2 = -31; end
		3101: begin l_1 = +24;
				 l_2 = +32; end
		5788: begin l_1 = +24;
				 l_2 = -32; end
		523: begin l_1 = -24;
				 l_2 = +32; end
		3210: begin l_1 = -24;
				 l_2 = -32; end
		4913: begin l_1 = +24;
				 l_2 = +33; end
		3976: begin l_1 = +24;
				 l_2 = -33; end
		2335: begin l_1 = -24;
				 l_2 = +33; end
		1398: begin l_1 = -24;
				 l_2 = -33; end
		1423: begin l_1 = -25;
				 l_2 = +27; end
		4888: begin l_1 = -25;
				 l_2 = -26; end
		268: begin l_1 = +25;
				 l_2 = +27; end
		6043: begin l_1 = -25;
				 l_2 = -27; end
		4269: begin l_1 = +25;
				 l_2 = +28; end
		887: begin l_1 = +25;
				 l_2 = -28; end
		5424: begin l_1 = -25;
				 l_2 = +28; end
		2042: begin l_1 = -25;
				 l_2 = -28; end
		5960: begin l_1 = +25;
				 l_2 = +29; end
		5507: begin l_1 = +25;
				 l_2 = -29; end
		804: begin l_1 = -25;
				 l_2 = +29; end
		351: begin l_1 = -25;
				 l_2 = -29; end
		3031: begin l_1 = +25;
				 l_2 = +30; end
		2125: begin l_1 = +25;
				 l_2 = -30; end
		4186: begin l_1 = -25;
				 l_2 = +30; end
		3280: begin l_1 = -25;
				 l_2 = -30; end
		3484: begin l_1 = +25;
				 l_2 = +31; end
		1672: begin l_1 = +25;
				 l_2 = -31; end
		4639: begin l_1 = -25;
				 l_2 = +31; end
		2827: begin l_1 = -25;
				 l_2 = -31; end
		4390: begin l_1 = +25;
				 l_2 = +32; end
		766: begin l_1 = +25;
				 l_2 = -32; end
		5545: begin l_1 = -25;
				 l_2 = +32; end
		1921: begin l_1 = -25;
				 l_2 = -32; end
		6202: begin l_1 = +25;
				 l_2 = +33; end
		5265: begin l_1 = +25;
				 l_2 = -33; end
		1046: begin l_1 = -25;
				 l_2 = +33; end
		109: begin l_1 = -25;
				 l_2 = -33; end
		2846: begin l_1 = -26;
				 l_2 = +28; end
		3465: begin l_1 = -26;
				 l_2 = -27; end
		536: begin l_1 = +26;
				 l_2 = +28; end
		5775: begin l_1 = -26;
				 l_2 = -28; end
		2227: begin l_1 = +26;
				 l_2 = +29; end
		1774: begin l_1 = +26;
				 l_2 = -29; end
		4537: begin l_1 = -26;
				 l_2 = +29; end
		4084: begin l_1 = -26;
				 l_2 = -29; end
		5609: begin l_1 = +26;
				 l_2 = +30; end
		4703: begin l_1 = +26;
				 l_2 = -30; end
		1608: begin l_1 = -26;
				 l_2 = +30; end
		702: begin l_1 = -26;
				 l_2 = -30; end
		6062: begin l_1 = +26;
				 l_2 = +31; end
		4250: begin l_1 = +26;
				 l_2 = -31; end
		2061: begin l_1 = -26;
				 l_2 = +31; end
		249: begin l_1 = -26;
				 l_2 = -31; end
		657: begin l_1 = +26;
				 l_2 = +32; end
		3344: begin l_1 = +26;
				 l_2 = -32; end
		2967: begin l_1 = -26;
				 l_2 = +32; end
		5654: begin l_1 = -26;
				 l_2 = -32; end
		2469: begin l_1 = +26;
				 l_2 = +33; end
		1532: begin l_1 = +26;
				 l_2 = -33; end
		4779: begin l_1 = -26;
				 l_2 = +33; end
		3842: begin l_1 = -26;
				 l_2 = -33; end
		5692: begin l_1 = -27;
				 l_2 = +29; end
		619: begin l_1 = -27;
				 l_2 = -28; end
		1072: begin l_1 = +27;
				 l_2 = +29; end
		5239: begin l_1 = -27;
				 l_2 = -29; end
		4454: begin l_1 = +27;
				 l_2 = +30; end
		3548: begin l_1 = +27;
				 l_2 = -30; end
		2763: begin l_1 = -27;
				 l_2 = +30; end
		1857: begin l_1 = -27;
				 l_2 = -30; end
		4907: begin l_1 = +27;
				 l_2 = +31; end
		3095: begin l_1 = +27;
				 l_2 = -31; end
		3216: begin l_1 = -27;
				 l_2 = +31; end
		1404: begin l_1 = -27;
				 l_2 = -31; end
		5813: begin l_1 = +27;
				 l_2 = +32; end
		2189: begin l_1 = +27;
				 l_2 = -32; end
		4122: begin l_1 = -27;
				 l_2 = +32; end
		498: begin l_1 = -27;
				 l_2 = -32; end
		1314: begin l_1 = +27;
				 l_2 = +33; end
		377: begin l_1 = +27;
				 l_2 = -33; end
		5934: begin l_1 = -27;
				 l_2 = +33; end
		4997: begin l_1 = -27;
				 l_2 = -33; end
		5073: begin l_1 = -28;
				 l_2 = +30; end
		1238: begin l_1 = -28;
				 l_2 = -29; end
		2144: begin l_1 = +28;
				 l_2 = +30; end
		4167: begin l_1 = -28;
				 l_2 = -30; end
		2597: begin l_1 = +28;
				 l_2 = +31; end
		785: begin l_1 = +28;
				 l_2 = -31; end
		5526: begin l_1 = -28;
				 l_2 = +31; end
		3714: begin l_1 = -28;
				 l_2 = -31; end
		3503: begin l_1 = +28;
				 l_2 = +32; end
		6190: begin l_1 = +28;
				 l_2 = -32; end
		121: begin l_1 = -28;
				 l_2 = +32; end
		2808: begin l_1 = -28;
				 l_2 = -32; end
		5315: begin l_1 = +28;
				 l_2 = +33; end
		4378: begin l_1 = +28;
				 l_2 = -33; end
		1933: begin l_1 = -28;
				 l_2 = +33; end
		996: begin l_1 = -28;
				 l_2 = -33; end
		3835: begin l_1 = -29;
				 l_2 = +31; end
		2476: begin l_1 = -29;
				 l_2 = -30; end
		4288: begin l_1 = +29;
				 l_2 = +31; end
		2023: begin l_1 = -29;
				 l_2 = -31; end
		5194: begin l_1 = +29;
				 l_2 = +32; end
		1570: begin l_1 = +29;
				 l_2 = -32; end
		4741: begin l_1 = -29;
				 l_2 = +32; end
		1117: begin l_1 = -29;
				 l_2 = -32; end
		695: begin l_1 = +29;
				 l_2 = +33; end
		6069: begin l_1 = +29;
				 l_2 = -33; end
		242: begin l_1 = -29;
				 l_2 = +33; end
		5616: begin l_1 = -29;
				 l_2 = -33; end
		1359: begin l_1 = -30;
				 l_2 = +32; end
		4952: begin l_1 = -30;
				 l_2 = -31; end
		2265: begin l_1 = +30;
				 l_2 = +32; end
		4046: begin l_1 = -30;
				 l_2 = -32; end
		4077: begin l_1 = +30;
				 l_2 = +33; end
		3140: begin l_1 = +30;
				 l_2 = -33; end
		3171: begin l_1 = -30;
				 l_2 = +33; end
		2234: begin l_1 = -30;
				 l_2 = -33; end
		2718: begin l_1 = -31;
				 l_2 = +33; end
		3593: begin l_1 = -31;
				 l_2 = -32; end
		4530: begin l_1 = +31;
				 l_2 = +33; end
		1781: begin l_1 = -31;
				 l_2 = -33; end
		5436: begin l_1 = +32;
				 l_2 = +33; end
		875: begin l_1 = -32;
				 l_2 = -33; end
		default: begin l_1 = 0;
					   l_2 = 0; end
	endcase
end

endmodule

// Product (AN) Code DEC_LUT_Decoder
// DEC_LUT_Decoder4bits.v
// Received codeword W = AN + E, E is double AWE (E = e1 + e2), +2^i or -2^i.
module DEC_LUT_Decoder4bits(W, N);
input 	[13:0]	W;
output	[3:0]	N;
parameter A = 665;

wire 	[3:0]	Q;
wire 	[9:0]	R;
assign Q = W / A;
assign R = W - (A * Q);

reg	signed	[14:0]	Delta;
always@(*) begin
	case(R)
		1: Delta = 15'sb000000000000001;
		664: Delta = 15'sb111111111111111;
		2: Delta = 15'sb000000000000010;
		663: Delta = 15'sb111111111111110;
		4: Delta = 15'sb000000000000100;
		661: Delta = 15'sb111111111111100;
		8: Delta = 15'sb000000000001000;
		657: Delta = 15'sb111111111111000;
		16: Delta = 15'sb000000000010000;
		649: Delta = 15'sb111111111110000;
		32: Delta = 15'sb000000000100000;
		633: Delta = 15'sb111111111100000;
		64: Delta = 15'sb000000001000000;
		601: Delta = 15'sb111111111000000;
		128: Delta = 15'sb000000010000000;
		537: Delta = 15'sb111111110000000;
		256: Delta = 15'sb000000100000000;
		409: Delta = 15'sb111111100000000;
		512: Delta = 15'sb000001000000000;
		153: Delta = 15'sb111111000000000;
		359: Delta = 15'sb000010000000000;
		306: Delta = 15'sb111110000000000;
		53: Delta = 15'sb000100000000000;
		612: Delta = 15'sb111100000000000;
		106: Delta = 15'sb001000000000000;
		559: Delta = 15'sb111000000000000;
		212: Delta = 15'sb010000000000000;
		453: Delta = 15'sb110000000000000;
		3: Delta = 15'sb000000000000011;
		662: Delta = 15'sb111111111111101;
		5: Delta = 15'sb000000000000101;
		660: Delta = 15'sb111111111111011;
		9: Delta = 15'sb000000000001001;
		658: Delta = 15'sb111111111111001;
		7: Delta = 15'sb000000000000111;
		656: Delta = 15'sb111111111110111;
		17: Delta = 15'sb000000000010001;
		650: Delta = 15'sb111111111110001;
		15: Delta = 15'sb000000000001111;
		648: Delta = 15'sb111111111101111;
		33: Delta = 15'sb000000000100001;
		634: Delta = 15'sb111111111100001;
		31: Delta = 15'sb000000000011111;
		632: Delta = 15'sb111111111011111;
		65: Delta = 15'sb000000001000001;
		602: Delta = 15'sb111111111000001;
		63: Delta = 15'sb000000000111111;
		600: Delta = 15'sb111111110111111;
		129: Delta = 15'sb000000010000001;
		538: Delta = 15'sb111111110000001;
		127: Delta = 15'sb000000001111111;
		536: Delta = 15'sb111111101111111;
		257: Delta = 15'sb000000100000001;
		410: Delta = 15'sb111111100000001;
		255: Delta = 15'sb000000011111111;
		408: Delta = 15'sb111111011111111;
		513: Delta = 15'sb000001000000001;
		154: Delta = 15'sb111111000000001;
		511: Delta = 15'sb000000111111111;
		152: Delta = 15'sb111110111111111;
		360: Delta = 15'sb000010000000001;
		307: Delta = 15'sb111110000000001;
		358: Delta = 15'sb000001111111111;
		305: Delta = 15'sb111101111111111;
		54: Delta = 15'sb000100000000001;
		613: Delta = 15'sb111100000000001;
		52: Delta = 15'sb000011111111111;
		611: Delta = 15'sb111011111111111;
		107: Delta = 15'sb001000000000001;
		560: Delta = 15'sb111000000000001;
		105: Delta = 15'sb000111111111111;
		558: Delta = 15'sb110111111111111;
		213: Delta = 15'sb010000000000001;
		454: Delta = 15'sb110000000000001;
		211: Delta = 15'sb001111111111111;
		452: Delta = 15'sb101111111111111;
		6: Delta = 15'sb000000000000110;
		659: Delta = 15'sb111111111111010;
		10: Delta = 15'sb000000000001010;
		655: Delta = 15'sb111111111110110;
		18: Delta = 15'sb000000000010010;
		651: Delta = 15'sb111111111110010;
		14: Delta = 15'sb000000000001110;
		647: Delta = 15'sb111111111101110;
		34: Delta = 15'sb000000000100010;
		635: Delta = 15'sb111111111100010;
		30: Delta = 15'sb000000000011110;
		631: Delta = 15'sb111111111011110;
		66: Delta = 15'sb000000001000010;
		603: Delta = 15'sb111111111000010;
		62: Delta = 15'sb000000000111110;
		599: Delta = 15'sb111111110111110;
		130: Delta = 15'sb000000010000010;
		539: Delta = 15'sb111111110000010;
		126: Delta = 15'sb000000001111110;
		535: Delta = 15'sb111111101111110;
		258: Delta = 15'sb000000100000010;
		411: Delta = 15'sb111111100000010;
		254: Delta = 15'sb000000011111110;
		407: Delta = 15'sb111111011111110;
		514: Delta = 15'sb000001000000010;
		155: Delta = 15'sb111111000000010;
		510: Delta = 15'sb000000111111110;
		151: Delta = 15'sb111110111111110;
		361: Delta = 15'sb000010000000010;
		308: Delta = 15'sb111110000000010;
		357: Delta = 15'sb000001111111110;
		304: Delta = 15'sb111101111111110;
		55: Delta = 15'sb000100000000010;
		614: Delta = 15'sb111100000000010;
		51: Delta = 15'sb000011111111110;
		610: Delta = 15'sb111011111111110;
		108: Delta = 15'sb001000000000010;
		561: Delta = 15'sb111000000000010;
		104: Delta = 15'sb000111111111110;
		557: Delta = 15'sb110111111111110;
		214: Delta = 15'sb010000000000010;
		455: Delta = 15'sb110000000000010;
		210: Delta = 15'sb001111111111110;
		451: Delta = 15'sb101111111111110;
		12: Delta = 15'sb000000000001100;
		653: Delta = 15'sb111111111110100;
		20: Delta = 15'sb000000000010100;
		645: Delta = 15'sb111111111101100;
		36: Delta = 15'sb000000000100100;
		637: Delta = 15'sb111111111100100;
		28: Delta = 15'sb000000000011100;
		629: Delta = 15'sb111111111011100;
		68: Delta = 15'sb000000001000100;
		605: Delta = 15'sb111111111000100;
		60: Delta = 15'sb000000000111100;
		597: Delta = 15'sb111111110111100;
		132: Delta = 15'sb000000010000100;
		541: Delta = 15'sb111111110000100;
		124: Delta = 15'sb000000001111100;
		533: Delta = 15'sb111111101111100;
		260: Delta = 15'sb000000100000100;
		413: Delta = 15'sb111111100000100;
		252: Delta = 15'sb000000011111100;
		405: Delta = 15'sb111111011111100;
		516: Delta = 15'sb000001000000100;
		157: Delta = 15'sb111111000000100;
		508: Delta = 15'sb000000111111100;
		149: Delta = 15'sb111110111111100;
		363: Delta = 15'sb000010000000100;
		310: Delta = 15'sb111110000000100;
		355: Delta = 15'sb000001111111100;
		302: Delta = 15'sb111101111111100;
		57: Delta = 15'sb000100000000100;
		616: Delta = 15'sb111100000000100;
		49: Delta = 15'sb000011111111100;
		608: Delta = 15'sb111011111111100;
		110: Delta = 15'sb001000000000100;
		563: Delta = 15'sb111000000000100;
		102: Delta = 15'sb000111111111100;
		555: Delta = 15'sb110111111111100;
		216: Delta = 15'sb010000000000100;
		457: Delta = 15'sb110000000000100;
		208: Delta = 15'sb001111111111100;
		449: Delta = 15'sb101111111111100;
		24: Delta = 15'sb000000000011000;
		641: Delta = 15'sb111111111101000;
		40: Delta = 15'sb000000000101000;
		625: Delta = 15'sb111111111011000;
		72: Delta = 15'sb000000001001000;
		609: Delta = 15'sb111111111001000;
		56: Delta = 15'sb000000000111000;
		593: Delta = 15'sb111111110111000;
		136: Delta = 15'sb000000010001000;
		545: Delta = 15'sb111111110001000;
		120: Delta = 15'sb000000001111000;
		529: Delta = 15'sb111111101111000;
		264: Delta = 15'sb000000100001000;
		417: Delta = 15'sb111111100001000;
		248: Delta = 15'sb000000011111000;
		401: Delta = 15'sb111111011111000;
		520: Delta = 15'sb000001000001000;
		161: Delta = 15'sb111111000001000;
		504: Delta = 15'sb000000111111000;
		145: Delta = 15'sb111110111111000;
		367: Delta = 15'sb000010000001000;
		314: Delta = 15'sb111110000001000;
		351: Delta = 15'sb000001111111000;
		298: Delta = 15'sb111101111111000;
		61: Delta = 15'sb000100000001000;
		620: Delta = 15'sb111100000001000;
		45: Delta = 15'sb000011111111000;
		604: Delta = 15'sb111011111111000;
		114: Delta = 15'sb001000000001000;
		567: Delta = 15'sb111000000001000;
		98: Delta = 15'sb000111111111000;
		551: Delta = 15'sb110111111111000;
		220: Delta = 15'sb010000000001000;
		461: Delta = 15'sb110000000001000;
		204: Delta = 15'sb001111111111000;
		445: Delta = 15'sb101111111111000;
		48: Delta = 15'sb000000000110000;
		617: Delta = 15'sb111111111010000;
		80: Delta = 15'sb000000001010000;
		585: Delta = 15'sb111111110110000;
		144: Delta = 15'sb000000010010000;
		553: Delta = 15'sb111111110010000;
		112: Delta = 15'sb000000001110000;
		521: Delta = 15'sb111111101110000;
		272: Delta = 15'sb000000100010000;
		425: Delta = 15'sb111111100010000;
		240: Delta = 15'sb000000011110000;
		393: Delta = 15'sb111111011110000;
		528: Delta = 15'sb000001000010000;
		169: Delta = 15'sb111111000010000;
		496: Delta = 15'sb000000111110000;
		137: Delta = 15'sb111110111110000;
		375: Delta = 15'sb000010000010000;
		322: Delta = 15'sb111110000010000;
		343: Delta = 15'sb000001111110000;
		290: Delta = 15'sb111101111110000;
		69: Delta = 15'sb000100000010000;
		628: Delta = 15'sb111100000010000;
		37: Delta = 15'sb000011111110000;
		596: Delta = 15'sb111011111110000;
		122: Delta = 15'sb001000000010000;
		575: Delta = 15'sb111000000010000;
		90: Delta = 15'sb000111111110000;
		543: Delta = 15'sb110111111110000;
		228: Delta = 15'sb010000000010000;
		469: Delta = 15'sb110000000010000;
		196: Delta = 15'sb001111111110000;
		437: Delta = 15'sb101111111110000;
		96: Delta = 15'sb000000001100000;
		569: Delta = 15'sb111111110100000;
		160: Delta = 15'sb000000010100000;
		505: Delta = 15'sb111111101100000;
		288: Delta = 15'sb000000100100000;
		441: Delta = 15'sb111111100100000;
		224: Delta = 15'sb000000011100000;
		377: Delta = 15'sb111111011100000;
		544: Delta = 15'sb000001000100000;
		185: Delta = 15'sb111111000100000;
		480: Delta = 15'sb000000111100000;
		121: Delta = 15'sb111110111100000;
		391: Delta = 15'sb000010000100000;
		338: Delta = 15'sb111110000100000;
		327: Delta = 15'sb000001111100000;
		274: Delta = 15'sb111101111100000;
		85: Delta = 15'sb000100000100000;
		644: Delta = 15'sb111100000100000;
		21: Delta = 15'sb000011111100000;
		580: Delta = 15'sb111011111100000;
		138: Delta = 15'sb001000000100000;
		591: Delta = 15'sb111000000100000;
		74: Delta = 15'sb000111111100000;
		527: Delta = 15'sb110111111100000;
		244: Delta = 15'sb010000000100000;
		485: Delta = 15'sb110000000100000;
		180: Delta = 15'sb001111111100000;
		421: Delta = 15'sb101111111100000;
		192: Delta = 15'sb000000011000000;
		473: Delta = 15'sb111111101000000;
		320: Delta = 15'sb000000101000000;
		345: Delta = 15'sb111111011000000;
		576: Delta = 15'sb000001001000000;
		217: Delta = 15'sb111111001000000;
		448: Delta = 15'sb000000111000000;
		89: Delta = 15'sb111110111000000;
		423: Delta = 15'sb000010001000000;
		370: Delta = 15'sb111110001000000;
		295: Delta = 15'sb000001111000000;
		242: Delta = 15'sb111101111000000;
		117: Delta = 15'sb000100001000000;
		11: Delta = 15'sb111100001000000;
		654: Delta = 15'sb000011111000000;
		548: Delta = 15'sb111011111000000;
		170: Delta = 15'sb001000001000000;
		623: Delta = 15'sb111000001000000;
		42: Delta = 15'sb000111111000000;
		495: Delta = 15'sb110111111000000;
		276: Delta = 15'sb010000001000000;
		517: Delta = 15'sb110000001000000;
		148: Delta = 15'sb001111111000000;
		389: Delta = 15'sb101111111000000;
		384: Delta = 15'sb000000110000000;
		281: Delta = 15'sb111111010000000;
		640: Delta = 15'sb000001010000000;
		25: Delta = 15'sb111110110000000;
		487: Delta = 15'sb000010010000000;
		434: Delta = 15'sb111110010000000;
		231: Delta = 15'sb000001110000000;
		178: Delta = 15'sb111101110000000;
		181: Delta = 15'sb000100010000000;
		75: Delta = 15'sb111100010000000;
		590: Delta = 15'sb000011110000000;
		484: Delta = 15'sb111011110000000;
		234: Delta = 15'sb001000010000000;
		22: Delta = 15'sb111000010000000;
		643: Delta = 15'sb000111110000000;
		431: Delta = 15'sb110111110000000;
		340: Delta = 15'sb010000010000000;
		581: Delta = 15'sb110000010000000;
		84: Delta = 15'sb001111110000000;
		325: Delta = 15'sb101111110000000;
		103: Delta = 15'sb000001100000000;
		562: Delta = 15'sb111110100000000;
		615: Delta = 15'sb000010100000000;
		50: Delta = 15'sb111101100000000;
		309: Delta = 15'sb000100100000000;
		203: Delta = 15'sb111100100000000;
		462: Delta = 15'sb000011100000000;
		356: Delta = 15'sb111011100000000;
		362: Delta = 15'sb001000100000000;
		150: Delta = 15'sb111000100000000;
		515: Delta = 15'sb000111100000000;
		303: Delta = 15'sb110111100000000;
		468: Delta = 15'sb010000100000000;
		44: Delta = 15'sb110000100000000;
		621: Delta = 15'sb001111100000000;
		197: Delta = 15'sb101111100000000;
		206: Delta = 15'sb000011000000000;
		459: Delta = 15'sb111101000000000;
		565: Delta = 15'sb000101000000000;
		100: Delta = 15'sb111011000000000;
		618: Delta = 15'sb001001000000000;
		406: Delta = 15'sb111001000000000;
		259: Delta = 15'sb000111000000000;
		47: Delta = 15'sb110111000000000;
		59: Delta = 15'sb010001000000000;
		300: Delta = 15'sb110001000000000;
		365: Delta = 15'sb001111000000000;
		606: Delta = 15'sb101111000000000;
		412: Delta = 15'sb000110000000000;
		253: Delta = 15'sb111010000000000;
		465: Delta = 15'sb001010000000000;
		200: Delta = 15'sb110110000000000;
		571: Delta = 15'sb010010000000000;
		147: Delta = 15'sb110010000000000;
		518: Delta = 15'sb001110000000000;
		94: Delta = 15'sb101110000000000;
		159: Delta = 15'sb001100000000000;
		506: Delta = 15'sb110100000000000;
		265: Delta = 15'sb010100000000000;
		400: Delta = 15'sb101100000000000;
		318: Delta = 15'sb011000000000000;
		347: Delta = 15'sb101000000000000;
		default: Delta =15'sb0;
	endcase
end

assign N = (W - Delta) / A;

endmodule
